###############################################################################
#TSMC Library/IP Product
#Filename: tcbn40lpbwp_9lm6X2ZRDL.lef
#Technology: CLN40LP
#Product Type: Standard Cell
#Product Name: tcbn40lpbwp
#Version: 120c
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################
# DESIGN RULE DOCUMENT: T-N45-CL-DR-001 V1.2

#+
#+Note:
#+      1. Please use Encounter 7.1USR1(or above) for advanced rule modeling support.
#+      2. Antenna ratio defined in OXIDE2 is for OD25/OD33.
#+      3. Please use Captable to get the correct RC values.
#+	4. Set the following command in Encounter to get the correct RC values from 
#+	   Captable when executing NanoRoute.
#+	   setNanoRouteMode -envResistanceFromCapTable true
#+      5. Using TSMC utility for dummy fill is strongly recommended.
#+	6. Please refer to T-N40-CL-RP-020 for DFM via usage.
#+
VERSION	5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS 
        # Begin added by Michael Oduoza
	LAYER LEF58_TYPE STRING ;
	LAYER LEF58_WIDTH STRING ;
	LAYER LEF58_ENCLOSURE STRING ;
 	# End added by Michael Oduoza
	LAYER LEF58_ENCLOSUREEDGE STRING ;
	LAYER LEF58_SPACING STRING ;
	LAYER LEF58_AREA STRING ;
	LIBRARY LEF58_MAXVIASTACK STRING "MAXVIASTACK 4 NOSINGLE RANGE M1 M7 ;" ;
END PROPERTYDEFINITIONS

LAYER VTH_P
	TYPE IMPLANT ;
	WIDTH 0.18 ;
	SPACING 0.18 ;
END VTH_P

LAYER VTH_N
	TYPE IMPLANT ;
	WIDTH 0.18 ;
	SPACING 0.18 ;
END VTH_N

LAYER VTL_P
	TYPE IMPLANT ;
	WIDTH 0.18 ;
	SPACING 0.18 ;
END VTL_P

LAYER VTL_N
	TYPE IMPLANT ;
	WIDTH 0.18 ;
	SPACING 0.18 ;
END VTL_N

# Begin added by Michael Oduoza
LAYER RELAY_METAL
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END RELAY_METAL

LAYER RELAY_VIA
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END RELAY_VIA

LAYER NEMANC
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END NEMANC

LAYER NEMCHAN
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END NEMCHAN

LAYER NEMBODY
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END NEMBODY

LAYER NEMCONT
  TYPE MASTERSLICE ;
  #DIRECTION HORIZONTAL ;
  WIDTH 0.07 ;
  #AREA 0.0215 ;
  #SPACING 0.07 ;
END NEMCONT
# End added by Michael Oduoza

LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
END CO

LAYER M1
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 0.535 ;
	THICKNESS 0.125 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.08	0.08	0.08	0.08
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.14	0.14	0.14
	WIDTH 0.62		0.07	0.12	0.14	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.14	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.08 ENDOFLINE 0.09 WITHIN 0.025 PARALLELEDGE 0.08 WITHIN 0.07 MINLENGTH 0.07 ; " ;
	AREA 0.0215 ;
	MINENCLOSEDAREA 0.2 ;
	PROPERTY LEF58_AREA "AREA 0.055 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.3080000000 ;
        CAPACITANCE CPERSQDIST	0.0002317460 ;
        EDGECAPACITANCE	0.0000808000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.07119	1.14910	1.20519	1.21609	1.22155	1.22458 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	14.65003	13.51795	11.26055	10.53159	10.10889	9.85397 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	30.86577	33.11056	34.72680	35.04107	35.19820	35.28550 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.07119	1.14910	1.20519	1.21609	1.22155	1.22458 ;
END M1

LAYER VIA1
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;
	PROPERTY LEF58_ENCLOSUREEDGE "ENCLOSUREEDGE BELOW 0.015 WIDTH 0.11 PARALLEL 0.27 WITHIN 0.08 EXCEPTEXTRACUT ;" ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA1

LAYER M2
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.14 ;
	OFFSET 0.07 ;
        HEIGHT 0.735 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000730000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	8.07330	7.37682	6.00661	5.55933	5.29799	5.13953 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M2

LAYER VIA2
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA2

LAYER M3
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 0.935 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000730000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.78447	6.88453	5.13176	4.52648	4.15850	3.92851 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M3

LAYER VIA3
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA3

LAYER M4
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.14 ;
	OFFSET 0.07 ;
        HEIGHT 1.135 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000730000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.66324	6.67939	4.74864	4.05673	3.62354	3.34586 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M4

LAYER VIA4
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA4

LAYER M5
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 1.335 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000730000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.60419	6.57371	4.53752	3.78921	3.31016	2.99658 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M5

LAYER VIA5
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA5

LAYER M6
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.14 ;
	OFFSET 0.07 ;
        HEIGHT 1.535 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 ;
	MINIMUMCUT 2 WIDTH 0.21 LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 LENGTH 7.0 WITHIN 7.101 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000730000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.56754	6.50734	4.40119	3.61285	3.09928	2.75703 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M6

LAYER VIA6
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA6

LAYER M7
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 1.735 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 2 WIDTH 1.8 WITHIN 1.701 FROMABOVE ;
	MINIMUMCUT 2 WIDTH 0.21 FROMBELOW LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 FROMBELOW LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 FROMBELOW LENGTH 7.0 WITHIN 7.101 ;
	MINIMUMCUT 2 WIDTH 3.0 FROMABOVE LENGTH 10.0 WITHIN 5.001 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000732000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.54402	6.46312	4.30689	3.48854	2.94786	2.58199 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M7

# Begin edited by Michael Oduoza
LAYER VIA7
	TYPE CUT ;
	SPACING 0.095 ;
	SPACING 0.09 ADJACENTCUTS 3 WITHIN 0.098 ;
	SPACING 0.11 PARALLELOVERLAP ;
	SPACING 0.07 SAMENET ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	18.14059 ;
        DCCURRENTDENSITY	AVERAGE	18.14059 ;
END VIA7

LAYER M8
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 1.735 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 2 WIDTH 1.8 WITHIN 1.701 FROMABOVE ;
	MINIMUMCUT 2 WIDTH 0.21 FROMBELOW LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 FROMBELOW LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 FROMBELOW LENGTH 7.0 WITHIN 7.101 ;
	MINIMUMCUT 2 WIDTH 3.0 FROMABOVE LENGTH 10.0 WITHIN 5.001 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000732000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.54402	6.46312	4.30689	3.48854	2.94786	2.58199 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M8

LAYER VIA8
	TYPE CUT ;
	SPACING 0.34 ;
	SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	29.31146 ;
        DCCURRENTDENSITY	AVERAGE	29.31146 ;
END VIA8

LAYER M9
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.14 ;
	OFFSET 0 ;
        HEIGHT 1.735 ;
	THICKNESS 0.14 ;
	FILLACTIVESPACING 0.6 ;
	WIDTH 0.07 ;
	MAXWIDTH 4.50 ;
	SPACINGTABLE
	PARALLELRUNLENGTH 	0.00	0.27	0.40	0.62	1.50
	WIDTH 0.00		0.07	0.07	0.07	0.07	0.07
	WIDTH 0.17		0.07	0.10	0.10	0.10	0.10
	WIDTH 0.24		0.07	0.12	0.12	0.12	0.12
	WIDTH 0.31		0.07	0.12	0.15	0.15	0.15
	WIDTH 0.62		0.07	0.12	0.15	0.21	0.21
	WIDTH 1.50		0.07	0.12	0.15	0.21	0.50 ;
	PROPERTY LEF58_SPACING "SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.10 WITHIN 0.10 MINLENGTH 0.07 ; SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.10 MINLENGTH 0.07 ENCLOSECUT BELOW 0.05 CUTSPACING 0.15 ; " ;
	AREA 0.027 ;
	MINENCLOSEDAREA 0.20 ;
	PROPERTY LEF58_AREA "AREA 0.06 EXCEPTEDGELENGTH 0.17 EXCEPTMINSIZE 0.07 0.17 ;" ;

	MINSTEP 0.07 MAXEDGES 1 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 85.0 ;
	DENSITYCHECKWINDOW 125 125 ;
	DENSITYCHECKSTEP 62.5 ;

	MINIMUMCUT 2 WIDTH 0.21 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 4 WIDTH 0.55 WITHIN 0.141 FROMBELOW ;
	MINIMUMCUT 2 WIDTH 1.8 WITHIN 1.701 FROMABOVE ;
	MINIMUMCUT 2 WIDTH 0.21 FROMBELOW LENGTH 0.21 WITHIN 1.141 ;
	MINIMUMCUT 2 WIDTH 1.4 FROMBELOW LENGTH 1.4 WITHIN 2.801 ;
	MINIMUMCUT 2 WIDTH 2.1 FROMBELOW LENGTH 7.0 WITHIN 7.101 ;
	MINIMUMCUT 2 WIDTH 3.0 FROMABOVE LENGTH 10.0 WITHIN 5.001 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

        RESISTANCE RPERSQ	0.2780000000 ;
        CAPACITANCE CPERSQDIST	0.0003444444 ;
        EDGECAPACITANCE	0.0000732000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	7.54402	6.46312	4.30689	3.48854	2.94786	2.58199 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	17.28483	18.54191	19.44701	19.62300	19.71099	19.75988 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	0.07000	0.14000	0.50000	1.00000	2.00000	4.50000 ;
              TABLEENTRIES	1.16024	1.24462	1.30537	1.31719	1.32309	1.32637 ;
END M9
# End edited by Michael Oduoza

LAYER RV
	TYPE CUT ;
	SPACING 2.0 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 200 ) ( 0.000025 400.00207 ) ( 0.2 416.6 ) ( 0.5 441.5 ) ( 1 483 ) ( 1.5 524.5 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 400.00207 ) ( 0.2 416.6 ) ( 0.5 441.5 ) ( 1 483 ) ( 1.5 524.5 ) ) ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              TABLEENTRIES	1.66667 ;
        DCCURRENTDENSITY	AVERAGE	1.66667 ;
END RV

LAYER AP
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	OFFSET 0.07 ;
	PITCH 5.0 ;
	WIDTH 2.0 ;
	MAXWIDTH 35.0 ;
	SPACING 2.0 ;
        HEIGHT 5.035 ;
	THICKNESS 1.45 ;

	MINIMUMDENSITY 10.0 ;
	MAXIMUMDENSITY 70.0 ;
	DENSITYCHECKWINDOW 100 100 ;
	DENSITYCHECKSTEP 50 ;

	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0 2000 ) ( 0.000025 30000.2 ) ( 0.2 31600.0 ) ( 0.5 34000.0 ) ( 1 38000 ) ( 1.5 42000.0 ) ) ;
	ANTENNAMODEL OXIDE2 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.000025 30000.2 ) ( 0.2 31600.0 ) ( 0.5 34000.0 ) ( 1 38000 ) ( 1.5 42000.0 ) ) ;

        RESISTANCE RPERSQ	0.0210000000 ;
        CAPACITANCE CPERSQDIST	0.0000611111 ;
        EDGECAPACITANCE	0.0000595000 ;

        ACCURRENTDENSITY	AVERAGE
              FREQUENCY	500 ;
              WIDTH    	2.00000	5.00000	8.00000	15.00000	20.00000	35.00000 ;
              TABLEENTRIES	3.00000	3.00000	3.00000	3.00000	3.00000	3.00000 ;
        ACCURRENTDENSITY	RMS
              FREQUENCY	500 ;
              WIDTH    	2.00000	5.00000	8.00000	15.00000	20.00000	35.00000 ;
              TABLEENTRIES	5.77325	4.57735	4.22583	3.93074	3.84227	3.72544 ;
        ACCURRENTDENSITY	PEAK
              FREQUENCY	500 ;
              WIDTH    	2.00000	5.00000	8.00000	15.00000	20.00000	35.00000 ;
              TABLEENTRIES	82.02439	82.02439	82.02439	82.02439	82.02439	82.02439 ;
        DCCURRENTDENSITY	AVERAGE
              WIDTH    	2.00000	5.00000	8.00000	15.00000	20.00000	35.00000 ;
              TABLEENTRIES	3.00000	3.00000	3.00000	3.00000	3.00000	3.00000 ;
END AP

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP
VIA VIA12_pin
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.035  0.035  0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035  0.035  0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.035  0.035  0.035 ;
END VIA12_pin

VIA CONT1 DEFAULT
        RESISTANCE 44.0000000000 ;
	LAYER PO ;
		RECT -0.04 -0.05 0.04 0.05 ;
	LAYER CO ;
		RECT -0.03 -0.03 0.03 0.03 ;
	LAYER M1 ;
		RECT -0.06 -0.035 0.06 0.035 ;
END CONT1

VIA VIA9AP_1cutA DEFAULT
        RESISTANCE 0.0640000000 ;
	LAYER M9 ;
		RECT -2.0 -2.0 2.0 2.0 ;
	LAYER RV ;
		RECT -1.5 -1.5 1.5 1.5 ;
	LAYER AP ;
		RECT -2.0 -2.0 2.0 2.0 ;
END VIA9AP_1cutA

VIA VIA12_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA12_1cut

VIA VIA12_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.035 0.085 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.085 0.035 0.085 ;
END VIA12_1cut_FAT_C

VIA VIA12_1cut_FAT_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.085 0.035 0.085 ;
END VIA12_1cut_FAT_V

VIA VIA12_1cut_FAT_VN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.105 ;
	LAYER VIA1 ;
		RECT -0.035 -0.015 0.035 0.055 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.105 ;
END VIA12_1cut_FAT_VN

VIA VIA12_1cut_FAT_VS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.105 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.055 0.035 0.015 ;
	LAYER M2 ;
		RECT -0.035 -0.105 0.035 0.065 ;
END VIA12_1cut_FAT_VS

VIA VIA12_1cut_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA12_1cut_H

VIA VIA12_1cut_R90 DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA12_1cut_R90

VIA VIA12_1cut_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA12_1cut_V

VIA VIA12_2cut_p1_CV DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.135 0.035 0.135 ;
	LAYER VIA1 ;
		RECT -0.035 -0.105 0.035 -0.035 ;
		RECT -0.035 0.035 0.035 0.105 ;
	LAYER M2 ;
		RECT -0.065 -0.105 0.065 0.105 ;
END VIA12_2cut_p1_CV

VIA VIA12_2cut_p1_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.065 -0.035 0.205 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.175 0.065 ;
END VIA12_2cut_p1_E

VIA VIA12_2cut_p1_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.205 -0.035 0.065 0.035 ;
	LAYER VIA1 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.175 -0.065 0.035 0.065 ;
END VIA12_2cut_p1_W

VIA VIA12_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.135 0.035 0.135 ;
	LAYER VIA1 ;
		RECT -0.035 -0.105 0.035 -0.035 ;
		RECT -0.035 0.035 0.035 0.105 ;
	LAYER M2 ;
		RECT -0.035 -0.26 0.035 0.26 ;
END VIA12_2cut_p2_BLC

VIA VIA12_2cut_p2_BLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M2 ;
		RECT -0.035 -0.19 0.035 0.33 ;
END VIA12_2cut_p2_BLN

VIA VIA12_2cut_p2_BLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.33 0.035 0.19 ;
END VIA12_2cut_p2_BLS

VIA VIA12_2cut_p2_SLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M2 ;
		RECT -0.035 -0.085 0.035 0.435 ;
END VIA12_2cut_p2_SLN

VIA VIA12_2cut_p2_SLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.435 0.035 0.085 ;
END VIA12_2cut_p2_SLS

VIA VIA12_2cut_p3_DN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.205 ;
END VIA12_2cut_p3_DN

VIA VIA12_2cut_p3_DS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.205 0.035 0.065 ;
END VIA12_2cut_p3_DS

VIA VIA12_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA1 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA12_FBD_YEN

VIA VIA12_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA1 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M2 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA12_FBD_YES

VIA VIA12_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA1 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M2 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA12_FBD_YWN

VIA VIA12_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA1 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M2 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA12_FBD_YWS

VIA VIA12_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA12_FBS

VIA VIA12_FBS_E DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.095 0.065 ;
	LAYER VIA1 ;
		RECT -0.005 -0.035 0.065 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.095 0.065 ;
END VIA12_FBS_E

VIA VIA12_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA1 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA12_FBS_EN

VIA VIA12_FBS_W DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.095 -0.065 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M2 ;
		RECT -0.095 -0.065 0.035 0.065 ;
END VIA12_FBS_W

VIA VIA12_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA1 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M2 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA12_PBD_N

VIA VIA12_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M1 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M2 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA12_PBD_S

VIA VIA12_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA12_PBS_H

VIA VIA12_PBS_HE DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.035 0.095 0.035 ;
	LAYER VIA1 ;
		RECT -0.005 -0.035 0.065 0.035 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.095 0.065 ;
END VIA12_PBS_HE

VIA VIA12_PBS_HW DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.095 -0.035 0.035 0.035 ;
	LAYER VIA1 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M2 ;
		RECT -0.095 -0.065 0.035 0.065 ;
END VIA12_PBS_HW

VIA VIA12_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M2 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA12_PBS_V

VIA VIA23_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA23_1cut

VIA VIA23_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.085 -0.035 0.085 0.035 ;
END VIA23_1cut_FAT_C

VIA VIA23_1stack_N DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.325 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA23_1stack_N

VIA VIA23_1stack_S DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.325 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA23_1stack_S

VIA VIA23_2cut_p1_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.175 ;
END VIA23_2cut_p1_N

VIA VIA23_2cut_p1_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.175 0.065 0.035 ;
END VIA23_2cut_p1_S

VIA VIA23_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.105 -0.065 0.105 0.065 ;
	LAYER VIA2 ;
		RECT -0.105 -0.035 -0.035 0.035 ;
		RECT 0.035 -0.035 0.105 0.035 ;
	LAYER M3 ;
		RECT -0.26 -0.035 0.26 0.035 ;
END VIA23_2cut_p2_BLC

VIA VIA23_2cut_p2_BLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M3 ;
		RECT -0.19 -0.035 0.33 0.035 ;
END VIA23_2cut_p2_BLE

VIA VIA23_2cut_p2_BLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.33 -0.035 0.19 0.035 ;
END VIA23_2cut_p2_BLW

VIA VIA23_2cut_p2_SLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M3 ;
		RECT -0.085 -0.035 0.435 0.035 ;
END VIA23_2cut_p2_SLE

VIA VIA23_2cut_p2_SLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.435 -0.035 0.085 0.035 ;
END VIA23_2cut_p2_SLW

VIA VIA23_2cut_p3_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.205 0.035 ;
END VIA23_2cut_p3_E

VIA VIA23_2cut_p3_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.205 -0.035 0.065 0.035 ;
END VIA23_2cut_p3_W

VIA VIA23_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA2 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA23_FBD_XEN

VIA VIA23_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA2 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M3 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA23_FBD_XES

VIA VIA23_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA2 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M3 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA23_FBD_XWN

VIA VIA23_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA2 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M3 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA23_FBD_XWS

VIA VIA23_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA2 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA23_FBD_YEN

VIA VIA23_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA2 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M3 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA23_FBD_YES

VIA VIA23_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA2 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M3 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA23_FBD_YWN

VIA VIA23_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA2 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M3 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA23_FBD_YWS

VIA VIA23_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA23_FBS

VIA VIA23_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA2 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA23_FBS_EN

VIA VIA23_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA2 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M3 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA23_FBS_ES

VIA VIA23_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA2 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M3 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA23_FBS_WN

VIA VIA23_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA2 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M3 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA23_FBS_WS

VIA VIA23_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA2 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M3 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA23_PBD_E

VIA VIA23_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA2 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA23_PBD_N

VIA VIA23_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA2 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M3 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA23_PBD_S

VIA VIA23_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M2 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA2 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M3 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA23_PBD_W

VIA VIA23_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA23_PBS_H

VIA VIA23_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M3 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA23_PBS_V

VIA VIA34_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA34_1cut

VIA VIA34_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.035 0.085 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.085 0.035 0.085 ;
END VIA34_1cut_FAT_C

VIA VIA34_1stack_E DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.325 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA34_1stack_E

VIA VIA34_1stack_W DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.325 -0.035 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA34_1stack_W

VIA VIA34_2cut_p1_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.205 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.175 0.065 ;
END VIA34_2cut_p1_E

VIA VIA34_2cut_p1_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.205 -0.035 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.175 -0.065 0.035 0.065 ;
END VIA34_2cut_p1_W

VIA VIA34_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.105 0.065 0.105 ;
	LAYER VIA3 ;
		RECT -0.035 -0.105 0.035 -0.035 ;
		RECT -0.035 0.035 0.035 0.105 ;
	LAYER M4 ;
		RECT -0.035 -0.26 0.035 0.26 ;
END VIA34_2cut_p2_BLC

VIA VIA34_2cut_p2_BLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M4 ;
		RECT -0.035 -0.19 0.035 0.33 ;
END VIA34_2cut_p2_BLN

VIA VIA34_2cut_p2_BLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.33 0.035 0.19 ;
END VIA34_2cut_p2_BLS

VIA VIA34_2cut_p2_SLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M4 ;
		RECT -0.035 -0.085 0.035 0.435 ;
END VIA34_2cut_p2_SLN

VIA VIA34_2cut_p2_SLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.435 0.035 0.085 ;
END VIA34_2cut_p2_SLS

VIA VIA34_2cut_p3_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.205 ;
END VIA34_2cut_p3_N

VIA VIA34_2cut_p3_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.205 0.035 0.065 ;
END VIA34_2cut_p3_S

VIA VIA34_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA3 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA34_FBD_XEN

VIA VIA34_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA3 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M4 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA34_FBD_XES

VIA VIA34_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA3 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M4 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA34_FBD_XWN

VIA VIA34_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA3 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M4 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA34_FBD_XWS

VIA VIA34_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA3 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA34_FBD_YEN

VIA VIA34_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA3 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M4 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA34_FBD_YES

VIA VIA34_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA3 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M4 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA34_FBD_YWN

VIA VIA34_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA3 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M4 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA34_FBD_YWS

VIA VIA34_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA34_FBS

VIA VIA34_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA3 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA34_FBS_EN

VIA VIA34_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA3 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M4 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA34_FBS_ES

VIA VIA34_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA3 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M4 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA34_FBS_WN

VIA VIA34_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA3 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M4 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA34_FBS_WS

VIA VIA34_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA3 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA34_PBD_E

VIA VIA34_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA3 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M4 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA34_PBD_N

VIA VIA34_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M4 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA34_PBD_S

VIA VIA34_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M3 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA3 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M4 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA34_PBD_W

VIA VIA34_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA34_PBS_H

VIA VIA34_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M4 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA34_PBS_V

VIA VIA45_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA45_1cut

VIA VIA45_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.085 -0.035 0.085 0.035 ;
END VIA45_1cut_FAT_C

VIA VIA45_1stack_N DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.325 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA45_1stack_N

VIA VIA45_1stack_S DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.325 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA45_1stack_S

VIA VIA45_2cut_p1_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.175 ;
END VIA45_2cut_p1_N

VIA VIA45_2cut_p1_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.175 0.065 0.035 ;
END VIA45_2cut_p1_S

VIA VIA45_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.105 -0.065 0.105 0.065 ;
	LAYER VIA4 ;
		RECT -0.105 -0.035 -0.035 0.035 ;
		RECT 0.035 -0.035 0.105 0.035 ;
	LAYER M5 ;
		RECT -0.26 -0.035 0.26 0.035 ;
END VIA45_2cut_p2_BLC

VIA VIA45_2cut_p2_BLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M5 ;
		RECT -0.19 -0.035 0.33 0.035 ;
END VIA45_2cut_p2_BLE

VIA VIA45_2cut_p2_BLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.33 -0.035 0.19 0.035 ;
END VIA45_2cut_p2_BLW

VIA VIA45_2cut_p2_SLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M5 ;
		RECT -0.085 -0.035 0.435 0.035 ;
END VIA45_2cut_p2_SLE

VIA VIA45_2cut_p2_SLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.435 -0.035 0.085 0.035 ;
END VIA45_2cut_p2_SLW

VIA VIA45_2cut_p3_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.205 0.035 ;
END VIA45_2cut_p3_E

VIA VIA45_2cut_p3_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.205 -0.035 0.065 0.035 ;
END VIA45_2cut_p3_W

VIA VIA45_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA4 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA45_FBD_XEN

VIA VIA45_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA4 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M5 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA45_FBD_XES

VIA VIA45_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA4 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M5 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA45_FBD_XWN

VIA VIA45_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA4 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M5 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA45_FBD_XWS

VIA VIA45_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA4 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA45_FBD_YEN

VIA VIA45_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA4 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M5 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA45_FBD_YES

VIA VIA45_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA4 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M5 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA45_FBD_YWN

VIA VIA45_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA4 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M5 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA45_FBD_YWS

VIA VIA45_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA45_FBS

VIA VIA45_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA4 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA45_FBS_EN

VIA VIA45_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA4 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M5 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA45_FBS_ES

VIA VIA45_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA4 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M5 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA45_FBS_WN

VIA VIA45_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA4 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M5 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA45_FBS_WS

VIA VIA45_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA4 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M5 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA45_PBD_E

VIA VIA45_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA4 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA45_PBD_N

VIA VIA45_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA4 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M5 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA45_PBD_S

VIA VIA45_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M4 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA4 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M5 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA45_PBD_W

VIA VIA45_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA45_PBS_H

VIA VIA45_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M5 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA45_PBS_V

VIA VIA56_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA56_1cut

VIA VIA56_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.035 0.085 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.085 0.035 0.085 ;
END VIA56_1cut_FAT_C

VIA VIA56_1stack_E DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.325 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA56_1stack_E

VIA VIA56_1stack_W DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.325 -0.035 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.065 ;
END VIA56_1stack_W

VIA VIA56_2cut_p1_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.205 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.175 0.065 ;
END VIA56_2cut_p1_E

VIA VIA56_2cut_p1_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.205 -0.035 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.175 -0.065 0.035 0.065 ;
END VIA56_2cut_p1_W

VIA VIA56_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.105 0.065 0.105 ;
	LAYER VIA5 ;
		RECT -0.035 -0.105 0.035 -0.035 ;
		RECT -0.035 0.035 0.035 0.105 ;
	LAYER M6 ;
		RECT -0.035 -0.26 0.035 0.26 ;
END VIA56_2cut_p2_BLC

VIA VIA56_2cut_p2_BLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M6 ;
		RECT -0.035 -0.19 0.035 0.33 ;
END VIA56_2cut_p2_BLN

VIA VIA56_2cut_p2_BLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.33 0.035 0.19 ;
END VIA56_2cut_p2_BLS

VIA VIA56_2cut_p2_SLN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M6 ;
		RECT -0.035 -0.085 0.035 0.435 ;
END VIA56_2cut_p2_SLN

VIA VIA56_2cut_p2_SLS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.435 0.035 0.085 ;
END VIA56_2cut_p2_SLS

VIA VIA56_2cut_p3_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.175 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.205 ;
END VIA56_2cut_p3_N

VIA VIA56_2cut_p3_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.065 -0.175 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.205 0.035 0.065 ;
END VIA56_2cut_p3_S

VIA VIA56_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA5 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA56_FBD_XEN

VIA VIA56_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA5 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M6 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA56_FBD_XES

VIA VIA56_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA5 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M6 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA56_FBD_XWN

VIA VIA56_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA5 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M6 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA56_FBD_XWS

VIA VIA56_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA5 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA56_FBD_YEN

VIA VIA56_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA5 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M6 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA56_FBD_YES

VIA VIA56_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA5 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M6 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA56_FBD_YWN

VIA VIA56_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA5 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M6 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA56_FBD_YWS

VIA VIA56_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA56_FBS

VIA VIA56_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA5 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA56_FBS_EN

VIA VIA56_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA5 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M6 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA56_FBS_ES

VIA VIA56_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA5 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M6 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA56_FBS_WN

VIA VIA56_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA5 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M6 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA56_FBS_WS

VIA VIA56_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA5 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA56_PBD_E

VIA VIA56_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA5 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M6 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA56_PBD_N

VIA VIA56_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M6 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA56_PBD_S

VIA VIA56_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M5 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA5 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M6 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA56_PBD_W

VIA VIA56_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA56_PBS_H

VIA VIA56_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M6 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA56_PBS_V

VIA VIA67_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA67_1cut

VIA VIA67_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.085 -0.035 0.085 0.035 ;
END VIA67_1cut_FAT_C

VIA VIA67_1stack_N DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.325 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA67_1stack_N

VIA VIA67_1stack_S DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.325 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA67_1stack_S

VIA VIA67_2cut_p1_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.175 ;
END VIA67_2cut_p1_N

VIA VIA67_2cut_p1_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.175 0.065 0.035 ;
END VIA67_2cut_p1_S

VIA VIA67_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.105 -0.065 0.105 0.065 ;
	LAYER VIA6 ;
		RECT -0.105 -0.035 -0.035 0.035 ;
		RECT 0.035 -0.035 0.105 0.035 ;
	LAYER M7 ;
		RECT -0.26 -0.035 0.26 0.035 ;
END VIA67_2cut_p2_BLC

VIA VIA67_2cut_p2_BLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M7 ;
		RECT -0.19 -0.035 0.33 0.035 ;
END VIA67_2cut_p2_BLE

VIA VIA67_2cut_p2_BLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.33 -0.035 0.19 0.035 ;
END VIA67_2cut_p2_BLW

VIA VIA67_2cut_p2_SLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M7 ;
		RECT -0.085 -0.035 0.435 0.035 ;
END VIA67_2cut_p2_SLE

VIA VIA67_2cut_p2_SLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.435 -0.035 0.085 0.035 ;
END VIA67_2cut_p2_SLW

VIA VIA67_2cut_p3_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.205 0.035 ;
END VIA67_2cut_p3_E

VIA VIA67_2cut_p3_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.205 -0.035 0.065 0.035 ;
END VIA67_2cut_p3_W

VIA VIA67_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA6 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA67_FBD_XEN

VIA VIA67_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA6 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M7 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA67_FBD_XES

VIA VIA67_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA6 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M7 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA67_FBD_XWN

VIA VIA67_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA6 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M7 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA67_FBD_XWS

VIA VIA67_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA6 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA67_FBD_YEN

VIA VIA67_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA6 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M7 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA67_FBD_YES

VIA VIA67_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA6 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M7 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA67_FBD_YWN

VIA VIA67_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA6 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M7 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA67_FBD_YWS

VIA VIA67_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA67_FBS

VIA VIA67_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA6 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA67_FBS_EN

VIA VIA67_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA6 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M7 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA67_FBS_ES

VIA VIA67_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA6 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M7 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA67_FBS_WN

VIA VIA67_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA6 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M7 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA67_FBS_WS

VIA VIA67_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA6 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA67_PBD_E

VIA VIA67_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA6 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA67_PBD_N

VIA VIA67_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA6 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M7 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA67_PBD_S

VIA VIA67_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M6 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA6 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M7 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA67_PBD_W

VIA VIA67_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA67_PBS_H

VIA VIA67_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M6 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M7 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA67_PBS_V

# Begin added by Michael Oduoza
VIA VIA78_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA78_1cut

VIA VIA78_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.085 -0.035 0.085 0.035 ;
END VIA78_1cut_FAT_C

VIA VIA78_1stack_N DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.035 0.325 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA78_1stack_N

VIA VIA78_1stack_S DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.325 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA78_1stack_S

VIA VIA78_2cut_p1_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.175 ;
END VIA78_2cut_p1_N

VIA VIA78_2cut_p1_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.175 0.065 0.035 ;
END VIA78_2cut_p1_S

VIA VIA78_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.105 -0.065 0.105 0.065 ;
	LAYER VIA7 ;
		RECT -0.105 -0.035 -0.035 0.035 ;
		RECT 0.035 -0.035 0.105 0.035 ;
	LAYER M8 ;
		RECT -0.26 -0.035 0.26 0.035 ;
END VIA78_2cut_p2_BLC

VIA VIA78_2cut_p2_BLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M8 ;
		RECT -0.19 -0.035 0.33 0.035 ;
END VIA78_2cut_p2_BLE

VIA VIA78_2cut_p2_BLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.33 -0.035 0.19 0.035 ;
END VIA78_2cut_p2_BLW

VIA VIA78_2cut_p2_SLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M8 ;
		RECT -0.085 -0.035 0.435 0.035 ;
END VIA78_2cut_p2_SLE

VIA VIA78_2cut_p2_SLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.435 -0.035 0.085 0.035 ;
END VIA78_2cut_p2_SLW

VIA VIA78_2cut_p3_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.205 0.035 ;
END VIA78_2cut_p3_E

VIA VIA78_2cut_p3_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.205 -0.035 0.065 0.035 ;
END VIA78_2cut_p3_W

VIA VIA78_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA7 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA78_FBD_XEN

VIA VIA78_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA7 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M8 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA78_FBD_XES

VIA VIA78_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA7 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M8 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA78_FBD_XWN

VIA VIA78_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA7 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M8 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA78_FBD_XWS

VIA VIA78_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA7 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA78_FBD_YEN

VIA VIA78_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA7 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M8 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA78_FBD_YES

VIA VIA78_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA7 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M8 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA78_FBD_YWN

VIA VIA78_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA7 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M8 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA78_FBD_YWS

VIA VIA78_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA78_FBS

VIA VIA78_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA7 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA78_FBS_EN

VIA VIA78_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA7 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M8 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA78_FBS_ES

VIA VIA78_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA7 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M8 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA78_FBS_WN

VIA VIA78_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA7 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M8 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA78_FBS_WS

VIA VIA78_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA7 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA78_PBD_E

VIA VIA78_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA7 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA78_PBD_N

VIA VIA78_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA7 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M8 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA78_PBD_S

VIA VIA78_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M7 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA7 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M8 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA78_PBD_W

VIA VIA78_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA78_PBS_H

VIA VIA78_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M7 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M8 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA78_PBS_V

VIA VIA89_1cut DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA89_1cut

VIA VIA89_1cut_FAT_C DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.085 0.035 0.085 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.085 -0.035 0.085 0.035 ;
END VIA89_1cut_FAT_C

VIA VIA89_1stack_N DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.035 0.325 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA89_1stack_N

VIA VIA89_1stack_S DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.325 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.065 0.035 ;
END VIA89_1stack_S

VIA VIA89_2cut_p1_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.035 0.205 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT -0.035 0.105 0.035 0.175 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.065 0.175 ;
END VIA89_2cut_p1_N

VIA VIA89_2cut_p1_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.205 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.175 0.035 -0.105 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.175 0.065 0.035 ;
END VIA89_2cut_p1_S

VIA VIA89_2cut_p2_BLC DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.105 -0.065 0.105 0.065 ;
	LAYER VIA8 ;
		RECT -0.105 -0.035 -0.035 0.035 ;
		RECT 0.035 -0.035 0.105 0.035 ;
	LAYER M9 ;
		RECT -0.26 -0.035 0.26 0.035 ;
END VIA89_2cut_p2_BLC

VIA VIA89_2cut_p2_BLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M9 ;
		RECT -0.19 -0.035 0.33 0.035 ;
END VIA89_2cut_p2_BLE

VIA VIA89_2cut_p2_BLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.33 -0.035 0.19 0.035 ;
END VIA89_2cut_p2_BLW

VIA VIA89_2cut_p2_SLE DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M9 ;
		RECT -0.085 -0.035 0.435 0.035 ;
END VIA89_2cut_p2_SLE

VIA VIA89_2cut_p2_SLW DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.435 -0.035 0.085 0.035 ;
END VIA89_2cut_p2_SLW

VIA VIA89_2cut_p3_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.175 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		RECT 0.105 -0.035 0.175 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.205 0.035 ;
END VIA89_2cut_p3_E

VIA VIA89_2cut_p3_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.175 -0.065 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.175 -0.035 -0.105 0.035 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.205 -0.035 0.065 0.035 ;
END VIA89_2cut_p3_W

VIA VIA89_FBD_XEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.235 0.095 ;
	LAYER VIA8 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT 0.135 -0.005 0.205 0.065 ;
	LAYER M9 ;
		RECT -0.035 -0.035 0.235 0.095 ;
END VIA89_FBD_XEN

VIA VIA89_FBD_XES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.095 0.235 0.035 ;
	LAYER VIA8 ;
		RECT -0.005 -0.065 0.065 0.005 ;
		RECT 0.135 -0.065 0.205 0.005 ;
	LAYER M9 ;
		RECT -0.035 -0.095 0.235 0.035 ;
END VIA89_FBD_XES

VIA VIA89_FBD_XWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.235 -0.035 0.035 0.095 ;
	LAYER VIA8 ;
		RECT -0.205 -0.005 -0.135 0.065 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M9 ;
		RECT -0.235 -0.035 0.035 0.095 ;
END VIA89_FBD_XWN

VIA VIA89_FBD_XWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.235 -0.095 0.035 0.035 ;
	LAYER VIA8 ;
		RECT -0.205 -0.065 -0.135 0.005 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M9 ;
		RECT -0.235 -0.095 0.035 0.035 ;
END VIA89_FBD_XWS

VIA VIA89_FBD_YEN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.095 0.235 ;
	LAYER VIA8 ;
		RECT -0.005 -0.005 0.065 0.065 ;
		RECT -0.005 0.135 0.065 0.205 ;
	LAYER M9 ;
		RECT -0.035 -0.035 0.095 0.235 ;
END VIA89_FBD_YEN

VIA VIA89_FBD_YES DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.235 0.095 0.035 ;
	LAYER VIA8 ;
		RECT -0.005 -0.205 0.065 -0.135 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M9 ;
		RECT -0.035 -0.235 0.095 0.035 ;
END VIA89_FBD_YES

VIA VIA89_FBD_YWN DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.095 -0.035 0.035 0.235 ;
	LAYER VIA8 ;
		RECT -0.065 -0.005 0.005 0.065 ;
		RECT -0.065 0.135 0.005 0.205 ;
	LAYER M9 ;
		RECT -0.095 -0.035 0.035 0.235 ;
END VIA89_FBD_YWN

VIA VIA89_FBD_YWS DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.095 -0.235 0.035 0.035 ;
	LAYER VIA8 ;
		RECT -0.065 -0.205 0.005 -0.135 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M9 ;
		RECT -0.095 -0.235 0.035 0.035 ;
END VIA89_FBD_YWS

VIA VIA89_FBS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.065 -0.065 0.065 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA89_FBS

VIA VIA89_FBS_EN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.095 0.095 ;
	LAYER VIA8 ;
		RECT -0.005 -0.005 0.065 0.065 ;
	LAYER M9 ;
		RECT -0.035 -0.035 0.095 0.095 ;
END VIA89_FBS_EN

VIA VIA89_FBS_ES DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.095 0.095 0.035 ;
	LAYER VIA8 ;
		RECT -0.005 -0.065 0.065 0.005 ;
	LAYER M9 ;
		RECT -0.035 -0.095 0.095 0.035 ;
END VIA89_FBS_ES

VIA VIA89_FBS_WN DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.095 -0.035 0.035 0.095 ;
	LAYER VIA8 ;
		RECT -0.065 -0.005 0.005 0.065 ;
	LAYER M9 ;
		RECT -0.095 -0.035 0.035 0.095 ;
END VIA89_FBS_WN

VIA VIA89_FBS_WS DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.095 -0.095 0.035 0.035 ;
	LAYER VIA8 ;
		RECT -0.065 -0.065 0.005 0.005 ;
	LAYER M9 ;
		RECT -0.095 -0.095 0.035 0.035 ;
END VIA89_FBS_WS

VIA VIA89_PBD_E DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.235 0.035 ;
	LAYER VIA8 ;
		RECT -0.005 -0.035 0.065 0.035 ;
		RECT 0.135 -0.035 0.205 0.035 ;
	LAYER M9 ;
		RECT -0.035 -0.065 0.235 0.065 ;
END VIA89_PBD_E

VIA VIA89_PBD_N DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.035 0.035 0.235 ;
	LAYER VIA8 ;
		RECT -0.035 -0.005 0.035 0.065 ;
		RECT -0.035 0.135 0.035 0.205 ;
	LAYER M9 ;
		RECT -0.065 -0.035 0.065 0.235 ;
END VIA89_PBD_N

VIA VIA89_PBD_S DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.035 -0.235 0.035 0.035 ;
	LAYER VIA8 ;
		RECT -0.035 -0.205 0.035 -0.135 ;
		RECT -0.035 -0.065 0.035 0.005 ;
	LAYER M9 ;
		RECT -0.065 -0.235 0.065 0.035 ;
END VIA89_PBD_S

VIA VIA89_PBD_W DEFAULT
        RESISTANCE 3.3500000000 ;
	LAYER M8 ;
		RECT -0.235 -0.035 0.035 0.035 ;
	LAYER VIA8 ;
		RECT -0.205 -0.035 -0.135 0.035 ;
		RECT -0.065 -0.035 0.005 0.035 ;
	LAYER M9 ;
		RECT -0.235 -0.065 0.035 0.065 ;
END VIA89_PBD_W

VIA VIA89_PBS_H DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.065 -0.035 0.065 0.035 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA89_PBS_H

VIA VIA89_PBS_V DEFAULT
        RESISTANCE 6.7000000000 ;
	LAYER M8 ;
		RECT -0.035 -0.065 0.035 0.065 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
	LAYER M9 ;
		RECT -0.065 -0.065 0.065 0.065 ;
END VIA89_PBS_V
# End added by Michael Oduoza

VIARULE VIAGEN12 GENERATE
	LAYER M1 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M2 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA1 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN12

VIARULE VIAGEN23 GENERATE
	LAYER M2 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M3 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA2 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN23

VIARULE VIAGEN34 GENERATE
	LAYER M3 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M4 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA3 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN34

VIARULE VIAGEN45 GENERATE
	LAYER M4 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M5 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA4 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN45

VIARULE VIAGEN56 GENERATE
	LAYER M5 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M6 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA5 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN56

VIARULE VIAGEN67 GENERATE
	LAYER M6 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M7 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA6 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN67

# Begin edited by Michael Oduoza
VIARULE VIAGEN78 GENERATE
	LAYER M7 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M8 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA7 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN78

VIARULE VIAGEN89 GENERATE
	LAYER M8 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER M9 ;
		ENCLOSURE 0.03 0 ;
		WIDTH 0.07 TO 4.50 ;
	LAYER VIA8 ;
		RECT -0.035 -0.035 0.035 0.035 ;
		SPACING 0.16 BY 0.16 ;
END VIAGEN89
# End edited by Michael Oduoza

VIARULE VIAGEN9AP GENERATE
	LAYER M9 ;
		ENCLOSURE 0.5 0.5 ;
		WIDTH 0.40 TO 12.0 ;
	LAYER AP ;
		ENCLOSURE 0.5 0.5 ;
		WIDTH 2.0 TO 35.0 ;
	LAYER RV ;
		RECT -1.5 -1.5 1.5 1.5 ;
		SPACING 5.0 BY 5.0 ;
END VIAGEN9AP

SITE core
	SIZE 0.140 BY 1.260 ;
	CLASS CORE ;
	SYMMETRY Y ;
END core

SITE bcore
	SIZE 0.140 BY 2.520 ;
	CLASS CORE ;
	SYMMETRY Y ;
END bcore

SITE bcoreExt
	SIZE 0.140 BY 2.520 ;
    CLASS CORE ;
END bcoreExt

SITE ccore
	SIZE 0.140 BY 3.780 ;
	CLASS CORE ;
	SYMMETRY Y ;
END ccore

SITE dcore
	SIZE 0.140 BY 5.040 ;
	CLASS CORE ;
	SYMMETRY Y ;
END dcore

SITE gacore
	SIZE 0.700 BY 1.260 ;
	CLASS CORE ;
	SYMMETRY Y ;
END gacore

SITE gabcore
	SIZE 0.700 BY 2.520 ;
	CLASS CORE ;
	SYMMETRY Y ;
END gabcore

# Begin added by Michael Oduoza
SITE tentoone
	SIZE 3.78 BY 3.78 ;
	CLASS CORE ;
	SYMMETRY Y ; 
END tentoone
# End added by Michael Oduoza

MACRO AN2D0BWP
    CLASS CORE ;
    FOREIGN AN2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.695 0.185 0.735 0.305 ;
        RECT  0.695 0.920 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.410 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.580 0.135 ;
        RECT  0.000 -0.115 0.460 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.990 0.580 1.375 ;
        RECT  0.150 1.145 0.460 1.375 ;
        RECT  0.070 0.960 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.650 0.640 ;
        RECT  0.515 0.205 0.585 0.915 ;
        RECT  0.150 0.205 0.515 0.275 ;
        RECT  0.340 0.845 0.515 0.915 ;
        RECT  0.260 0.845 0.340 1.045 ;
        RECT  0.070 0.205 0.150 0.335 ;
    END
END AN2D0BWP

MACRO AN2D1BWP
    CLASS CORE ;
    FOREIGN AN2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.765 0.355 0.805 0.905 ;
        RECT  0.735 0.185 0.765 1.045 ;
        RECT  0.695 0.185 0.735 0.465 ;
        RECT  0.695 0.745 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.410 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.580 0.135 ;
        RECT  0.000 -0.115 0.460 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.990 0.580 1.375 ;
        RECT  0.150 1.145 0.460 1.375 ;
        RECT  0.070 0.960 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.650 0.640 ;
        RECT  0.515 0.205 0.585 0.915 ;
        RECT  0.150 0.205 0.515 0.275 ;
        RECT  0.340 0.845 0.515 0.915 ;
        RECT  0.260 0.845 0.340 1.050 ;
        RECT  0.070 0.205 0.150 0.325 ;
    END
END AN2D1BWP

MACRO AN2D2BWP
    CLASS CORE ;
    FOREIGN AN2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.905 ;
        RECT  0.725 0.355 0.735 0.475 ;
        RECT  0.725 0.765 0.735 0.905 ;
        RECT  0.655 0.185 0.725 0.475 ;
        RECT  0.655 0.765 0.725 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.280 ;
        RECT  0.540 -0.115 0.830 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.985 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.545 0.650 0.615 ;
        RECT  0.490 0.205 0.560 0.915 ;
        RECT  0.125 0.205 0.490 0.275 ;
        RECT  0.330 0.845 0.490 0.915 ;
        RECT  0.210 0.845 0.330 1.055 ;
        RECT  0.055 0.205 0.125 0.345 ;
    END
END AN2D2BWP

MACRO AN2D4BWP
    CLASS CORE ;
    FOREIGN AN2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.485 ;
        RECT  1.375 0.700 1.445 1.030 ;
        RECT  1.295 0.355 1.375 0.485 ;
        RECT  1.295 0.700 1.375 0.820 ;
        RECT  1.085 0.355 1.295 0.820 ;
        RECT  1.015 0.185 1.085 0.475 ;
        RECT  1.015 0.700 1.085 1.030 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.740 0.640 ;
        RECT  0.595 0.520 0.665 0.790 ;
        RECT  0.245 0.720 0.595 0.790 ;
        RECT  0.170 0.495 0.245 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.355 0.525 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.475 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.280 ;
        RECT  0.900 -0.115 1.170 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.130 -0.115 0.780 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.675 1.630 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.890 1.290 1.375 ;
        RECT  0.880 1.145 1.170 1.375 ;
        RECT  0.800 1.000 0.880 1.375 ;
        RECT  0.490 1.145 0.800 1.375 ;
        RECT  0.410 1.000 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.485 ;
        RECT  1.375 0.700 1.445 1.030 ;
        RECT  1.365 0.355 1.375 0.485 ;
        RECT  1.365 0.700 1.375 0.820 ;
        RECT  0.885 0.545 0.995 0.615 ;
        RECT  0.815 0.205 0.885 0.930 ;
        RECT  0.390 0.205 0.815 0.275 ;
        RECT  0.690 0.860 0.815 0.930 ;
        RECT  0.570 0.860 0.690 1.065 ;
        RECT  0.330 0.860 0.570 0.930 ;
        RECT  0.210 0.860 0.330 1.065 ;
    END
END AN2D4BWP

MACRO AN2D8BWP
    CLASS CORE ;
    FOREIGN AN2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.185 2.570 0.445 ;
        RECT  2.490 0.700 2.570 0.990 ;
        RECT  2.190 0.325 2.490 0.445 ;
        RECT  2.190 0.700 2.490 0.820 ;
        RECT  2.110 0.185 2.190 0.445 ;
        RECT  2.110 0.700 2.190 0.990 ;
        RECT  1.995 0.325 2.110 0.445 ;
        RECT  1.995 0.700 2.110 0.820 ;
        RECT  1.810 0.325 1.995 0.820 ;
        RECT  1.785 0.185 1.810 1.045 ;
        RECT  1.715 0.185 1.785 0.445 ;
        RECT  1.715 0.700 1.785 1.045 ;
        RECT  1.430 0.325 1.715 0.445 ;
        RECT  1.430 0.700 1.715 0.820 ;
        RECT  1.350 0.185 1.430 0.445 ;
        RECT  1.350 0.700 1.430 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.110 0.770 ;
        RECT  0.535 0.700 1.015 0.770 ;
        RECT  0.445 0.495 0.535 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.545 0.875 0.625 ;
        RECT  0.730 0.350 0.805 0.625 ;
        RECT  0.265 0.350 0.730 0.420 ;
        RECT  0.195 0.350 0.265 0.640 ;
        RECT  0.125 0.495 0.195 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.445 ;
        RECT  2.400 -0.115 2.670 0.115 ;
        RECT  2.280 -0.115 2.400 0.255 ;
        RECT  2.020 -0.115 2.280 0.115 ;
        RECT  1.900 -0.115 2.020 0.255 ;
        RECT  1.640 -0.115 1.900 0.115 ;
        RECT  1.520 -0.115 1.640 0.255 ;
        RECT  1.240 -0.115 1.520 0.115 ;
        RECT  1.160 -0.115 1.240 0.265 ;
        RECT  0.520 -0.115 1.160 0.115 ;
        RECT  0.400 -0.115 0.520 0.140 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.685 2.750 1.375 ;
        RECT  2.400 1.145 2.670 1.375 ;
        RECT  2.280 0.890 2.400 1.375 ;
        RECT  2.020 1.145 2.280 1.375 ;
        RECT  1.900 0.890 2.020 1.375 ;
        RECT  1.640 1.145 1.900 1.375 ;
        RECT  1.520 0.890 1.640 1.375 ;
        RECT  1.240 1.145 1.520 1.375 ;
        RECT  1.160 0.980 1.240 1.375 ;
        RECT  0.870 1.145 1.160 1.375 ;
        RECT  0.790 0.980 0.870 1.375 ;
        RECT  0.500 1.145 0.790 1.375 ;
        RECT  0.420 0.980 0.500 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.185 2.570 0.445 ;
        RECT  2.490 0.700 2.570 0.990 ;
        RECT  2.190 0.325 2.490 0.445 ;
        RECT  2.190 0.700 2.490 0.820 ;
        RECT  2.110 0.185 2.190 0.445 ;
        RECT  2.110 0.700 2.190 0.990 ;
        RECT  2.065 0.325 2.110 0.445 ;
        RECT  2.065 0.700 2.110 0.820 ;
        RECT  1.430 0.325 1.715 0.445 ;
        RECT  1.430 0.700 1.715 0.820 ;
        RECT  1.350 0.185 1.430 0.445 ;
        RECT  1.350 0.700 1.430 0.990 ;
        RECT  2.085 0.545 2.585 0.615 ;
        RECT  1.260 0.545 1.695 0.615 ;
        RECT  1.190 0.345 1.260 0.910 ;
        RECT  1.045 0.345 1.190 0.415 ;
        RECT  1.070 0.840 1.190 0.910 ;
        RECT  0.590 0.840 0.710 1.050 ;
        RECT  0.305 0.840 0.590 0.910 ;
        RECT  0.235 0.735 0.305 1.035 ;
        RECT  0.055 0.210 0.125 0.380 ;
        RECT  0.950 0.840 1.070 1.050 ;
        RECT  0.975 0.210 1.045 0.415 ;
        RECT  0.125 0.210 0.975 0.280 ;
        RECT  0.710 0.840 0.950 0.910 ;
    END
END AN2D8BWP

MACRO AN2XD1BWP
    CLASS CORE ;
    FOREIGN AN2XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.700 0.185 0.735 0.465 ;
        RECT  0.700 0.735 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.580 0.135 ;
        RECT  0.000 -0.115 0.460 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 1.005 0.580 1.375 ;
        RECT  0.145 1.145 0.460 1.375 ;
        RECT  0.075 0.850 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.610 0.520 0.650 0.640 ;
        RECT  0.540 0.205 0.610 0.915 ;
        RECT  0.145 0.205 0.540 0.275 ;
        RECT  0.360 0.845 0.540 0.915 ;
        RECT  0.240 0.845 0.360 1.055 ;
        RECT  0.075 0.205 0.145 0.325 ;
    END
END AN2XD1BWP

MACRO AN3D0BWP
    CLASS CORE ;
    FOREIGN AN3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.045 ;
        RECT  0.840 0.190 0.875 0.320 ;
        RECT  0.840 0.920 0.875 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.000 -0.115 0.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 0.990 0.720 1.375 ;
        RECT  0.330 1.145 0.600 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.695 0.205 0.765 0.915 ;
        RECT  0.125 0.205 0.695 0.275 ;
        RECT  0.485 0.845 0.695 0.915 ;
        RECT  0.415 0.845 0.485 1.050 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.205 0.125 0.335 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END AN3D0BWP

MACRO AN3D1BWP
    CLASS CORE ;
    FOREIGN AN3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.045 ;
        RECT  0.840 0.190 0.875 0.480 ;
        RECT  0.840 0.735 0.875 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.000 -0.115 0.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 0.990 0.720 1.375 ;
        RECT  0.330 1.145 0.600 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.695 0.205 0.765 0.915 ;
        RECT  0.130 0.205 0.695 0.275 ;
        RECT  0.490 0.845 0.695 0.915 ;
        RECT  0.410 0.845 0.490 1.035 ;
        RECT  0.130 0.845 0.410 0.915 ;
        RECT  0.050 0.205 0.130 0.325 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END AN3D1BWP

MACRO AN3D2BWP
    CLASS CORE ;
    FOREIGN AN3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.905 ;
        RECT  0.805 0.185 0.875 0.470 ;
        RECT  0.805 0.765 0.875 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.115 1.120 0.115 ;
        RECT  0.990 -0.115 1.070 0.300 ;
        RECT  0.700 -0.115 0.990 0.115 ;
        RECT  0.580 -0.115 0.700 0.135 ;
        RECT  0.000 -0.115 0.580 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.960 1.070 1.375 ;
        RECT  0.700 1.145 0.990 1.375 ;
        RECT  0.580 0.985 0.700 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.725 0.545 0.795 0.615 ;
        RECT  0.655 0.205 0.725 0.915 ;
        RECT  0.130 0.205 0.655 0.275 ;
        RECT  0.485 0.845 0.655 0.915 ;
        RECT  0.415 0.845 0.485 1.075 ;
        RECT  0.130 0.845 0.415 0.915 ;
        RECT  0.050 0.205 0.130 0.325 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END AN3D2BWP

MACRO AN3D4BWP
    CLASS CORE ;
    FOREIGN AN3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.485 ;
        RECT  1.785 0.785 1.855 1.065 ;
        RECT  1.715 0.355 1.785 0.485 ;
        RECT  1.715 0.785 1.785 0.905 ;
        RECT  1.505 0.355 1.715 0.905 ;
        RECT  1.465 0.355 1.505 0.485 ;
        RECT  1.465 0.785 1.505 0.905 ;
        RECT  1.395 0.185 1.465 0.485 ;
        RECT  1.395 0.785 1.465 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.495 1.125 0.790 ;
        RECT  0.250 0.720 1.055 0.790 ;
        RECT  0.170 0.495 0.250 0.790 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.350 0.950 0.640 ;
        RECT  0.410 0.350 0.875 0.420 ;
        RECT  0.340 0.350 0.410 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.475 ;
        RECT  1.680 -0.115 1.970 0.115 ;
        RECT  1.560 -0.115 1.680 0.275 ;
        RECT  1.260 -0.115 1.560 0.115 ;
        RECT  1.180 -0.115 1.260 0.265 ;
        RECT  0.125 -0.115 1.180 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.675 2.050 1.375 ;
        RECT  1.680 1.145 1.970 1.375 ;
        RECT  1.560 0.985 1.680 1.375 ;
        RECT  1.260 1.145 1.560 1.375 ;
        RECT  1.180 1.000 1.260 1.375 ;
        RECT  0.870 1.145 1.180 1.375 ;
        RECT  0.790 1.000 0.870 1.375 ;
        RECT  0.490 1.145 0.790 1.375 ;
        RECT  0.410 1.000 0.490 1.375 ;
        RECT  0.125 1.145 0.410 1.375 ;
        RECT  0.055 0.920 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.485 ;
        RECT  1.785 0.785 1.855 1.065 ;
        RECT  1.395 0.185 1.435 0.485 ;
        RECT  1.395 0.785 1.435 1.065 ;
        RECT  1.245 0.345 1.315 0.930 ;
        RECT  1.095 0.345 1.245 0.415 ;
        RECT  1.070 0.860 1.245 0.930 ;
        RECT  1.025 0.210 1.095 0.415 ;
        RECT  0.950 0.860 1.070 1.070 ;
        RECT  0.580 0.210 1.025 0.280 ;
        RECT  0.700 0.860 0.950 0.930 ;
        RECT  0.580 0.860 0.700 1.070 ;
        RECT  0.330 0.860 0.580 0.930 ;
        RECT  0.210 0.860 0.330 1.070 ;
    END
END AN3D4BWP

MACRO AN3D8BWP
    CLASS CORE ;
    FOREIGN AN3D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.730 3.130 1.025 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  2.765 0.345 3.055 0.465 ;
        RECT  2.765 0.730 3.050 0.820 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.730 2.765 1.045 ;
        RECT  2.675 0.185 2.695 1.045 ;
        RECT  2.670 0.345 2.675 1.045 ;
        RECT  2.485 0.345 2.670 0.905 ;
        RECT  2.365 0.345 2.485 0.465 ;
        RECT  2.370 0.700 2.485 0.905 ;
        RECT  2.290 0.700 2.370 1.025 ;
        RECT  2.295 0.185 2.365 0.465 ;
        RECT  1.985 0.345 2.295 0.465 ;
        RECT  1.990 0.700 2.290 0.820 ;
        RECT  1.910 0.700 1.990 1.025 ;
        RECT  1.915 0.185 1.985 0.465 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.295 0.495 1.575 0.615 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.740 0.495 1.015 0.615 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.520 0.615 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.465 ;
        RECT  2.960 -0.115 3.230 0.115 ;
        RECT  2.840 -0.115 2.960 0.265 ;
        RECT  2.580 -0.115 2.840 0.115 ;
        RECT  2.460 -0.115 2.580 0.265 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.265 ;
        RECT  1.780 -0.115 2.080 0.115 ;
        RECT  1.700 -0.115 1.780 0.445 ;
        RECT  1.390 -0.115 1.700 0.115 ;
        RECT  1.310 -0.115 1.390 0.275 ;
        RECT  0.000 -0.115 1.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.675 3.310 1.375 ;
        RECT  2.960 1.145 3.230 1.375 ;
        RECT  2.840 0.890 2.960 1.375 ;
        RECT  2.580 1.145 2.840 1.375 ;
        RECT  2.460 0.985 2.580 1.375 ;
        RECT  2.200 1.145 2.460 1.375 ;
        RECT  2.080 0.890 2.200 1.375 ;
        RECT  1.780 1.145 2.080 1.375 ;
        RECT  1.700 0.985 1.780 1.375 ;
        RECT  1.390 1.145 1.700 1.375 ;
        RECT  1.310 0.985 1.390 1.375 ;
        RECT  1.030 1.145 1.310 1.375 ;
        RECT  0.950 0.985 1.030 1.375 ;
        RECT  0.670 1.145 0.950 1.375 ;
        RECT  0.590 0.985 0.670 1.375 ;
        RECT  0.310 1.145 0.590 1.375 ;
        RECT  0.230 0.985 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.730 3.130 1.025 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  2.765 0.345 3.055 0.465 ;
        RECT  2.765 0.730 3.050 0.820 ;
        RECT  2.365 0.345 2.415 0.465 ;
        RECT  2.370 0.700 2.415 0.905 ;
        RECT  2.290 0.700 2.370 1.025 ;
        RECT  2.295 0.185 2.365 0.465 ;
        RECT  1.985 0.345 2.295 0.465 ;
        RECT  1.990 0.700 2.290 0.820 ;
        RECT  1.910 0.700 1.990 1.025 ;
        RECT  1.915 0.185 1.985 0.465 ;
        RECT  2.800 0.545 3.130 0.615 ;
        RECT  1.810 0.545 2.395 0.615 ;
        RECT  1.720 0.545 1.810 0.915 ;
        RECT  1.565 0.845 1.720 0.915 ;
        RECT  1.470 0.205 1.590 0.415 ;
        RECT  1.495 0.845 1.565 1.075 ;
        RECT  1.205 0.845 1.495 0.915 ;
        RECT  1.205 0.345 1.470 0.415 ;
        RECT  1.135 0.185 1.205 0.415 ;
        RECT  1.135 0.845 1.205 1.075 ;
        RECT  0.750 0.345 1.135 0.415 ;
        RECT  0.845 0.845 1.135 0.915 ;
        RECT  0.210 0.205 1.050 0.275 ;
        RECT  0.775 0.845 0.845 1.075 ;
        RECT  0.670 0.845 0.775 0.915 ;
        RECT  0.590 0.345 0.670 0.915 ;
        RECT  0.125 0.345 0.590 0.415 ;
        RECT  0.485 0.845 0.590 0.915 ;
        RECT  0.415 0.845 0.485 1.075 ;
        RECT  0.130 0.845 0.415 0.915 ;
        RECT  0.050 0.845 0.130 0.975 ;
        RECT  0.055 0.255 0.125 0.415 ;
    END
END AN3D8BWP

MACRO AN3XD1BWP
    CLASS CORE ;
    FOREIGN AN3XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.185 0.945 1.045 ;
        RECT  0.840 0.185 0.865 0.475 ;
        RECT  0.840 0.735 0.865 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.200 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.000 -0.115 0.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.145 0.980 1.375 ;
        RECT  0.620 0.985 0.700 1.375 ;
        RECT  0.310 1.145 0.620 1.375 ;
        RECT  0.230 0.985 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.695 0.205 0.765 0.915 ;
        RECT  0.125 0.205 0.695 0.275 ;
        RECT  0.510 0.845 0.695 0.915 ;
        RECT  0.390 0.845 0.510 1.055 ;
        RECT  0.125 0.845 0.390 0.915 ;
        RECT  0.055 0.205 0.125 0.325 ;
        RECT  0.055 0.845 0.125 0.975 ;
    END
END AN3XD1BWP

MACRO AN4D0BWP
    CLASS CORE ;
    FOREIGN AN4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.195 1.085 1.055 ;
        RECT  0.980 0.195 1.015 0.315 ;
        RECT  0.980 0.930 1.015 1.055 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.505 0.735 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.695 0.580 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 0.985 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.960 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.205 0.910 0.915 ;
        RECT  0.125 0.205 0.840 0.275 ;
        RECT  0.670 0.845 0.840 0.915 ;
        RECT  0.590 0.845 0.670 1.045 ;
        RECT  0.310 0.845 0.590 0.915 ;
        RECT  0.230 0.845 0.310 1.045 ;
        RECT  0.055 0.205 0.125 0.345 ;
    END
END AN4D0BWP

MACRO AN4D1BWP
    CLASS CORE ;
    FOREIGN AN4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.195 1.085 1.045 ;
        RECT  0.995 0.195 1.015 0.475 ;
        RECT  0.995 0.735 1.015 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.505 0.735 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.695 0.580 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 0.985 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.960 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.205 0.920 0.915 ;
        RECT  0.130 0.205 0.850 0.275 ;
        RECT  0.670 0.845 0.850 0.915 ;
        RECT  0.590 0.845 0.670 1.045 ;
        RECT  0.310 0.845 0.590 0.915 ;
        RECT  0.230 0.845 0.310 1.045 ;
        RECT  0.050 0.205 0.130 0.330 ;
    END
END AN4D1BWP

MACRO AN4D2BWP
    CLASS CORE ;
    FOREIGN AN4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.355 1.085 0.905 ;
        RECT  1.015 0.185 1.025 1.065 ;
        RECT  0.955 0.185 1.015 0.465 ;
        RECT  0.955 0.785 1.015 1.065 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.765 ;
        RECT  0.595 0.635 0.665 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.585 0.565 ;
        RECT  0.455 0.355 0.525 0.635 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.300 ;
        RECT  0.850 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.850 0.290 ;
        RECT  0.000 -0.115 0.770 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.960 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.985 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.985 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.960 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.885 0.520 0.910 0.640 ;
        RECT  0.815 0.370 0.885 0.915 ;
        RECT  0.700 0.370 0.815 0.440 ;
        RECT  0.690 0.845 0.815 0.915 ;
        RECT  0.630 0.205 0.700 0.440 ;
        RECT  0.570 0.845 0.690 1.055 ;
        RECT  0.130 0.205 0.630 0.275 ;
        RECT  0.330 0.845 0.570 0.915 ;
        RECT  0.210 0.845 0.330 1.055 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AN4D2BWP

MACRO AN4D4BWP
    CLASS CORE ;
    FOREIGN AN4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2098 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.485 ;
        RECT  2.275 0.745 2.285 1.025 ;
        RECT  2.215 0.185 2.275 1.025 ;
        RECT  2.065 0.355 2.215 0.905 ;
        RECT  1.925 0.355 2.065 0.485 ;
        RECT  1.915 0.745 2.065 0.905 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.845 0.745 1.915 1.025 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.520 1.580 0.915 ;
        RECT  0.410 0.845 1.505 0.915 ;
        RECT  0.315 0.740 0.410 0.915 ;
        RECT  0.245 0.740 0.315 0.810 ;
        RECT  0.165 0.495 0.245 0.810 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.345 1.370 0.765 ;
        RECT  0.410 0.345 1.290 0.415 ;
        RECT  0.315 0.345 0.410 0.655 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.520 1.160 0.765 ;
        RECT  0.665 0.695 1.090 0.765 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.275 ;
        RECT  1.720 -0.115 2.010 0.115 ;
        RECT  1.640 -0.115 1.720 0.300 ;
        RECT  0.125 -0.115 1.640 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.985 2.130 1.375 ;
        RECT  1.720 1.145 2.010 1.375 ;
        RECT  1.600 1.125 1.720 1.375 ;
        RECT  1.300 1.145 1.600 1.375 ;
        RECT  1.180 1.125 1.300 1.375 ;
        RECT  0.900 1.145 1.180 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 1.125 0.520 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.970 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.355 1.995 0.485 ;
        RECT  1.915 0.745 1.995 0.905 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.845 0.745 1.915 1.025 ;
        RECT  1.705 0.370 1.775 1.055 ;
        RECT  1.530 0.370 1.705 0.440 ;
        RECT  0.210 0.985 1.705 1.055 ;
        RECT  1.460 0.205 1.530 0.440 ;
        RECT  0.810 0.205 1.460 0.275 ;
    END
END AN4D4BWP

MACRO AN4D8BWP
    CLASS CORE ;
    FOREIGN AN4D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 0.695 3.550 0.995 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.345 3.475 0.465 ;
        RECT  3.190 0.695 3.470 0.815 ;
        RECT  3.115 0.695 3.190 0.995 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.110 0.345 3.115 0.995 ;
        RECT  2.905 0.345 3.110 0.905 ;
        RECT  2.825 0.345 2.905 0.465 ;
        RECT  2.830 0.695 2.905 0.905 ;
        RECT  2.750 0.695 2.830 0.995 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.345 2.755 0.465 ;
        RECT  2.470 0.695 2.750 0.815 ;
        RECT  2.390 0.695 2.470 0.995 ;
        RECT  2.395 0.185 2.465 0.465 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.065 0.765 ;
        RECT  1.715 0.495 1.995 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.295 0.495 1.575 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.085 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.175 0.495 0.455 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.465 ;
        RECT  3.390 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.390 0.275 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.275 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.275 ;
        RECT  2.290 -0.115 2.550 0.115 ;
        RECT  2.210 -0.115 2.290 0.455 ;
        RECT  1.930 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.930 0.275 ;
        RECT  0.000 -0.115 1.850 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.675 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 0.885 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 0.985 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 0.885 2.670 1.375 ;
        RECT  2.290 1.145 2.550 1.375 ;
        RECT  2.210 0.985 2.290 1.375 ;
        RECT  1.930 1.145 2.210 1.375 ;
        RECT  1.850 0.985 1.930 1.375 ;
        RECT  1.570 1.145 1.850 1.375 ;
        RECT  1.490 0.985 1.570 1.375 ;
        RECT  1.210 1.145 1.490 1.375 ;
        RECT  1.130 0.985 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.985 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.985 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.810 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.470 0.695 3.550 0.995 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.345 3.475 0.465 ;
        RECT  3.190 0.695 3.470 0.815 ;
        RECT  3.185 0.695 3.190 0.995 ;
        RECT  2.825 0.345 2.835 0.465 ;
        RECT  2.830 0.695 2.835 0.905 ;
        RECT  2.750 0.695 2.830 0.995 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.345 2.755 0.465 ;
        RECT  2.470 0.695 2.750 0.815 ;
        RECT  2.390 0.695 2.470 0.995 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  3.220 0.545 3.550 0.615 ;
        RECT  2.280 0.545 2.815 0.615 ;
        RECT  2.200 0.545 2.280 0.915 ;
        RECT  2.130 0.845 2.200 0.915 ;
        RECT  2.010 0.205 2.130 0.415 ;
        RECT  2.010 0.845 2.130 1.055 ;
        RECT  1.750 0.345 2.010 0.415 ;
        RECT  1.770 0.845 2.010 0.915 ;
        RECT  1.650 0.845 1.770 1.055 ;
        RECT  1.670 0.205 1.750 0.415 ;
        RECT  1.290 0.205 1.670 0.275 ;
        RECT  1.410 0.845 1.650 0.915 ;
        RECT  1.205 0.345 1.590 0.415 ;
        RECT  1.290 0.845 1.410 1.055 ;
        RECT  1.050 0.845 1.290 0.915 ;
        RECT  1.135 0.185 1.205 0.415 ;
        RECT  0.750 0.345 1.135 0.415 ;
        RECT  0.210 0.205 1.050 0.275 ;
        RECT  0.930 0.845 1.050 1.055 ;
        RECT  0.690 0.845 0.930 0.915 ;
        RECT  0.665 0.845 0.690 1.055 ;
        RECT  0.595 0.345 0.665 1.055 ;
        RECT  0.125 0.345 0.595 0.415 ;
        RECT  0.570 0.845 0.595 1.055 ;
        RECT  0.330 0.845 0.570 0.915 ;
        RECT  0.210 0.845 0.330 1.055 ;
        RECT  0.055 0.255 0.125 0.415 ;
    END
END AN4D8BWP

MACRO AN4XD1BWP
    CLASS CORE ;
    FOREIGN AN4XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.165 0.355 1.225 0.765 ;
        RECT  1.155 0.195 1.165 0.765 ;
        RECT  1.095 0.195 1.155 0.475 ;
        RECT  1.150 0.675 1.155 0.765 ;
        RECT  1.080 0.675 1.150 1.075 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.830 0.640 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.495 0.665 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.390 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 -0.115 1.260 0.115 ;
        RECT  0.840 -0.115 0.960 0.130 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.840 0.985 0.960 1.375 ;
        RECT  0.540 1.145 0.840 1.375 ;
        RECT  0.420 0.985 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.540 1.050 0.610 ;
        RECT  0.930 0.200 1.000 0.915 ;
        RECT  0.125 0.200 0.930 0.275 ;
        RECT  0.740 0.845 0.930 0.915 ;
        RECT  0.620 0.845 0.740 1.055 ;
        RECT  0.340 0.845 0.620 0.915 ;
        RECT  0.220 0.845 0.340 1.055 ;
        RECT  0.055 0.200 0.125 0.320 ;
    END
END AN4XD1BWP

MACRO ANTENNABWP
    CLASS CORE ;
    FOREIGN ANTENNABWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN I
        ANTENNADIFFAREA 0.1184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.190 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
END ANTENNABWP

MACRO AO211D0BWP
    CLASS CORE ;
    FOREIGN AO211D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.190 1.085 1.045 ;
        RECT  0.990 0.190 1.015 0.310 ;
        RECT  0.990 0.890 1.015 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.520 0.755 0.705 ;
        RECT  0.665 0.635 0.685 0.705 ;
        RECT  0.595 0.635 0.665 0.905 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.485 0.600 0.555 ;
        RECT  0.455 0.485 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.145 1.120 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 0.930 0.640 ;
        RECT  0.850 0.205 0.920 1.055 ;
        RECT  0.130 0.205 0.850 0.275 ;
        RECT  0.210 0.985 0.850 1.055 ;
        RECT  0.130 0.845 0.515 0.915 ;
        RECT  0.050 0.205 0.130 0.335 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END AO211D0BWP

MACRO AO211D1BWP
    CLASS CORE ;
    FOREIGN AO211D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.190 1.085 1.045 ;
        RECT  0.990 0.190 1.015 0.470 ;
        RECT  0.990 0.735 1.015 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.520 0.755 0.905 ;
        RECT  0.595 0.775 0.685 0.905 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.145 1.120 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 0.930 0.640 ;
        RECT  0.850 0.205 0.920 1.055 ;
        RECT  0.685 0.205 0.850 0.275 ;
        RECT  0.210 0.985 0.850 1.055 ;
        RECT  0.615 0.205 0.685 0.440 ;
        RECT  0.130 0.205 0.615 0.275 ;
        RECT  0.130 0.845 0.510 0.915 ;
        RECT  0.050 0.205 0.130 0.325 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO211D1BWP

MACRO AO211D2BWP
    CLASS CORE ;
    FOREIGN AO211D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.355 1.085 0.905 ;
        RECT  1.015 0.185 1.025 1.055 ;
        RECT  0.955 0.185 1.015 0.465 ;
        RECT  0.955 0.770 1.015 1.055 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.765 ;
        RECT  0.595 0.635 0.665 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.580 0.565 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.300 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.250 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.250 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.960 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.000 1.145 0.750 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.885 0.520 0.910 0.640 ;
        RECT  0.815 0.345 0.885 0.915 ;
        RECT  0.665 0.345 0.815 0.415 ;
        RECT  0.670 0.845 0.815 0.915 ;
        RECT  0.600 0.845 0.670 1.055 ;
        RECT  0.595 0.255 0.665 0.415 ;
        RECT  0.210 0.985 0.600 1.055 ;
        RECT  0.290 0.345 0.595 0.415 ;
        RECT  0.130 0.845 0.510 0.915 ;
        RECT  0.220 0.215 0.290 0.415 ;
        RECT  0.140 0.215 0.220 0.290 ;
        RECT  0.040 0.190 0.140 0.290 ;
        RECT  0.050 0.845 0.130 1.000 ;
    END
END AO211D2BWP

MACRO AO211D4BWP
    CLASS CORE ;
    FOREIGN AO211D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.485 ;
        RECT  2.275 0.745 2.285 1.030 ;
        RECT  2.215 0.185 2.275 1.030 ;
        RECT  2.065 0.365 2.215 0.905 ;
        RECT  1.925 0.365 2.065 0.485 ;
        RECT  1.925 0.745 2.065 0.905 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.745 1.925 1.030 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.510 0.740 0.765 ;
        RECT  0.245 0.695 0.670 0.765 ;
        RECT  0.170 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.520 1.505 0.775 ;
        RECT  0.945 0.705 1.430 0.775 ;
        RECT  0.840 0.495 0.945 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.355 1.225 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.750 -0.115 2.010 0.115 ;
        RECT  1.670 -0.115 1.750 0.300 ;
        RECT  1.570 -0.115 1.670 0.115 ;
        RECT  1.490 -0.115 1.570 0.300 ;
        RECT  0.850 -0.115 1.490 0.115 ;
        RECT  0.770 -0.115 0.850 0.265 ;
        RECT  0.490 -0.115 0.770 0.115 ;
        RECT  0.410 -0.115 0.490 0.275 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.985 2.130 1.375 ;
        RECT  1.760 1.145 2.010 1.375 ;
        RECT  1.640 1.125 1.760 1.375 ;
        RECT  0.510 1.145 1.640 1.375 ;
        RECT  0.390 1.000 0.510 1.375 ;
        RECT  0.000 1.145 0.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.365 1.995 0.485 ;
        RECT  1.925 0.745 1.995 0.905 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.745 1.925 1.030 ;
        RECT  1.710 0.370 1.780 1.055 ;
        RECT  1.390 0.370 1.710 0.440 ;
        RECT  0.930 0.985 1.710 1.055 ;
        RECT  0.845 0.845 1.590 0.915 ;
        RECT  1.320 0.205 1.390 0.440 ;
        RECT  1.025 0.205 1.320 0.275 ;
        RECT  0.955 0.205 1.025 0.415 ;
        RECT  0.690 0.345 0.955 0.415 ;
        RECT  0.775 0.845 0.845 1.075 ;
        RECT  0.130 0.845 0.775 0.915 ;
        RECT  0.570 0.205 0.690 0.415 ;
        RECT  0.330 0.345 0.570 0.415 ;
        RECT  0.210 0.205 0.330 0.415 ;
        RECT  0.050 0.845 0.130 1.010 ;
    END
END AO211D4BWP

MACRO AO21D0BWP
    CLASS CORE ;
    FOREIGN AO21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0391 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 1.045 ;
        RECT  0.855 0.195 0.875 0.315 ;
        RECT  0.855 0.920 0.875 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.130 -0.115 0.620 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 1.000 0.740 1.375 ;
        RECT  0.000 1.145 0.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.775 0.520 0.805 0.640 ;
        RECT  0.705 0.205 0.775 0.925 ;
        RECT  0.400 0.205 0.705 0.275 ;
        RECT  0.210 0.855 0.705 0.925 ;
        RECT  0.130 0.995 0.520 1.065 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO21D0BWP

MACRO AO21D1BWP
    CLASS CORE ;
    FOREIGN AO21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 1.045 ;
        RECT  0.860 0.195 0.875 0.475 ;
        RECT  0.855 0.735 0.875 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.130 -0.115 0.620 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 1.005 0.740 1.375 ;
        RECT  0.000 1.145 0.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.775 0.520 0.805 0.640 ;
        RECT  0.705 0.205 0.775 0.915 ;
        RECT  0.400 0.205 0.705 0.275 ;
        RECT  0.210 0.845 0.705 0.915 ;
        RECT  0.130 0.995 0.510 1.065 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO21D1BWP

MACRO AO21D2BWP
    CLASS CORE ;
    FOREIGN AO21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.370 0.945 0.890 ;
        RECT  0.865 0.370 0.875 0.465 ;
        RECT  0.865 0.785 0.875 0.890 ;
        RECT  0.795 0.205 0.865 0.465 ;
        RECT  0.795 0.785 0.865 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.115 1.120 0.115 ;
        RECT  0.970 -0.115 1.050 0.300 ;
        RECT  0.700 -0.115 0.970 0.115 ;
        RECT  0.580 -0.115 0.700 0.135 ;
        RECT  0.130 -0.115 0.580 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.120 1.375 ;
        RECT  0.970 0.960 1.050 1.375 ;
        RECT  0.700 1.145 0.970 1.375 ;
        RECT  0.580 1.125 0.700 1.375 ;
        RECT  0.000 1.145 0.580 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.725 0.520 0.750 0.640 ;
        RECT  0.655 0.205 0.725 1.055 ;
        RECT  0.390 0.205 0.655 0.275 ;
        RECT  0.210 0.985 0.655 1.055 ;
        RECT  0.130 0.845 0.520 0.915 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO21D2BWP

MACRO AO21D4BWP
    CLASS CORE ;
    FOREIGN AO21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 0.185 1.845 0.485 ;
        RECT  1.775 0.745 1.845 1.030 ;
        RECT  1.715 0.355 1.775 0.485 ;
        RECT  1.715 0.745 1.775 0.905 ;
        RECT  1.505 0.355 1.715 0.905 ;
        RECT  1.465 0.355 1.505 0.485 ;
        RECT  1.465 0.745 1.505 0.905 ;
        RECT  1.395 0.185 1.465 0.485 ;
        RECT  1.395 0.745 1.465 1.030 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.520 1.130 0.780 ;
        RECT  0.245 0.710 1.050 0.780 ;
        RECT  0.145 0.495 0.245 0.780 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.970 0.640 ;
        RECT  0.410 0.345 0.875 0.415 ;
        RECT  0.315 0.345 0.410 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 -0.115 2.100 0.115 ;
        RECT  1.950 -0.115 2.030 0.475 ;
        RECT  1.680 -0.115 1.950 0.115 ;
        RECT  1.560 -0.115 1.680 0.280 ;
        RECT  1.280 -0.115 1.560 0.115 ;
        RECT  1.160 -0.115 1.280 0.135 ;
        RECT  0.700 -0.115 1.160 0.115 ;
        RECT  0.580 -0.115 0.700 0.135 ;
        RECT  0.125 -0.115 0.580 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.145 2.100 1.375 ;
        RECT  1.950 0.675 2.030 1.375 ;
        RECT  1.680 1.145 1.950 1.375 ;
        RECT  1.560 0.985 1.680 1.375 ;
        RECT  1.280 1.145 1.560 1.375 ;
        RECT  1.160 0.990 1.280 1.375 ;
        RECT  0.125 1.145 1.160 1.375 ;
        RECT  0.055 0.870 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.845 0.485 ;
        RECT  1.785 0.745 1.845 1.030 ;
        RECT  1.395 0.185 1.435 0.485 ;
        RECT  1.395 0.745 1.435 1.030 ;
        RECT  1.245 0.205 1.315 0.920 ;
        RECT  0.210 0.205 1.245 0.275 ;
        RECT  0.390 0.850 1.245 0.920 ;
        RECT  0.210 0.990 1.070 1.060 ;
    END
END AO21D4BWP

MACRO AO221D0BWP
    CLASS CORE ;
    FOREIGN AO221D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.045 ;
        RECT  1.400 0.185 1.435 0.290 ;
        RECT  1.415 0.920 1.435 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.635 1.225 0.905 ;
        RECT  1.065 0.635 1.155 0.755 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.805 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.530 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.540 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.710 -0.115 1.180 0.115 ;
        RECT  0.590 -0.115 0.710 0.135 ;
        RECT  0.130 -0.115 0.590 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.200 0.985 1.280 1.375 ;
        RECT  0.000 1.145 1.200 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.640 ;
        RECT  1.065 0.355 1.295 0.425 ;
        RECT  0.990 0.845 1.070 1.045 ;
        RECT  0.995 0.205 1.065 0.425 ;
        RECT  0.340 0.205 0.995 0.275 ;
        RECT  0.590 0.845 0.990 0.915 ;
        RECT  0.505 0.985 0.910 1.055 ;
        RECT  0.435 0.875 0.505 1.055 ;
        RECT  0.125 0.985 0.435 1.055 ;
        RECT  0.270 0.205 0.340 0.915 ;
        RECT  0.210 0.845 0.270 0.915 ;
        RECT  0.055 0.875 0.125 1.055 ;
    END
END AO221D0BWP

MACRO AO221D1BWP
    CLASS CORE ;
    FOREIGN AO221D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.195 1.505 1.045 ;
        RECT  1.410 0.195 1.435 0.475 ;
        RECT  1.410 0.735 1.435 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.520 1.165 0.640 ;
        RECT  1.015 0.355 1.085 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.760 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.495 0.525 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.115 1.540 0.115 ;
        RECT  1.170 -0.115 1.290 0.135 ;
        RECT  0.700 -0.115 1.170 0.115 ;
        RECT  0.620 -0.115 0.700 0.280 ;
        RECT  0.140 -0.115 0.620 0.115 ;
        RECT  0.040 -0.115 0.140 0.290 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.145 1.540 1.375 ;
        RECT  1.190 0.740 1.270 1.375 ;
        RECT  0.000 1.145 1.190 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.265 0.205 1.340 0.640 ;
        RECT  0.875 0.205 1.265 0.275 ;
        RECT  0.985 0.845 1.055 1.030 ;
        RECT  0.600 0.845 0.985 0.915 ;
        RECT  0.125 0.995 0.900 1.065 ;
        RECT  0.805 0.205 0.875 0.420 ;
        RECT  0.340 0.350 0.805 0.420 ;
        RECT  0.270 0.350 0.340 0.915 ;
        RECT  0.210 0.845 0.270 0.915 ;
        RECT  0.055 0.905 0.125 1.065 ;
    END
END AO221D1BWP

MACRO AO221D2BWP
    CLASS CORE ;
    FOREIGN AO221D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.355 1.505 0.765 ;
        RECT  1.435 0.205 1.445 1.075 ;
        RECT  1.375 0.205 1.435 0.465 ;
        RECT  1.375 0.675 1.435 1.075 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.105 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.300 ;
        RECT  1.260 -0.115 1.550 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.670 -0.115 1.140 0.115 ;
        RECT  0.590 -0.115 0.670 0.280 ;
        RECT  0.130 -0.115 0.590 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.840 1.630 1.375 ;
        RECT  1.240 1.145 1.550 1.375 ;
        RECT  1.160 0.820 1.240 1.375 ;
        RECT  0.000 1.145 1.160 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.235 0.205 1.305 0.640 ;
        RECT  0.850 0.205 1.235 0.275 ;
        RECT  0.955 0.845 1.025 1.030 ;
        RECT  0.570 0.845 0.955 0.915 ;
        RECT  0.125 0.985 0.870 1.055 ;
        RECT  0.780 0.205 0.850 0.420 ;
        RECT  0.485 0.350 0.780 0.420 ;
        RECT  0.415 0.185 0.485 0.420 ;
        RECT  0.330 0.350 0.415 0.420 ;
        RECT  0.260 0.350 0.330 0.915 ;
        RECT  0.210 0.845 0.260 0.915 ;
        RECT  0.055 0.845 0.125 1.055 ;
    END
END AO221D2BWP

MACRO AO221D4BWP
    CLASS CORE ;
    FOREIGN AO221D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.705 0.465 ;
        RECT  2.695 0.745 2.705 1.030 ;
        RECT  2.635 0.185 2.695 1.030 ;
        RECT  2.485 0.355 2.635 0.905 ;
        RECT  2.345 0.355 2.485 0.465 ;
        RECT  2.345 0.745 2.485 0.905 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.745 2.345 1.030 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.945 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.525 0.775 ;
        RECT  1.085 0.705 1.435 0.775 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.950 0.495 1.015 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.260 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.740 0.640 ;
        RECT  0.595 0.520 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 0.355 0.525 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.475 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.280 ;
        RECT  2.165 -0.115 2.430 0.115 ;
        RECT  2.095 -0.115 2.165 0.275 ;
        RECT  1.740 -0.115 2.095 0.115 ;
        RECT  1.740 0.205 1.830 0.275 ;
        RECT  1.620 -0.115 1.740 0.275 ;
        RECT  0.900 -0.115 1.620 0.115 ;
        RECT  1.530 0.205 1.620 0.275 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.130 -0.115 0.780 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.680 2.890 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 0.985 2.550 1.375 ;
        RECT  2.170 1.145 2.430 1.375 ;
        RECT  2.090 0.695 2.170 1.375 ;
        RECT  1.810 1.145 2.090 1.375 ;
        RECT  1.730 0.985 1.810 1.375 ;
        RECT  0.000 1.145 1.730 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.465 ;
        RECT  2.345 0.745 2.415 0.905 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.745 2.345 1.030 ;
        RECT  2.205 0.545 2.395 0.615 ;
        RECT  2.135 0.345 2.205 0.615 ;
        RECT  1.985 0.345 2.135 0.415 ;
        RECT  1.915 0.185 1.985 0.415 ;
        RECT  1.915 0.845 1.985 1.035 ;
        RECT  1.440 0.345 1.915 0.415 ;
        RECT  0.990 0.845 1.915 0.915 ;
        RECT  0.130 0.985 1.650 1.055 ;
        RECT  1.370 0.205 1.440 0.415 ;
        RECT  0.880 0.205 1.370 0.275 ;
        RECT  0.810 0.205 0.880 0.915 ;
        RECT  0.390 0.205 0.810 0.275 ;
        RECT  0.210 0.845 0.810 0.915 ;
        RECT  0.050 0.875 0.130 1.055 ;
    END
END AO221D4BWP

MACRO AO222D0BWP
    CLASS CORE ;
    FOREIGN AO222D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.045 ;
        RECT  1.540 0.185 1.575 0.290 ;
        RECT  1.555 0.895 1.575 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.495 1.365 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.520 1.150 0.640 ;
        RECT  1.015 0.355 1.085 0.640 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.630 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.800 0.495 0.875 0.620 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 -0.115 1.680 0.115 ;
        RECT  1.350 -0.115 1.470 0.250 ;
        RECT  0.520 -0.115 1.350 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.145 1.680 1.375 ;
        RECT  1.370 0.895 1.450 1.375 ;
        RECT  1.090 1.145 1.370 1.375 ;
        RECT  0.990 0.990 1.090 1.375 ;
        RECT  0.000 1.145 0.990 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.515 ;
        RECT  1.260 0.355 1.435 0.425 ;
        RECT  1.190 0.845 1.270 1.020 ;
        RECT  1.190 0.205 1.260 0.425 ;
        RECT  0.720 0.205 1.190 0.275 ;
        RECT  0.315 0.845 1.190 0.915 ;
        RECT  0.130 0.985 0.910 1.055 ;
        RECT  0.650 0.205 0.720 0.765 ;
        RECT  0.125 0.205 0.650 0.275 ;
        RECT  0.600 0.695 0.650 0.765 ;
        RECT  0.245 0.765 0.315 0.915 ;
        RECT  0.050 0.935 0.130 1.055 ;
        RECT  0.055 0.205 0.125 0.325 ;
    END
END AO222D0BWP

MACRO AO222D1BWP
    CLASS CORE ;
    FOREIGN AO222D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.045 ;
        RECT  1.555 0.185 1.575 0.465 ;
        RECT  1.555 0.735 1.575 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.675 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.650 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.610 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.800 0.495 0.875 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 1.680 0.115 ;
        RECT  1.340 -0.115 1.460 0.250 ;
        RECT  0.520 -0.115 1.340 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.145 1.680 1.375 ;
        RECT  1.360 0.740 1.440 1.375 ;
        RECT  1.090 1.145 1.360 1.375 ;
        RECT  0.970 1.000 1.090 1.375 ;
        RECT  0.000 1.145 0.970 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.485 0.520 1.505 0.640 ;
        RECT  1.415 0.320 1.485 0.640 ;
        RECT  1.260 0.320 1.415 0.390 ;
        RECT  0.210 0.855 1.270 0.925 ;
        RECT  1.190 0.205 1.260 0.390 ;
        RECT  0.730 0.205 1.190 0.275 ;
        RECT  0.130 0.995 0.890 1.065 ;
        RECT  0.660 0.205 0.730 0.785 ;
        RECT  0.125 0.205 0.660 0.275 ;
        RECT  0.600 0.685 0.660 0.785 ;
        RECT  0.050 0.925 0.130 1.065 ;
        RECT  0.055 0.205 0.125 0.355 ;
    END
END AO222D1BWP

MACRO AO222D2BWP
    CLASS CORE ;
    FOREIGN AO222D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.585 0.355 1.645 0.905 ;
        RECT  1.575 0.185 1.585 1.045 ;
        RECT  1.515 0.185 1.575 0.465 ;
        RECT  1.515 0.785 1.575 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.295 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.675 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.610 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.800 0.495 0.875 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.300 ;
        RECT  1.430 -0.115 1.690 0.115 ;
        RECT  1.310 -0.115 1.430 0.250 ;
        RECT  0.520 -0.115 1.310 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.960 1.770 1.375 ;
        RECT  1.410 1.145 1.690 1.375 ;
        RECT  1.330 0.740 1.410 1.375 ;
        RECT  1.050 1.145 1.330 1.375 ;
        RECT  0.970 1.000 1.050 1.375 ;
        RECT  0.000 1.145 0.970 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.445 0.520 1.470 0.640 ;
        RECT  1.375 0.320 1.445 0.640 ;
        RECT  1.235 0.320 1.375 0.390 ;
        RECT  0.205 0.855 1.250 0.925 ;
        RECT  1.165 0.205 1.235 0.390 ;
        RECT  0.730 0.205 1.165 0.275 ;
        RECT  0.125 0.995 0.890 1.065 ;
        RECT  0.660 0.205 0.730 0.785 ;
        RECT  0.125 0.205 0.660 0.275 ;
        RECT  0.600 0.685 0.660 0.785 ;
        RECT  0.055 0.205 0.125 0.345 ;
        RECT  0.055 0.945 0.125 1.065 ;
    END
END AO222D2BWP

MACRO AO222D4BWP
    CLASS CORE ;
    FOREIGN AO222D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.485 ;
        RECT  3.115 0.710 3.125 1.045 ;
        RECT  3.055 0.185 3.115 1.045 ;
        RECT  2.905 0.355 3.055 0.830 ;
        RECT  2.765 0.355 2.905 0.485 ;
        RECT  2.765 0.710 2.905 0.830 ;
        RECT  2.695 0.185 2.765 0.485 ;
        RECT  2.695 0.710 2.765 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.520 2.420 0.640 ;
        RECT  2.275 0.520 2.345 0.775 ;
        RECT  1.810 0.705 2.275 0.775 ;
        RECT  1.715 0.495 1.810 0.775 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.105 0.355 2.205 0.630 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.495 1.645 0.775 ;
        RECT  1.085 0.705 1.550 0.775 ;
        RECT  1.015 0.520 1.085 0.775 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.255 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.640 ;
        RECT  0.595 0.520 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 0.355 0.525 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.475 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.280 ;
        RECT  2.580 -0.115 2.850 0.115 ;
        RECT  2.460 -0.115 2.580 0.135 ;
        RECT  1.740 -0.115 2.460 0.115 ;
        RECT  1.740 0.205 1.840 0.275 ;
        RECT  1.620 -0.115 1.740 0.275 ;
        RECT  0.900 -0.115 1.620 0.115 ;
        RECT  1.520 0.205 1.620 0.275 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.130 -0.115 0.780 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.680 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.900 2.970 1.375 ;
        RECT  2.560 1.145 2.850 1.375 ;
        RECT  2.480 0.750 2.560 1.375 ;
        RECT  2.170 1.145 2.480 1.375 ;
        RECT  2.090 0.985 2.170 1.375 ;
        RECT  1.810 1.145 2.090 1.375 ;
        RECT  1.730 0.985 1.810 1.375 ;
        RECT  0.000 1.145 1.730 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.485 ;
        RECT  2.765 0.710 2.835 0.830 ;
        RECT  2.695 0.185 2.765 0.485 ;
        RECT  2.695 0.710 2.765 1.045 ;
        RECT  2.545 0.205 2.615 0.640 ;
        RECT  2.025 0.205 2.545 0.275 ;
        RECT  2.250 0.845 2.370 1.055 ;
        RECT  2.010 0.845 2.250 0.915 ;
        RECT  1.955 0.205 2.025 0.415 ;
        RECT  1.890 0.845 2.010 1.055 ;
        RECT  1.440 0.345 1.955 0.415 ;
        RECT  0.990 0.845 1.890 0.915 ;
        RECT  0.130 0.985 1.650 1.055 ;
        RECT  1.370 0.205 1.440 0.415 ;
        RECT  0.875 0.205 1.370 0.275 ;
        RECT  0.805 0.205 0.875 0.915 ;
        RECT  0.390 0.205 0.805 0.275 ;
        RECT  0.210 0.845 0.805 0.915 ;
        RECT  0.050 0.875 0.130 1.055 ;
    END
END AO222D4BWP

MACRO AO22D0BWP
    CLASS CORE ;
    FOREIGN AO22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.185 1.225 1.045 ;
        RECT  1.135 0.185 1.155 0.315 ;
        RECT  1.135 0.895 1.155 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.440 0.190 0.565 ;
        RECT  0.035 0.440 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.670 0.900 0.740 ;
        RECT  0.735 0.345 0.805 0.740 ;
        RECT  0.405 0.345 0.735 0.415 ;
        RECT  0.315 0.345 0.405 0.485 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.495 0.665 0.765 ;
        RECT  0.545 0.685 0.575 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.600 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.960 -0.115 1.260 0.115 ;
        RECT  0.840 -0.115 0.960 0.135 ;
        RECT  0.125 -0.115 0.840 0.115 ;
        RECT  0.055 -0.115 0.125 0.290 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.145 1.260 1.375 ;
        RECT  0.880 0.995 1.000 1.375 ;
        RECT  0.125 1.145 0.880 1.375 ;
        RECT  0.055 0.925 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.460 1.065 0.925 ;
        RECT  0.985 0.460 0.995 0.530 ;
        RECT  0.465 0.855 0.995 0.925 ;
        RECT  0.910 0.205 0.985 0.530 ;
        RECT  0.420 0.205 0.910 0.275 ;
        RECT  0.210 0.995 0.780 1.065 ;
    END
END AO22D0BWP

MACRO AO22D1BWP
    CLASS CORE ;
    FOREIGN AO22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.185 1.225 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.355 0.550 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.115 1.260 0.115 ;
        RECT  0.930 -0.115 1.050 0.270 ;
        RECT  0.850 -0.115 0.930 0.115 ;
        RECT  0.775 -0.115 0.850 0.260 ;
        RECT  0.130 -0.115 0.775 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.025 1.145 1.260 1.375 ;
        RECT  0.955 0.990 1.025 1.375 ;
        RECT  0.330 1.145 0.955 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.345 1.065 0.915 ;
        RECT  0.700 0.345 0.995 0.415 ;
        RECT  0.570 0.845 0.995 0.915 ;
        RECT  0.485 0.995 0.870 1.065 ;
        RECT  0.630 0.205 0.700 0.415 ;
        RECT  0.380 0.205 0.630 0.275 ;
        RECT  0.415 0.845 0.485 1.065 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO22D1BWP

MACRO AO22D2BWP
    CLASS CORE ;
    FOREIGN AO22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 0.365 1.365 0.765 ;
        RECT  1.295 0.185 1.305 1.075 ;
        RECT  1.235 0.185 1.295 0.465 ;
        RECT  1.235 0.675 1.295 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.405 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.670 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.310 ;
        RECT  1.150 -0.115 1.410 0.115 ;
        RECT  1.030 -0.115 1.150 0.270 ;
        RECT  0.950 -0.115 1.030 0.115 ;
        RECT  0.880 -0.115 0.950 0.260 ;
        RECT  0.130 -0.115 0.880 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.850 1.490 1.375 ;
        RECT  1.125 1.145 1.410 1.375 ;
        RECT  1.055 0.990 1.125 1.375 ;
        RECT  0.340 1.145 1.055 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.095 0.345 1.165 0.915 ;
        RECT  0.810 0.345 1.095 0.415 ;
        RECT  0.630 0.845 1.095 0.915 ;
        RECT  0.515 0.985 0.970 1.055 ;
        RECT  0.740 0.205 0.810 0.415 ;
        RECT  0.400 0.205 0.740 0.275 ;
        RECT  0.445 0.845 0.515 1.055 ;
        RECT  0.125 0.845 0.445 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO22D2BWP

MACRO AO22D4BWP
    CLASS CORE ;
    FOREIGN AO22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.485 ;
        RECT  2.275 0.710 2.285 1.045 ;
        RECT  2.215 0.185 2.275 1.045 ;
        RECT  2.065 0.355 2.215 0.830 ;
        RECT  1.925 0.355 2.065 0.485 ;
        RECT  1.925 0.710 2.065 0.830 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.710 1.925 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.640 ;
        RECT  0.595 0.520 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 0.355 0.525 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.775 ;
        RECT  0.945 0.705 1.435 0.775 ;
        RECT  0.875 0.495 0.945 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.355 1.225 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.770 -0.115 2.010 0.115 ;
        RECT  1.650 -0.115 1.770 0.260 ;
        RECT  1.565 -0.115 1.650 0.115 ;
        RECT  1.495 -0.115 1.565 0.260 ;
        RECT  0.845 -0.115 1.495 0.115 ;
        RECT  0.775 -0.115 0.845 0.275 ;
        RECT  0.130 -0.115 0.775 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.680 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.900 2.130 1.375 ;
        RECT  1.745 1.145 2.010 1.375 ;
        RECT  1.675 0.990 1.745 1.375 ;
        RECT  0.670 1.145 1.675 1.375 ;
        RECT  0.590 0.985 0.670 1.375 ;
        RECT  0.310 1.145 0.590 1.375 ;
        RECT  0.230 0.985 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.355 1.995 0.485 ;
        RECT  1.925 0.710 1.995 0.830 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.710 1.925 1.045 ;
        RECT  1.700 0.345 1.780 0.915 ;
        RECT  1.395 0.345 1.700 0.415 ;
        RECT  0.930 0.845 1.700 0.915 ;
        RECT  0.845 0.985 1.590 1.055 ;
        RECT  1.325 0.205 1.395 0.415 ;
        RECT  1.025 0.205 1.325 0.275 ;
        RECT  0.955 0.205 1.025 0.415 ;
        RECT  0.680 0.345 0.955 0.415 ;
        RECT  0.775 0.845 0.845 1.055 ;
        RECT  0.510 0.845 0.775 0.915 ;
        RECT  0.610 0.205 0.680 0.415 ;
        RECT  0.380 0.205 0.610 0.275 ;
        RECT  0.390 0.845 0.510 1.055 ;
        RECT  0.125 0.845 0.390 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO22D4BWP

MACRO AO31D0BWP
    CLASS CORE ;
    FOREIGN AO31D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.190 1.085 1.045 ;
        RECT  0.995 0.190 1.015 0.310 ;
        RECT  0.995 0.920 1.015 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.525 0.770 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.695 0.600 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.130 -0.115 0.780 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 1.120 1.375 ;
        RECT  0.790 0.995 0.910 1.375 ;
        RECT  0.000 1.145 0.790 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.925 0.520 0.945 0.640 ;
        RECT  0.855 0.205 0.925 0.925 ;
        RECT  0.570 0.205 0.855 0.275 ;
        RECT  0.125 0.855 0.855 0.925 ;
        RECT  0.210 0.995 0.710 1.065 ;
        RECT  0.055 0.855 0.125 1.005 ;
    END
END AO31D0BWP

MACRO AO31D1BWP
    CLASS CORE ;
    FOREIGN AO31D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.190 1.085 1.045 ;
        RECT  0.980 0.190 1.015 0.470 ;
        RECT  0.980 0.760 1.015 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.640 ;
        RECT  0.595 0.355 0.665 0.485 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.555 0.580 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.880 0.145 ;
        RECT  0.140 -0.115 0.760 0.115 ;
        RECT  0.040 -0.115 0.140 0.290 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 1.145 1.120 1.375 ;
        RECT  0.770 0.985 0.870 1.375 ;
        RECT  0.000 1.145 0.770 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 0.520 0.925 0.640 ;
        RECT  0.835 0.215 0.905 0.915 ;
        RECT  0.570 0.215 0.835 0.285 ;
        RECT  0.125 0.845 0.835 0.915 ;
        RECT  0.210 0.985 0.690 1.055 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO31D1BWP

MACRO AO31D2BWP
    CLASS CORE ;
    FOREIGN AO31D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.355 1.085 0.905 ;
        RECT  1.015 0.185 1.025 1.045 ;
        RECT  0.955 0.185 1.015 0.465 ;
        RECT  0.955 0.785 1.015 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.510 0.735 0.765 ;
        RECT  0.595 0.635 0.665 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.215 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.580 0.565 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.300 ;
        RECT  0.860 -0.115 1.130 0.115 ;
        RECT  0.760 -0.115 0.860 0.265 ;
        RECT  0.130 -0.115 0.760 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.960 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.985 0.850 1.375 ;
        RECT  0.000 1.145 0.770 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.875 0.520 0.910 0.640 ;
        RECT  0.805 0.335 0.875 0.915 ;
        RECT  0.690 0.335 0.805 0.405 ;
        RECT  0.125 0.845 0.805 0.915 ;
        RECT  0.570 0.195 0.690 0.405 ;
        RECT  0.210 0.985 0.690 1.055 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO31D2BWP

MACRO AO31D4BWP
    CLASS CORE ;
    FOREIGN AO31D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.485 ;
        RECT  2.275 0.700 2.285 1.035 ;
        RECT  2.215 0.185 2.275 1.035 ;
        RECT  2.065 0.355 2.215 0.820 ;
        RECT  1.925 0.355 2.065 0.485 ;
        RECT  1.925 0.700 2.065 0.820 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.700 1.925 1.035 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.070 0.495 1.130 0.640 ;
        RECT  1.000 0.495 1.070 0.780 ;
        RECT  0.245 0.710 1.000 0.780 ;
        RECT  0.125 0.495 0.245 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.345 0.930 0.640 ;
        RECT  0.385 0.345 0.840 0.415 ;
        RECT  0.315 0.345 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.760 -0.115 2.010 0.115 ;
        RECT  1.660 -0.115 1.760 0.270 ;
        RECT  1.580 -0.115 1.660 0.115 ;
        RECT  1.480 -0.115 1.580 0.270 ;
        RECT  1.230 -0.115 1.480 0.115 ;
        RECT  1.140 -0.115 1.230 0.280 ;
        RECT  0.130 -0.115 1.140 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.890 2.130 1.375 ;
        RECT  1.770 1.145 2.010 1.375 ;
        RECT  1.670 0.850 1.770 1.375 ;
        RECT  1.290 0.850 1.670 0.920 ;
        RECT  0.000 1.145 1.670 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.355 1.995 0.485 ;
        RECT  1.925 0.700 1.995 0.820 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.700 1.925 1.035 ;
        RECT  1.705 0.350 1.775 0.780 ;
        RECT  1.070 0.350 1.705 0.420 ;
        RECT  1.210 0.710 1.705 0.780 ;
        RECT  0.125 0.990 1.590 1.060 ;
        RECT  1.140 0.710 1.210 0.920 ;
        RECT  0.210 0.850 1.140 0.920 ;
        RECT  1.000 0.205 1.070 0.420 ;
        RECT  0.570 0.205 1.000 0.275 ;
        RECT  0.055 0.880 0.125 1.060 ;
    END
END AO31D4BWP

MACRO AO32D0BWP
    CLASS CORE ;
    FOREIGN AO32D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.190 1.505 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.970 0.495 1.015 0.645 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.830 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.115 1.540 0.115 ;
        RECT  1.235 -0.115 1.305 0.270 ;
        RECT  1.105 -0.115 1.235 0.115 ;
        RECT  1.035 -0.115 1.105 0.270 ;
        RECT  0.130 -0.115 1.035 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.540 1.375 ;
        RECT  1.210 0.995 1.330 1.375 ;
        RECT  0.940 1.145 1.210 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.345 1.345 0.915 ;
        RECT  0.725 0.345 1.275 0.415 ;
        RECT  0.125 0.845 1.275 0.915 ;
        RECT  0.220 0.985 1.130 1.055 ;
        RECT  0.655 0.195 0.725 0.415 ;
        RECT  0.055 0.845 0.125 1.045 ;
    END
END AO32D0BWP

MACRO AO32D1BWP
    CLASS CORE ;
    FOREIGN AO32D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.190 1.505 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.970 0.495 1.015 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.830 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.115 1.540 0.115 ;
        RECT  1.210 -0.115 1.330 0.260 ;
        RECT  1.110 -0.115 1.210 0.115 ;
        RECT  1.040 -0.115 1.110 0.260 ;
        RECT  0.130 -0.115 1.040 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.540 1.375 ;
        RECT  1.210 1.005 1.330 1.375 ;
        RECT  0.940 1.145 1.210 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.345 1.345 0.915 ;
        RECT  0.970 0.345 1.275 0.415 ;
        RECT  0.125 0.845 1.275 0.915 ;
        RECT  0.220 0.985 1.130 1.055 ;
        RECT  0.900 0.205 0.970 0.415 ;
        RECT  0.600 0.205 0.900 0.275 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO32D1BWP

MACRO AO32D2BWP
    CLASS CORE ;
    FOREIGN AO32D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.355 1.505 0.905 ;
        RECT  1.435 0.185 1.445 1.045 ;
        RECT  1.375 0.185 1.435 0.465 ;
        RECT  1.375 0.785 1.435 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.950 0.495 1.015 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.355 0.810 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.280 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.260 ;
        RECT  1.090 -0.115 1.170 0.115 ;
        RECT  1.020 -0.115 1.090 0.260 ;
        RECT  0.130 -0.115 1.020 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.980 1.630 1.375 ;
        RECT  1.305 1.145 1.550 1.375 ;
        RECT  1.190 0.985 1.305 1.375 ;
        RECT  0.920 1.145 1.190 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.000 1.145 0.800 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.235 0.345 1.305 0.915 ;
        RECT  0.950 0.345 1.235 0.415 ;
        RECT  0.125 0.845 1.235 0.915 ;
        RECT  0.220 0.985 1.110 1.055 ;
        RECT  0.880 0.205 0.950 0.415 ;
        RECT  0.600 0.205 0.880 0.275 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO32D2BWP

MACRO AO32D4BWP
    CLASS CORE ;
    FOREIGN AO32D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.705 0.485 ;
        RECT  2.695 0.710 2.705 1.050 ;
        RECT  2.635 0.185 2.695 1.050 ;
        RECT  2.485 0.355 2.635 0.830 ;
        RECT  2.345 0.355 2.485 0.485 ;
        RECT  2.345 0.710 2.485 0.830 ;
        RECT  2.275 0.185 2.345 0.485 ;
        RECT  2.275 0.710 2.345 1.050 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.495 1.925 0.770 ;
        RECT  1.365 0.700 1.850 0.770 ;
        RECT  1.265 0.495 1.365 0.770 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.355 1.645 0.630 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.135 0.640 ;
        RECT  1.015 0.495 1.085 0.770 ;
        RECT  0.190 0.700 1.015 0.770 ;
        RECT  0.120 0.520 0.190 0.770 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.345 0.945 0.630 ;
        RECT  0.385 0.345 0.850 0.415 ;
        RECT  0.295 0.345 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.475 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.280 ;
        RECT  2.165 -0.115 2.430 0.115 ;
        RECT  2.095 -0.115 2.165 0.260 ;
        RECT  2.010 -0.115 2.095 0.115 ;
        RECT  1.890 -0.115 2.010 0.250 ;
        RECT  1.290 -0.115 1.890 0.115 ;
        RECT  1.170 -0.115 1.290 0.265 ;
        RECT  0.130 -0.115 1.170 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.675 2.890 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 0.900 2.550 1.375 ;
        RECT  1.820 1.145 2.430 1.375 ;
        RECT  1.700 1.120 1.820 1.375 ;
        RECT  1.440 1.145 1.700 1.375 ;
        RECT  1.320 1.120 1.440 1.375 ;
        RECT  0.000 1.145 1.320 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.485 ;
        RECT  2.345 0.710 2.415 0.830 ;
        RECT  2.275 0.185 2.345 0.485 ;
        RECT  2.275 0.710 2.345 1.050 ;
        RECT  2.125 0.345 2.195 0.910 ;
        RECT  1.810 0.345 2.125 0.415 ;
        RECT  0.210 0.840 2.125 0.910 ;
        RECT  0.125 0.980 2.010 1.050 ;
        RECT  1.740 0.205 1.810 0.415 ;
        RECT  1.445 0.205 1.740 0.275 ;
        RECT  1.375 0.205 1.445 0.415 ;
        RECT  1.100 0.345 1.375 0.415 ;
        RECT  1.030 0.205 1.100 0.415 ;
        RECT  0.570 0.205 1.030 0.275 ;
        RECT  0.055 0.900 0.125 1.050 ;
    END
END AO32D4BWP

MACRO AO33D0BWP
    CLASS CORE ;
    FOREIGN AO33D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.195 1.505 1.045 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.520 1.150 0.640 ;
        RECT  1.015 0.355 1.085 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.680 0.520 0.735 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.575 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.540 0.115 ;
        RECT  1.180 -0.115 1.300 0.135 ;
        RECT  0.130 -0.115 1.180 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 0.985 1.300 1.375 ;
        RECT  0.900 1.145 1.180 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.205 1.345 0.915 ;
        RECT  0.580 0.205 1.275 0.275 ;
        RECT  0.125 0.845 1.275 0.915 ;
        RECT  0.210 0.985 1.100 1.055 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO33D0BWP

MACRO AO33D1BWP
    CLASS CORE ;
    FOREIGN AO33D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.195 1.505 1.075 ;
        RECT  1.400 0.195 1.435 0.475 ;
        RECT  1.400 0.665 1.435 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.520 1.150 0.640 ;
        RECT  1.015 0.355 1.085 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.680 0.520 0.735 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.540 0.115 ;
        RECT  1.180 -0.115 1.300 0.135 ;
        RECT  0.130 -0.115 1.180 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 0.985 1.300 1.375 ;
        RECT  0.900 1.145 1.180 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.205 1.330 0.915 ;
        RECT  0.580 0.205 1.260 0.275 ;
        RECT  0.130 0.845 1.260 0.915 ;
        RECT  0.210 0.985 1.100 1.055 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO33D1BWP

MACRO AO33D2BWP
    CLASS CORE ;
    FOREIGN AO33D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.355 1.505 0.765 ;
        RECT  1.435 0.195 1.450 1.075 ;
        RECT  1.380 0.195 1.435 0.475 ;
        RECT  1.380 0.675 1.435 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.520 1.130 0.640 ;
        RECT  1.015 0.355 1.085 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.670 0.520 0.735 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.300 ;
        RECT  1.260 -0.115 1.550 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.130 -0.115 1.140 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.840 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 0.985 1.280 1.375 ;
        RECT  0.880 1.145 1.160 1.375 ;
        RECT  0.760 1.125 0.880 1.375 ;
        RECT  0.000 1.145 0.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.205 1.310 0.915 ;
        RECT  0.560 0.205 1.240 0.275 ;
        RECT  0.125 0.845 1.240 0.915 ;
        RECT  0.210 0.985 1.080 1.055 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO33D2BWP

MACRO AO33D4BWP
    CLASS CORE ;
    FOREIGN AO33D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.485 ;
        RECT  3.115 0.710 3.125 1.050 ;
        RECT  3.055 0.185 3.115 1.050 ;
        RECT  2.905 0.355 3.055 0.830 ;
        RECT  2.765 0.355 2.905 0.485 ;
        RECT  2.765 0.710 2.905 0.830 ;
        RECT  2.695 0.185 2.765 0.485 ;
        RECT  2.695 0.710 2.765 1.050 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.495 2.345 0.780 ;
        RECT  1.390 0.710 2.270 0.780 ;
        RECT  1.295 0.495 1.390 0.780 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.520 2.120 0.640 ;
        RECT  1.995 0.345 2.065 0.640 ;
        RECT  1.595 0.345 1.995 0.415 ;
        RECT  1.505 0.345 1.595 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 1.925 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.780 ;
        RECT  1.080 0.495 1.155 0.615 ;
        RECT  0.195 0.710 1.155 0.780 ;
        RECT  0.125 0.520 0.195 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.965 0.640 ;
        RECT  0.385 0.345 0.875 0.415 ;
        RECT  0.295 0.345 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.475 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.280 ;
        RECT  2.610 -0.115 2.850 0.115 ;
        RECT  2.490 -0.115 2.610 0.280 ;
        RECT  2.405 -0.115 2.490 0.115 ;
        RECT  2.335 -0.115 2.405 0.280 ;
        RECT  1.285 -0.115 2.335 0.115 ;
        RECT  1.215 -0.115 1.285 0.275 ;
        RECT  0.130 -0.115 1.215 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.680 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.900 2.970 1.375 ;
        RECT  2.585 1.145 2.850 1.375 ;
        RECT  2.515 0.990 2.585 1.375 ;
        RECT  2.240 1.145 2.515 1.375 ;
        RECT  2.120 1.130 2.240 1.375 ;
        RECT  1.860 1.145 2.120 1.375 ;
        RECT  1.740 1.130 1.860 1.375 ;
        RECT  1.480 1.145 1.740 1.375 ;
        RECT  1.360 1.130 1.480 1.375 ;
        RECT  0.000 1.145 1.360 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.485 ;
        RECT  2.765 0.710 2.835 0.830 ;
        RECT  2.695 0.185 2.765 0.485 ;
        RECT  2.695 0.710 2.765 1.050 ;
        RECT  2.545 0.350 2.615 0.920 ;
        RECT  2.235 0.350 2.545 0.420 ;
        RECT  0.210 0.850 2.545 0.920 ;
        RECT  0.125 0.990 2.430 1.060 ;
        RECT  2.165 0.205 2.235 0.420 ;
        RECT  1.435 0.205 2.165 0.275 ;
        RECT  1.365 0.205 1.435 0.415 ;
        RECT  1.115 0.345 1.365 0.415 ;
        RECT  1.045 0.205 1.115 0.415 ;
        RECT  0.610 0.205 1.045 0.275 ;
        RECT  0.055 0.910 0.125 1.060 ;
    END
END AO33D4BWP

MACRO AOI211D0BWP
    CLASS CORE ;
    FOREIGN AOI211D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0723 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.770 0.275 ;
        RECT  0.455 0.205 0.525 0.925 ;
        RECT  0.125 0.205 0.455 0.275 ;
        RECT  0.210 0.855 0.455 0.925 ;
        RECT  0.035 0.205 0.125 0.345 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.310 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.135 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.920 0.930 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.995 0.570 1.065 ;
        RECT  0.055 0.915 0.125 1.065 ;
    END
END AOI211D0BWP

MACRO AOI211D1BWP
    CLASS CORE ;
    FOREIGN AOI211D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1431 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.770 0.275 ;
        RECT  0.455 0.205 0.525 0.905 ;
        RECT  0.125 0.205 0.455 0.275 ;
        RECT  0.210 0.825 0.455 0.905 ;
        RECT  0.035 0.205 0.125 0.345 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.420 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.135 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.840 0.850 0.940 1.375 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.570 1.055 ;
        RECT  0.055 0.905 0.125 1.055 ;
    END
END AOI211D1BWP

MACRO AOI211D2BWP
    CLASS CORE ;
    FOREIGN AOI211D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.845 1.470 0.915 ;
        RECT  0.875 0.205 1.290 0.275 ;
        RECT  0.875 0.775 0.945 0.915 ;
        RECT  0.805 0.205 0.875 0.915 ;
        RECT  0.670 0.345 0.805 0.415 ;
        RECT  0.735 0.775 0.805 0.915 ;
        RECT  0.590 0.185 0.670 0.415 ;
        RECT  0.330 0.345 0.590 0.415 ;
        RECT  0.210 0.205 0.330 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.640 ;
        RECT  0.595 0.520 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.130 0.495 0.245 0.775 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.550 0.640 ;
        RECT  1.435 0.495 1.505 0.775 ;
        RECT  1.085 0.705 1.435 0.775 ;
        RECT  1.015 0.520 1.085 0.775 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.255 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.420 ;
        RECT  0.900 -0.115 1.550 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.485 -0.115 0.780 0.115 ;
        RECT  0.415 -0.115 0.485 0.275 ;
        RECT  0.130 -0.115 0.415 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 1.680 1.375 ;
        RECT  0.390 0.990 0.510 1.375 ;
        RECT  0.000 1.145 0.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.555 0.905 1.625 1.055 ;
        RECT  0.665 0.985 1.555 1.055 ;
        RECT  0.595 0.845 0.665 1.055 ;
        RECT  0.125 0.845 0.595 0.915 ;
        RECT  0.055 0.845 0.125 0.995 ;
    END
END AOI211D2BWP

MACRO AOI211D4BWP
    CLASS CORE ;
    FOREIGN AOI211D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5352 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.020 0.190 3.140 0.415 ;
        RECT  2.740 0.345 3.020 0.415 ;
        RECT  2.620 0.190 2.740 0.415 ;
        RECT  2.370 0.345 2.620 0.415 ;
        RECT  2.250 0.190 2.370 0.415 ;
        RECT  2.010 0.345 2.250 0.415 ;
        RECT  1.890 0.190 2.010 0.415 ;
        RECT  0.735 0.345 1.890 0.415 ;
        RECT  0.735 0.775 1.610 0.905 ;
        RECT  0.525 0.345 0.735 0.905 ;
        RECT  0.210 0.345 0.525 0.415 ;
        RECT  0.125 0.775 0.525 0.905 ;
        RECT  0.055 0.775 0.125 1.070 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 3.100 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.415 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.460 ;
        RECT  2.920 -0.115 3.230 0.115 ;
        RECT  2.840 -0.115 2.920 0.275 ;
        RECT  2.530 -0.115 2.840 0.115 ;
        RECT  2.450 -0.115 2.530 0.275 ;
        RECT  2.170 -0.115 2.450 0.115 ;
        RECT  2.090 -0.115 2.170 0.275 ;
        RECT  1.810 -0.115 2.090 0.115 ;
        RECT  1.730 -0.115 1.810 0.275 ;
        RECT  1.440 -0.115 1.730 0.115 ;
        RECT  1.320 -0.115 1.440 0.130 ;
        RECT  1.060 -0.115 1.320 0.115 ;
        RECT  0.940 -0.115 1.060 0.130 ;
        RECT  0.000 -0.115 0.940 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.145 3.360 1.375 ;
        RECT  3.040 0.860 3.120 1.375 ;
        RECT  2.720 1.145 3.040 1.375 ;
        RECT  2.640 0.860 2.720 1.375 ;
        RECT  0.000 1.145 2.640 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 0.190 3.140 0.415 ;
        RECT  2.740 0.345 3.020 0.415 ;
        RECT  2.620 0.190 2.740 0.415 ;
        RECT  2.370 0.345 2.620 0.415 ;
        RECT  2.250 0.190 2.370 0.415 ;
        RECT  2.010 0.345 2.250 0.415 ;
        RECT  1.890 0.190 2.010 0.415 ;
        RECT  0.805 0.345 1.890 0.415 ;
        RECT  0.805 0.775 1.610 0.905 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.125 0.775 0.455 0.905 ;
        RECT  0.055 0.775 0.125 1.070 ;
        RECT  3.230 0.720 3.310 1.010 ;
        RECT  2.920 0.720 3.230 0.790 ;
        RECT  2.840 0.720 2.920 1.010 ;
        RECT  2.530 0.720 2.840 0.790 ;
        RECT  2.450 0.720 2.530 1.010 ;
        RECT  2.190 0.720 2.450 0.790 ;
        RECT  0.210 0.995 2.370 1.065 ;
        RECT  2.070 0.720 2.190 0.925 ;
        RECT  1.710 0.720 2.070 0.790 ;
        RECT  0.130 0.205 1.630 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI211D4BWP

MACRO AOI211XD0BWP
    CLASS CORE ;
    FOREIGN AOI211XD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1043 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.770 0.275 ;
        RECT  0.455 0.205 0.525 0.905 ;
        RECT  0.125 0.205 0.455 0.275 ;
        RECT  0.210 0.825 0.455 0.905 ;
        RECT  0.035 0.205 0.125 0.345 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.325 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.135 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.840 0.850 0.940 1.375 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.570 1.055 ;
        RECT  0.055 0.905 0.125 1.055 ;
    END
END AOI211XD0BWP

MACRO AOI211XD1BWP
    CLASS CORE ;
    FOREIGN AOI211XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1923 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.835 1.470 0.905 ;
        RECT  1.225 0.205 1.450 0.275 ;
        RECT  1.150 0.205 1.225 0.905 ;
        RECT  0.685 0.345 1.150 0.415 ;
        RECT  0.990 0.835 1.150 0.905 ;
        RECT  0.615 0.215 0.685 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 0.355 0.525 0.630 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.485 0.805 0.775 ;
        RECT  0.245 0.705 0.715 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        RECT  0.130 0.495 0.175 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.035 0.640 ;
        RECT  0.875 0.495 0.950 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.115 1.680 0.115 ;
        RECT  0.970 -0.115 1.050 0.260 ;
        RECT  0.890 -0.115 0.970 0.115 ;
        RECT  0.770 -0.115 0.890 0.260 ;
        RECT  0.510 -0.115 0.770 0.115 ;
        RECT  0.430 -0.115 0.510 0.280 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 1.680 1.375 ;
        RECT  0.410 1.125 0.550 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.555 0.755 1.625 1.055 ;
        RECT  0.125 0.985 1.555 1.055 ;
        RECT  0.220 0.845 0.750 0.915 ;
        RECT  0.055 0.875 0.125 1.055 ;
    END
END AOI211XD1BWP

MACRO AOI211XD2BWP
    CLASS CORE ;
    FOREIGN AOI211XD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3598 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.185 2.750 0.415 ;
        RECT  2.105 0.345 2.630 0.415 ;
        RECT  2.035 0.185 2.105 0.415 ;
        RECT  0.875 0.345 2.035 0.415 ;
        RECT  0.875 0.775 1.415 0.905 ;
        RECT  0.665 0.345 0.875 0.905 ;
        RECT  0.520 0.345 0.665 0.415 ;
        RECT  0.205 0.775 0.665 0.905 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 2.205 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.555 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.910 -0.115 3.360 0.115 ;
        RECT  2.830 -0.115 2.910 0.425 ;
        RECT  2.560 -0.115 2.830 0.115 ;
        RECT  2.440 -0.115 2.560 0.275 ;
        RECT  2.310 -0.115 2.440 0.115 ;
        RECT  2.190 -0.115 2.310 0.275 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.275 ;
        RECT  1.030 -0.115 1.830 0.115 ;
        RECT  0.890 -0.115 1.030 0.135 ;
        RECT  0.000 -0.115 0.890 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.145 3.360 1.375 ;
        RECT  3.210 0.735 3.290 1.375 ;
        RECT  2.930 1.145 3.210 1.375 ;
        RECT  2.830 0.850 2.930 1.375 ;
        RECT  2.560 1.145 2.830 1.375 ;
        RECT  2.460 0.850 2.560 1.375 ;
        RECT  0.000 1.145 2.460 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.630 0.185 2.750 0.415 ;
        RECT  2.105 0.345 2.630 0.415 ;
        RECT  2.035 0.185 2.105 0.415 ;
        RECT  0.945 0.345 2.035 0.415 ;
        RECT  0.945 0.775 1.415 0.905 ;
        RECT  0.520 0.345 0.595 0.415 ;
        RECT  0.205 0.775 0.595 0.905 ;
        RECT  3.035 0.710 3.105 1.035 ;
        RECT  2.725 0.710 3.035 0.780 ;
        RECT  2.655 0.710 2.725 1.035 ;
        RECT  1.650 0.710 2.655 0.780 ;
        RECT  2.190 0.850 2.310 1.055 ;
        RECT  1.950 0.985 2.190 1.055 ;
        RECT  1.830 0.850 1.950 1.055 ;
        RECT  1.565 0.985 1.830 1.055 ;
        RECT  1.495 0.670 1.565 1.055 ;
        RECT  0.125 0.985 1.495 1.055 ;
        RECT  0.350 0.205 1.210 0.275 ;
        RECT  0.055 0.740 0.125 1.055 ;
    END
END AOI211XD2BWP

MACRO AOI211XD4BWP
    CLASS CORE ;
    FOREIGN AOI211XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7196 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.470 0.205 5.590 0.415 ;
        RECT  4.985 0.345 5.470 0.415 ;
        RECT  4.915 0.185 4.985 0.415 ;
        RECT  4.085 0.345 4.915 0.415 ;
        RECT  4.015 0.185 4.085 0.415 ;
        RECT  3.545 0.345 4.015 0.415 ;
        RECT  3.475 0.185 3.545 0.415 ;
        RECT  1.575 0.345 3.475 0.415 ;
        RECT  1.575 0.715 2.850 0.895 ;
        RECT  1.365 0.345 1.575 0.895 ;
        RECT  0.930 0.345 1.365 0.415 ;
        RECT  0.210 0.715 1.365 0.895 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.495 5.845 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.495 4.305 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.685 0.495 2.765 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 1.255 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.750 -0.115 6.160 0.115 ;
        RECT  5.670 -0.115 5.750 0.420 ;
        RECT  5.390 -0.115 5.670 0.115 ;
        RECT  5.310 -0.115 5.390 0.260 ;
        RECT  5.190 -0.115 5.310 0.115 ;
        RECT  5.070 -0.115 5.190 0.260 ;
        RECT  4.830 -0.115 5.070 0.115 ;
        RECT  4.710 -0.115 4.830 0.275 ;
        RECT  4.290 -0.115 4.710 0.115 ;
        RECT  4.170 -0.115 4.290 0.275 ;
        RECT  3.910 -0.115 4.170 0.115 ;
        RECT  3.830 -0.115 3.910 0.260 ;
        RECT  3.750 -0.115 3.830 0.115 ;
        RECT  3.630 -0.115 3.750 0.275 ;
        RECT  3.390 -0.115 3.630 0.115 ;
        RECT  3.270 -0.115 3.390 0.275 ;
        RECT  2.280 -0.115 3.270 0.115 ;
        RECT  2.160 -0.115 2.280 0.135 ;
        RECT  1.800 -0.115 2.160 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.000 -0.115 1.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.925 1.145 6.160 1.375 ;
        RECT  5.855 0.850 5.925 1.375 ;
        RECT  5.565 1.145 5.855 1.375 ;
        RECT  5.495 0.850 5.565 1.375 ;
        RECT  5.195 1.145 5.495 1.375 ;
        RECT  5.125 0.850 5.195 1.375 ;
        RECT  4.815 1.145 5.125 1.375 ;
        RECT  4.745 0.850 4.815 1.375 ;
        RECT  0.000 1.145 4.745 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.470 0.205 5.590 0.415 ;
        RECT  4.985 0.345 5.470 0.415 ;
        RECT  4.915 0.185 4.985 0.415 ;
        RECT  4.085 0.345 4.915 0.415 ;
        RECT  4.015 0.185 4.085 0.415 ;
        RECT  3.545 0.345 4.015 0.415 ;
        RECT  3.475 0.185 3.545 0.415 ;
        RECT  1.645 0.345 3.475 0.415 ;
        RECT  1.645 0.715 2.850 0.895 ;
        RECT  0.930 0.345 1.295 0.415 ;
        RECT  0.210 0.715 1.295 0.895 ;
        RECT  6.035 0.710 6.105 1.045 ;
        RECT  5.745 0.710 6.035 0.780 ;
        RECT  5.675 0.710 5.745 1.045 ;
        RECT  5.385 0.710 5.675 0.780 ;
        RECT  5.315 0.710 5.385 1.045 ;
        RECT  5.005 0.710 5.315 0.780 ;
        RECT  4.935 0.710 5.005 1.045 ;
        RECT  4.625 0.710 4.935 0.780 ;
        RECT  4.555 0.710 4.625 1.045 ;
        RECT  3.090 0.835 4.555 0.905 ;
        RECT  3.005 0.985 4.470 1.055 ;
        RECT  2.935 0.755 3.005 1.055 ;
        RECT  0.125 0.985 2.935 1.055 ;
        RECT  0.750 0.205 2.490 0.275 ;
        RECT  0.055 0.730 0.125 1.055 ;
    END
END AOI211XD4BWP

MACRO AOI21D0BWP
    CLASS CORE ;
    FOREIGN AOI21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0635 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.195 0.540 0.915 ;
        RECT  0.230 0.845 0.455 0.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.640 0.495 0.735 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.840 0.115 ;
        RECT  0.660 -0.115 0.740 0.280 ;
        RECT  0.130 -0.115 0.660 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.660 0.930 0.740 1.375 ;
        RECT  0.000 1.145 0.660 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.580 1.055 ;
        RECT  0.055 0.895 0.125 1.055 ;
    END
END AOI21D0BWP

MACRO AOI21D1BWP
    CLASS CORE ;
    FOREIGN AOI21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1254 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.195 0.540 0.905 ;
        RECT  0.230 0.825 0.455 0.905 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.640 0.495 0.735 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.840 0.115 ;
        RECT  0.650 -0.115 0.730 0.410 ;
        RECT  0.130 -0.115 0.650 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.145 0.840 1.375 ;
        RECT  0.650 0.845 0.730 1.375 ;
        RECT  0.000 1.145 0.650 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.570 1.055 ;
        RECT  0.055 0.885 0.125 1.055 ;
    END
END AOI21D1BWP

MACRO AOI21D2BWP
    CLASS CORE ;
    FOREIGN AOI21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2268 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.185 1.220 0.285 ;
        RECT  1.010 0.215 1.120 0.285 ;
        RECT  0.580 0.845 1.050 0.915 ;
        RECT  0.940 0.215 1.010 0.415 ;
        RECT  0.525 0.345 0.940 0.415 ;
        RECT  0.510 0.710 0.580 0.915 ;
        RECT  0.415 0.185 0.525 0.415 ;
        RECT  0.390 0.710 0.510 0.780 ;
        RECT  0.390 0.345 0.415 0.415 ;
        RECT  0.310 0.345 0.390 0.780 ;
        RECT  0.125 0.345 0.310 0.415 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 0.495 1.000 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 0.355 1.225 0.630 ;
        RECT  1.135 0.355 1.140 0.765 ;
        RECT  1.070 0.520 1.135 0.765 ;
        RECT  0.720 0.695 1.070 0.765 ;
        RECT  0.650 0.495 0.720 0.765 ;
        RECT  0.530 0.495 0.650 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 -0.115 1.260 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.330 -0.115 0.750 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.145 1.260 1.375 ;
        RECT  0.230 1.010 0.300 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.915 1.205 1.055 ;
        RECT  0.440 0.985 1.135 1.055 ;
        RECT  0.370 0.860 0.440 1.055 ;
        RECT  0.125 0.860 0.370 0.930 ;
        RECT  0.055 0.860 0.125 1.015 ;
    END
END AOI21D2BWP

MACRO AOI21D4BWP
    CLASS CORE ;
    FOREIGN AOI21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.205 2.310 0.415 ;
        RECT  1.925 0.345 2.190 0.415 ;
        RECT  1.855 0.185 1.925 0.415 ;
        RECT  1.775 0.345 1.855 0.415 ;
        RECT  1.705 0.345 1.775 0.765 ;
        RECT  1.450 0.695 1.705 0.765 ;
        RECT  1.380 0.695 1.450 0.905 ;
        RECT  0.735 0.775 1.380 0.905 ;
        RECT  0.525 0.350 0.735 0.905 ;
        RECT  0.210 0.350 0.525 0.420 ;
        RECT  0.125 0.775 0.525 0.905 ;
        RECT  0.055 0.775 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.205 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.495 1.370 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.415 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.470 ;
        RECT  2.110 -0.115 2.390 0.115 ;
        RECT  2.030 -0.115 2.110 0.270 ;
        RECT  1.760 -0.115 2.030 0.115 ;
        RECT  1.660 -0.115 1.760 0.270 ;
        RECT  1.390 -0.115 1.660 0.115 ;
        RECT  1.310 -0.115 1.390 0.265 ;
        RECT  1.025 -0.115 1.310 0.115 ;
        RECT  0.955 -0.115 1.025 0.265 ;
        RECT  0.000 -0.115 0.955 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.110 1.145 2.390 1.375 ;
        RECT  2.030 0.840 2.110 1.375 ;
        RECT  1.750 1.145 2.030 1.375 ;
        RECT  1.680 0.980 1.750 1.375 ;
        RECT  0.000 1.145 1.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.190 0.205 2.310 0.415 ;
        RECT  1.925 0.345 2.190 0.415 ;
        RECT  1.855 0.185 1.925 0.415 ;
        RECT  1.775 0.345 1.855 0.415 ;
        RECT  1.705 0.345 1.775 0.765 ;
        RECT  1.450 0.695 1.705 0.765 ;
        RECT  1.380 0.695 1.450 0.905 ;
        RECT  0.805 0.775 1.380 0.905 ;
        RECT  0.210 0.350 0.455 0.420 ;
        RECT  0.125 0.775 0.455 0.905 ;
        RECT  0.055 0.775 0.125 1.045 ;
        RECT  2.215 0.700 2.285 1.020 ;
        RECT  1.925 0.700 2.215 0.770 ;
        RECT  1.855 0.700 1.925 1.020 ;
        RECT  1.600 0.840 1.855 0.910 ;
        RECT  1.530 0.840 1.600 1.045 ;
        RECT  1.490 0.290 1.570 0.415 ;
        RECT  0.210 0.975 1.530 1.045 ;
        RECT  1.230 0.345 1.490 0.415 ;
        RECT  1.110 0.205 1.230 0.415 ;
        RECT  0.885 0.345 1.110 0.415 ;
        RECT  0.815 0.205 0.885 0.415 ;
        RECT  0.130 0.205 0.815 0.280 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI21D4BWP

MACRO AOI221D0BWP
    CLASS CORE ;
    FOREIGN AOI221D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0674 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.205 1.060 0.275 ;
        RECT  0.735 0.205 0.805 0.415 ;
        RECT  0.385 0.345 0.735 0.415 ;
        RECT  0.340 0.345 0.385 0.735 ;
        RECT  0.315 0.345 0.340 0.915 ;
        RECT  0.125 0.345 0.315 0.415 ;
        RECT  0.270 0.665 0.315 0.915 ;
        RECT  0.210 0.845 0.270 0.915 ;
        RECT  0.035 0.185 0.125 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.070 0.495 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.965 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.485 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.305 ;
        RECT  0.665 -0.115 1.130 0.115 ;
        RECT  0.595 -0.115 0.665 0.260 ;
        RECT  0.510 -0.115 0.595 0.115 ;
        RECT  0.390 -0.115 0.510 0.260 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.920 1.210 1.375 ;
        RECT  0.000 1.145 1.130 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.905 1.025 1.065 ;
        RECT  0.690 0.995 0.955 1.065 ;
        RECT  0.750 0.835 0.870 0.925 ;
        RECT  0.490 0.835 0.750 0.905 ;
        RECT  0.570 0.980 0.690 1.065 ;
        RECT  0.420 0.835 0.490 1.055 ;
        RECT  0.125 0.985 0.420 1.055 ;
        RECT  0.055 0.890 0.125 1.055 ;
    END
END AOI221D0BWP

MACRO AOI221D1BWP
    CLASS CORE ;
    FOREIGN AOI221D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1349 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.205 1.060 0.275 ;
        RECT  0.735 0.205 0.805 0.415 ;
        RECT  0.385 0.345 0.735 0.415 ;
        RECT  0.310 0.345 0.385 0.915 ;
        RECT  0.125 0.345 0.310 0.415 ;
        RECT  0.210 0.845 0.310 0.915 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.070 0.495 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.485 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.965 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.485 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.400 ;
        RECT  0.665 -0.115 1.130 0.115 ;
        RECT  0.595 -0.115 0.665 0.260 ;
        RECT  0.510 -0.115 0.595 0.115 ;
        RECT  0.390 -0.115 0.510 0.260 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.910 1.210 1.375 ;
        RECT  0.000 1.145 1.130 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.570 0.845 1.050 0.915 ;
        RECT  0.125 0.985 0.870 1.055 ;
        RECT  0.055 0.895 0.125 1.055 ;
    END
END AOI221D1BWP

MACRO AOI221D2BWP
    CLASS CORE ;
    FOREIGN AOI221D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3212 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.905 0.205 2.025 0.275 ;
        RECT  1.835 0.205 1.905 0.415 ;
        RECT  1.430 0.345 1.835 0.415 ;
        RECT  1.295 0.205 1.430 0.415 ;
        RECT  0.865 0.345 1.295 0.415 ;
        RECT  0.130 0.845 0.890 0.915 ;
        RECT  0.735 0.185 0.865 0.415 ;
        RECT  0.125 0.345 0.735 0.415 ;
        RECT  0.105 0.845 0.130 1.045 ;
        RECT  0.105 0.215 0.125 0.415 ;
        RECT  0.035 0.215 0.105 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.355 2.075 0.630 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.655 0.775 ;
        RECT  1.225 0.705 1.575 0.775 ;
        RECT  1.150 0.495 1.225 0.775 ;
        RECT  1.015 0.495 1.150 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.775 ;
        RECT  0.245 0.705 0.735 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.280 ;
        RECT  1.765 -0.115 2.110 0.115 ;
        RECT  1.695 -0.115 1.765 0.265 ;
        RECT  1.070 -0.115 1.695 0.115 ;
        RECT  0.950 -0.115 1.070 0.275 ;
        RECT  0.530 -0.115 0.950 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.145 2.240 1.375 ;
        RECT  1.910 0.840 1.990 1.375 ;
        RECT  0.000 1.145 1.910 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.115 0.700 2.185 1.025 ;
        RECT  1.830 0.700 2.115 0.770 ;
        RECT  1.760 0.700 1.830 0.915 ;
        RECT  1.045 0.845 1.760 0.915 ;
        RECT  0.210 0.985 1.610 1.055 ;
        RECT  0.975 0.775 1.045 0.915 ;
    END
END AOI221D2BWP

MACRO AOI221D4BWP
    CLASS CORE ;
    FOREIGN AOI221D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2078 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.830 0.475 ;
        RECT  1.690 0.700 1.760 1.045 ;
        RECT  1.575 0.700 1.690 0.820 ;
        RECT  1.405 0.355 1.575 0.820 ;
        RECT  1.365 0.355 1.405 1.045 ;
        RECT  1.295 0.355 1.365 0.485 ;
        RECT  1.295 0.700 1.365 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.640 ;
        RECT  1.060 0.520 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 -0.115 2.240 0.115 ;
        RECT  1.900 -0.115 2.020 0.135 ;
        RECT  1.620 -0.115 1.900 0.115 ;
        RECT  1.500 -0.115 1.620 0.135 ;
        RECT  1.240 -0.115 1.500 0.115 ;
        RECT  1.120 -0.115 1.240 0.135 ;
        RECT  0.600 -0.115 1.120 0.115 ;
        RECT  0.600 0.205 0.690 0.275 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.000 -0.115 0.480 0.115 ;
        RECT  0.390 0.205 0.480 0.275 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.145 2.240 1.375 ;
        RECT  1.900 0.860 1.980 1.375 ;
        RECT  1.610 1.145 1.900 1.375 ;
        RECT  1.490 0.890 1.610 1.375 ;
        RECT  1.215 1.145 1.490 1.375 ;
        RECT  1.145 0.750 1.215 1.375 ;
        RECT  0.000 1.145 1.145 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.355 1.830 0.475 ;
        RECT  1.690 0.700 1.760 1.045 ;
        RECT  1.645 0.700 1.690 0.820 ;
        RECT  2.120 0.185 2.190 1.075 ;
        RECT  2.115 0.720 2.120 1.075 ;
        RECT  1.900 0.720 2.115 0.790 ;
        RECT  2.040 0.520 2.050 0.640 ;
        RECT  1.970 0.205 2.040 0.640 ;
        RECT  1.030 0.205 1.970 0.275 ;
        RECT  1.830 0.545 1.900 0.790 ;
        RECT  1.675 0.545 1.830 0.615 ;
        RECT  0.570 0.845 1.050 0.915 ;
        RECT  0.950 0.205 1.030 0.415 ;
        RECT  0.385 0.345 0.950 0.415 ;
        RECT  0.130 0.985 0.870 1.055 ;
        RECT  0.310 0.345 0.385 0.915 ;
        RECT  0.125 0.345 0.310 0.415 ;
        RECT  0.210 0.845 0.310 0.915 ;
        RECT  0.050 0.895 0.130 1.055 ;
        RECT  0.055 0.255 0.125 0.415 ;
    END
END AOI221D4BWP

MACRO AOI221XD4BWP
    CLASS CORE ;
    FOREIGN AOI221XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5476 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.705 4.145 1.010 ;
        RECT  3.785 0.705 4.075 0.775 ;
        RECT  3.580 0.345 3.990 0.415 ;
        RECT  3.715 0.705 3.785 0.915 ;
        RECT  3.580 0.705 3.715 0.775 ;
        RECT  3.510 0.345 3.580 0.775 ;
        RECT  3.425 0.705 3.510 0.775 ;
        RECT  3.355 0.705 3.425 0.915 ;
        RECT  3.065 0.705 3.355 0.775 ;
        RECT  2.995 0.705 3.065 0.915 ;
        RECT  2.705 0.705 2.995 0.775 ;
        RECT  2.635 0.705 2.705 0.915 ;
        RECT  2.555 0.705 2.635 0.775 ;
        RECT  2.345 0.345 2.555 0.775 ;
        RECT  1.890 0.345 2.345 0.415 ;
        RECT  1.225 0.705 2.345 0.775 ;
        RECT  1.155 0.550 1.225 0.775 ;
        RECT  0.845 0.550 1.155 0.620 ;
        RECT  0.775 0.185 0.845 0.620 ;
        RECT  0.510 0.345 0.775 0.415 ;
        RECT  0.390 0.205 0.510 0.415 ;
        RECT  0.125 0.345 0.390 0.415 ;
        RECT  0.055 0.275 0.125 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.665 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.645 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.235 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.665 0.495 3.325 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.495 4.025 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.250 -0.115 4.200 0.115 ;
        RECT  3.170 -0.115 3.250 0.275 ;
        RECT  2.890 -0.115 3.170 0.115 ;
        RECT  2.810 -0.115 2.890 0.275 ;
        RECT  1.620 -0.115 2.810 0.115 ;
        RECT  1.540 -0.115 1.620 0.275 ;
        RECT  1.220 -0.115 1.540 0.115 ;
        RECT  1.140 -0.115 1.220 0.275 ;
        RECT  0.670 -0.115 1.140 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.310 -0.115 0.590 0.115 ;
        RECT  0.230 -0.115 0.310 0.275 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 4.200 1.375 ;
        RECT  0.650 0.850 0.720 1.375 ;
        RECT  0.315 1.145 0.650 1.375 ;
        RECT  0.245 0.850 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.075 0.705 4.145 1.010 ;
        RECT  3.785 0.705 4.075 0.775 ;
        RECT  3.580 0.345 3.990 0.415 ;
        RECT  3.715 0.705 3.785 0.915 ;
        RECT  3.580 0.705 3.715 0.775 ;
        RECT  3.510 0.345 3.580 0.775 ;
        RECT  3.425 0.705 3.510 0.775 ;
        RECT  3.355 0.705 3.425 0.915 ;
        RECT  3.065 0.705 3.355 0.775 ;
        RECT  2.995 0.705 3.065 0.915 ;
        RECT  2.705 0.705 2.995 0.775 ;
        RECT  2.635 0.705 2.705 0.915 ;
        RECT  2.625 0.705 2.635 0.775 ;
        RECT  1.890 0.345 2.275 0.415 ;
        RECT  1.225 0.705 2.275 0.775 ;
        RECT  1.155 0.550 1.225 0.775 ;
        RECT  0.845 0.550 1.155 0.620 ;
        RECT  0.775 0.185 0.845 0.620 ;
        RECT  0.510 0.345 0.775 0.415 ;
        RECT  0.390 0.205 0.510 0.415 ;
        RECT  0.125 0.345 0.390 0.415 ;
        RECT  0.055 0.275 0.125 0.415 ;
        RECT  4.075 0.205 4.145 0.345 ;
        RECT  3.425 0.205 4.075 0.275 ;
        RECT  3.870 0.845 3.990 1.055 ;
        RECT  3.630 0.985 3.870 1.055 ;
        RECT  3.510 0.845 3.630 1.055 ;
        RECT  3.270 0.985 3.510 1.055 ;
        RECT  3.355 0.205 3.425 0.415 ;
        RECT  3.090 0.345 3.355 0.415 ;
        RECT  3.150 0.845 3.270 1.055 ;
        RECT  2.910 0.985 3.150 1.055 ;
        RECT  2.970 0.205 3.090 0.415 ;
        RECT  2.705 0.345 2.970 0.415 ;
        RECT  2.790 0.845 2.910 1.055 ;
        RECT  1.170 0.985 2.790 1.055 ;
        RECT  2.635 0.235 2.705 0.415 ;
        RECT  1.805 0.205 2.555 0.275 ;
        RECT  1.085 0.845 2.550 0.915 ;
        RECT  1.735 0.205 1.805 0.415 ;
        RECT  1.440 0.345 1.735 0.415 ;
        RECT  1.320 0.205 1.440 0.415 ;
        RECT  0.930 0.345 1.320 0.415 ;
        RECT  1.015 0.705 1.085 1.010 ;
        RECT  0.905 0.705 1.015 0.775 ;
        RECT  0.835 0.705 0.905 1.010 ;
        RECT  0.515 0.705 0.835 0.775 ;
        RECT  0.445 0.705 0.515 1.010 ;
        RECT  0.125 0.705 0.445 0.775 ;
        RECT  0.055 0.705 0.125 1.010 ;
    END
END AOI221XD4BWP

MACRO AOI222D0BWP
    CLASS CORE ;
    FOREIGN AOI222D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0857 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.125 0.415 ;
        RECT  0.525 0.345 1.015 0.415 ;
        RECT  0.455 0.195 0.525 0.905 ;
        RECT  0.210 0.825 0.455 0.905 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.495 1.435 0.640 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.270 ;
        RECT  0.130 -0.115 1.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.290 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.905 1.490 1.375 ;
        RECT  0.000 1.145 1.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.845 1.330 0.915 ;
        RECT  0.125 0.985 0.930 1.055 ;
        RECT  0.055 0.915 0.125 1.055 ;
    END
END AOI222D0BWP

MACRO AOI222D1BWP
    CLASS CORE ;
    FOREIGN AOI222D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1617 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.345 1.150 0.415 ;
        RECT  0.455 0.195 0.525 0.905 ;
        RECT  0.210 0.825 0.455 0.905 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.520 1.435 0.640 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.270 ;
        RECT  0.130 -0.115 1.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.750 1.490 1.375 ;
        RECT  0.000 1.145 1.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.845 1.330 1.055 ;
        RECT  0.660 0.845 1.210 0.915 ;
        RECT  0.130 0.985 0.970 1.055 ;
        RECT  0.050 0.895 0.130 1.055 ;
    END
END AOI222D1BWP

MACRO AOI222D2BWP
    CLASS CORE ;
    FOREIGN AOI222D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3026 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.205 2.130 0.275 ;
        RECT  1.850 0.205 1.920 0.415 ;
        RECT  1.570 0.345 1.850 0.415 ;
        RECT  1.500 0.205 1.570 0.415 ;
        RECT  1.200 0.205 1.500 0.275 ;
        RECT  1.130 0.205 1.200 0.415 ;
        RECT  0.945 0.345 1.130 0.415 ;
        RECT  0.870 0.345 0.945 0.775 ;
        RECT  0.125 0.345 0.870 0.415 ;
        RECT  0.850 0.705 0.870 0.775 ;
        RECT  0.735 0.705 0.850 0.915 ;
        RECT  0.130 0.845 0.735 0.915 ;
        RECT  0.035 0.845 0.130 1.045 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.495 2.390 0.640 ;
        RECT  2.275 0.495 2.345 0.775 ;
        RECT  1.925 0.705 2.275 0.775 ;
        RECT  1.855 0.495 1.925 0.775 ;
        RECT  1.790 0.495 1.855 0.640 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.095 0.630 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.650 0.775 ;
        RECT  1.090 0.705 1.570 0.775 ;
        RECT  1.015 0.495 1.090 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.545 0.760 0.615 ;
        RECT  0.595 0.545 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.420 ;
        RECT  1.745 -0.115 2.390 0.115 ;
        RECT  1.675 -0.115 1.745 0.275 ;
        RECT  1.050 -0.115 1.675 0.115 ;
        RECT  0.930 -0.115 1.050 0.275 ;
        RECT  0.510 -0.115 0.930 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.145 2.520 1.375 ;
        RECT  2.210 0.985 2.290 1.375 ;
        RECT  1.930 1.145 2.210 1.375 ;
        RECT  1.850 0.985 1.930 1.375 ;
        RECT  0.000 1.145 1.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.845 2.470 1.005 ;
        RECT  2.130 0.845 2.390 0.915 ;
        RECT  2.010 0.845 2.130 1.055 ;
        RECT  1.760 0.845 2.010 0.915 ;
        RECT  1.660 0.845 1.760 1.070 ;
        RECT  0.930 0.845 1.660 0.915 ;
        RECT  0.210 0.995 1.590 1.065 ;
    END
END AOI222D2BWP

MACRO AOI222D4BWP
    CLASS CORE ;
    FOREIGN AOI222D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.350 2.110 0.470 ;
        RECT  2.015 0.860 2.085 1.045 ;
        RECT  1.855 0.860 2.015 0.960 ;
        RECT  1.725 0.350 1.855 0.960 ;
        RECT  1.645 0.350 1.725 1.045 ;
        RECT  1.610 0.350 1.645 0.470 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.355 1.515 0.625 ;
        RECT  1.340 0.545 1.425 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.830 0.495 0.875 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.200 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.905 ;
        RECT  0.410 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.115 2.520 0.115 ;
        RECT  2.180 -0.115 2.300 0.140 ;
        RECT  1.920 -0.115 2.180 0.115 ;
        RECT  1.800 -0.115 1.920 0.140 ;
        RECT  1.540 -0.115 1.800 0.115 ;
        RECT  1.420 -0.115 1.540 0.140 ;
        RECT  0.190 -0.115 1.420 0.115 ;
        RECT  0.110 -0.115 0.190 0.420 ;
        RECT  0.000 -0.115 0.110 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.145 2.520 1.375 ;
        RECT  2.205 0.895 2.275 1.375 ;
        RECT  1.930 1.145 2.205 1.375 ;
        RECT  1.810 1.030 1.930 1.375 ;
        RECT  1.535 1.145 1.810 1.375 ;
        RECT  1.465 0.735 1.535 1.375 ;
        RECT  0.000 1.145 1.465 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.350 2.110 0.470 ;
        RECT  2.015 0.860 2.085 1.045 ;
        RECT  1.925 0.860 2.015 0.960 ;
        RECT  2.415 0.185 2.485 1.045 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.720 2.415 1.045 ;
        RECT  2.160 0.720 2.395 0.790 ;
        RECT  2.310 0.520 2.345 0.640 ;
        RECT  2.240 0.210 2.310 0.640 ;
        RECT  1.145 0.210 2.240 0.280 ;
        RECT  2.090 0.545 2.160 0.790 ;
        RECT  1.955 0.545 2.090 0.615 ;
        RECT  1.275 0.845 1.345 1.035 ;
        RECT  0.630 0.845 1.275 0.915 ;
        RECT  1.075 0.210 1.145 0.415 ;
        RECT  0.570 0.345 1.075 0.415 ;
        RECT  0.190 0.985 0.950 1.055 ;
        RECT  0.450 0.205 0.570 0.415 ;
        RECT  0.340 0.345 0.450 0.415 ;
        RECT  0.340 0.790 0.365 0.915 ;
        RECT  0.270 0.345 0.340 0.915 ;
        RECT  0.110 0.895 0.190 1.055 ;
    END
END AOI222D4BWP

MACRO AOI222XD4BWP
    CLASS CORE ;
    FOREIGN AOI222XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5228 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.770 0.710 4.850 1.035 ;
        RECT  4.290 0.710 4.770 0.780 ;
        RECT  4.290 0.345 4.700 0.415 ;
        RECT  4.210 0.345 4.290 0.780 ;
        RECT  3.255 0.710 4.210 0.780 ;
        RECT  3.045 0.345 3.255 0.780 ;
        RECT  1.740 0.345 3.045 0.415 ;
        RECT  1.670 0.345 1.740 0.475 ;
        RECT  1.415 0.405 1.670 0.475 ;
        RECT  1.345 0.345 1.415 0.475 ;
        RECT  0.930 0.345 1.345 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.495 0.735 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.225 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.495 2.955 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.930 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.495 4.725 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 -0.115 4.900 0.115 ;
        RECT  3.870 -0.115 3.950 0.275 ;
        RECT  3.590 -0.115 3.870 0.115 ;
        RECT  3.510 -0.115 3.590 0.275 ;
        RECT  2.340 -0.115 3.510 0.115 ;
        RECT  2.220 -0.115 2.340 0.135 ;
        RECT  1.960 -0.115 2.220 0.115 ;
        RECT  1.840 -0.115 1.960 0.135 ;
        RECT  0.670 -0.115 1.840 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.310 -0.115 0.590 0.115 ;
        RECT  0.230 -0.115 0.310 0.275 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.420 1.145 4.900 1.375 ;
        RECT  1.340 0.840 1.420 1.375 ;
        RECT  1.050 1.145 1.340 1.375 ;
        RECT  0.970 0.840 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.840 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.840 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.770 0.710 4.850 1.035 ;
        RECT  4.290 0.710 4.770 0.780 ;
        RECT  4.290 0.345 4.700 0.415 ;
        RECT  4.210 0.345 4.290 0.780 ;
        RECT  3.325 0.710 4.210 0.780 ;
        RECT  1.740 0.345 2.975 0.415 ;
        RECT  1.670 0.345 1.740 0.475 ;
        RECT  1.415 0.405 1.670 0.475 ;
        RECT  1.345 0.345 1.415 0.475 ;
        RECT  0.930 0.345 1.345 0.415 ;
        RECT  4.770 0.195 4.850 0.335 ;
        RECT  4.125 0.195 4.770 0.265 ;
        RECT  4.570 0.850 4.690 1.060 ;
        RECT  4.330 0.990 4.570 1.060 ;
        RECT  4.210 0.850 4.330 1.060 ;
        RECT  3.970 0.990 4.210 1.060 ;
        RECT  4.055 0.195 4.125 0.465 ;
        RECT  3.790 0.345 4.055 0.415 ;
        RECT  3.850 0.850 3.970 1.060 ;
        RECT  3.610 0.990 3.850 1.060 ;
        RECT  3.670 0.205 3.790 0.415 ;
        RECT  3.405 0.345 3.670 0.415 ;
        RECT  3.490 0.850 3.610 1.060 ;
        RECT  1.870 0.990 3.490 1.060 ;
        RECT  3.335 0.195 3.405 0.465 ;
        RECT  1.650 0.205 3.250 0.275 ;
        RECT  2.530 0.850 3.250 0.920 ;
        RECT  2.410 0.700 2.530 0.920 ;
        RECT  2.170 0.700 2.410 0.770 ;
        RECT  2.050 0.700 2.170 0.910 ;
        RECT  1.785 0.700 2.050 0.770 ;
        RECT  1.715 0.700 1.785 1.010 ;
        RECT  1.605 0.700 1.715 0.770 ;
        RECT  1.535 0.700 1.605 1.010 ;
        RECT  1.495 0.205 1.565 0.325 ;
        RECT  1.225 0.700 1.535 0.770 ;
        RECT  0.845 0.205 1.495 0.275 ;
        RECT  1.155 0.700 1.225 1.010 ;
        RECT  0.865 0.700 1.155 0.770 ;
        RECT  0.795 0.700 0.865 1.010 ;
        RECT  0.775 0.205 0.845 0.415 ;
        RECT  0.505 0.700 0.795 0.770 ;
        RECT  0.485 0.345 0.775 0.415 ;
        RECT  0.435 0.700 0.505 1.010 ;
        RECT  0.415 0.185 0.485 0.415 ;
        RECT  0.125 0.700 0.435 0.770 ;
        RECT  0.125 0.345 0.415 0.415 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.700 0.125 1.010 ;
    END
END AOI222XD4BWP

MACRO AOI22D0BWP
    CLASS CORE ;
    FOREIGN AOI22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0702 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.710 0.735 0.915 ;
        RECT  0.525 0.710 0.665 0.780 ;
        RECT  0.455 0.195 0.525 0.780 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.310 ;
        RECT  0.130 -0.115 0.850 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.980 1.375 ;
        RECT  0.240 1.010 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.855 0.915 0.925 1.055 ;
        RECT  0.545 0.985 0.855 1.055 ;
        RECT  0.475 0.870 0.545 1.055 ;
        RECT  0.125 0.870 0.475 0.940 ;
        RECT  0.055 0.870 0.125 1.055 ;
    END
END AOI22D0BWP

MACRO AOI22D1BWP
    CLASS CORE ;
    FOREIGN AOI22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1194 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.720 0.770 0.790 ;
        RECT  0.455 0.195 0.525 0.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.420 ;
        RECT  0.130 -0.115 0.850 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.980 1.375 ;
        RECT  0.240 1.015 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.865 0.930 1.005 ;
        RECT  0.580 0.865 0.850 0.935 ;
        RECT  0.460 0.865 0.580 1.075 ;
        RECT  0.130 0.865 0.460 0.935 ;
        RECT  0.050 0.865 0.130 1.005 ;
    END
END AOI22D1BWP

MACRO AOI22D2BWP
    CLASS CORE ;
    FOREIGN AOI22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2408 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.205 1.645 0.815 ;
        RECT  1.555 0.205 1.575 0.395 ;
        RECT  1.445 0.745 1.575 0.815 ;
        RECT  0.130 0.205 1.555 0.275 ;
        RECT  1.375 0.745 1.445 0.915 ;
        RECT  0.970 0.845 1.375 0.915 ;
        RECT  0.035 0.205 0.130 0.345 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.425 0.355 0.525 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.775 ;
        RECT  0.245 0.705 0.715 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.225 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.520 1.505 0.640 ;
        RECT  1.295 0.345 1.365 0.640 ;
        RECT  0.970 0.345 1.295 0.415 ;
        RECT  0.875 0.345 0.970 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 -0.115 1.680 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.520 -0.115 1.140 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.145 1.680 1.375 ;
        RECT  0.590 0.985 0.710 1.375 ;
        RECT  0.330 1.145 0.590 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.550 0.895 1.630 1.055 ;
        RECT  0.880 0.985 1.550 1.055 ;
        RECT  0.800 0.845 0.880 1.055 ;
        RECT  0.495 0.845 0.800 0.915 ;
        RECT  0.425 0.845 0.495 1.075 ;
        RECT  0.130 0.845 0.425 0.915 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END AOI22D2BWP

MACRO AOI22D4BWP
    CLASS CORE ;
    FOREIGN AOI22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4504 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.355 3.140 0.425 ;
        RECT  2.470 0.355 2.540 0.775 ;
        RECT  1.205 0.705 2.470 0.775 ;
        RECT  1.135 0.705 1.205 0.905 ;
        RECT  0.735 0.775 1.135 0.905 ;
        RECT  0.525 0.350 0.735 0.905 ;
        RECT  0.210 0.350 0.525 0.420 ;
        RECT  0.125 0.775 0.525 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.425 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.360 -0.115 3.360 0.115 ;
        RECT  2.240 -0.115 2.360 0.145 ;
        RECT  1.960 -0.115 2.240 0.115 ;
        RECT  1.880 -0.115 1.960 0.275 ;
        RECT  1.390 -0.115 1.880 0.115 ;
        RECT  1.310 -0.115 1.390 0.265 ;
        RECT  1.040 -0.115 1.310 0.115 ;
        RECT  0.960 -0.115 1.040 0.265 ;
        RECT  0.000 -0.115 0.960 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.685 3.310 1.375 ;
        RECT  2.920 1.145 3.230 1.375 ;
        RECT  2.840 0.860 2.920 1.375 ;
        RECT  2.540 1.145 2.840 1.375 ;
        RECT  2.460 0.990 2.540 1.375 ;
        RECT  2.140 1.145 2.460 1.375 ;
        RECT  2.060 0.990 2.140 1.375 ;
        RECT  1.780 1.145 2.060 1.375 ;
        RECT  1.680 0.990 1.780 1.375 ;
        RECT  0.000 1.145 1.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.540 0.355 3.140 0.425 ;
        RECT  2.470 0.355 2.540 0.775 ;
        RECT  1.205 0.705 2.470 0.775 ;
        RECT  1.135 0.705 1.205 0.905 ;
        RECT  0.805 0.775 1.135 0.905 ;
        RECT  0.210 0.350 0.455 0.420 ;
        RECT  0.125 0.775 0.455 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        RECT  3.230 0.215 3.310 0.375 ;
        RECT  2.170 0.215 3.230 0.285 ;
        RECT  3.045 0.710 3.115 1.000 ;
        RECT  2.725 0.710 3.045 0.790 ;
        RECT  2.655 0.710 2.725 1.025 ;
        RECT  2.360 0.850 2.655 0.920 ;
        RECT  2.240 0.850 2.360 1.060 ;
        RECT  1.970 0.850 2.240 0.920 ;
        RECT  2.050 0.215 2.170 0.415 ;
        RECT  1.790 0.345 2.050 0.415 ;
        RECT  1.850 0.850 1.970 1.060 ;
        RECT  1.385 0.850 1.850 0.920 ;
        RECT  1.670 0.205 1.790 0.415 ;
        RECT  1.470 0.205 1.590 0.415 ;
        RECT  1.230 0.345 1.470 0.415 ;
        RECT  1.315 0.850 1.385 1.045 ;
        RECT  0.210 0.975 1.315 1.045 ;
        RECT  1.110 0.205 1.230 0.415 ;
        RECT  0.890 0.345 1.110 0.415 ;
        RECT  0.820 0.210 0.890 0.415 ;
        RECT  0.130 0.210 0.820 0.280 ;
        RECT  0.050 0.210 0.130 0.370 ;
    END
END AOI22D4BWP

MACRO AOI31D0BWP
    CLASS CORE ;
    FOREIGN AOI31D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.215 0.740 0.285 ;
        RECT  0.525 0.855 0.570 0.925 ;
        RECT  0.455 0.215 0.525 0.925 ;
        RECT  0.125 0.855 0.455 0.925 ;
        RECT  0.035 0.855 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.640 ;
        RECT  0.790 0.520 0.875 0.640 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.940 0.270 ;
        RECT  0.130 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.130 0.290 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.910 0.930 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.220 0.995 0.770 1.065 ;
    END
END AOI31D0BWP

MACRO AOI31D1BWP
    CLASS CORE ;
    FOREIGN AOI31D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1541 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.205 0.760 0.275 ;
        RECT  0.130 0.855 0.545 0.925 ;
        RECT  0.315 0.205 0.385 0.375 ;
        RECT  0.105 0.305 0.315 0.375 ;
        RECT  0.105 0.855 0.130 1.045 ;
        RECT  0.035 0.305 0.105 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.790 0.495 0.875 0.640 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.455 0.245 0.775 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.450 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.355 0.670 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.410 ;
        RECT  0.170 -0.115 0.850 0.115 ;
        RECT  0.050 -0.115 0.170 0.225 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.845 0.930 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.650 0.805 0.720 1.065 ;
        RECT  0.220 0.995 0.650 1.065 ;
    END
END AOI31D1BWP

MACRO AOI31D2BWP
    CLASS CORE ;
    FOREIGN AOI31D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2656 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.335 1.450 0.405 ;
        RECT  1.290 0.335 1.365 0.920 ;
        RECT  1.090 0.335 1.290 0.405 ;
        RECT  0.210 0.850 1.290 0.920 ;
        RECT  1.020 0.205 1.090 0.405 ;
        RECT  0.570 0.205 1.020 0.275 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.645 0.625 ;
        RECT  1.435 0.540 1.575 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.065 0.495 1.135 0.780 ;
        RECT  0.245 0.710 1.065 0.780 ;
        RECT  0.170 0.495 0.245 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.950 0.630 ;
        RECT  0.430 0.345 0.875 0.415 ;
        RECT  0.315 0.345 0.430 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.510 -0.115 1.630 0.275 ;
        RECT  1.230 -0.115 1.510 0.115 ;
        RECT  1.160 -0.115 1.230 0.255 ;
        RECT  0.130 -0.115 1.160 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.145 1.680 1.375 ;
        RECT  1.320 1.130 1.440 1.375 ;
        RECT  0.000 1.145 1.320 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.770 1.605 1.060 ;
        RECT  0.130 0.990 1.535 1.060 ;
        RECT  0.050 0.880 0.130 1.060 ;
    END
END AOI31D2BWP

MACRO AOI31D4BWP
    CLASS CORE ;
    FOREIGN AOI31D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5714 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.020 0.205 3.140 0.415 ;
        RECT  2.740 0.345 3.020 0.415 ;
        RECT  2.620 0.205 2.740 0.415 ;
        RECT  2.545 0.345 2.620 0.415 ;
        RECT  2.415 0.345 2.545 0.905 ;
        RECT  0.735 0.775 2.415 0.905 ;
        RECT  0.525 0.350 0.735 0.905 ;
        RECT  0.210 0.350 0.525 0.420 ;
        RECT  0.125 0.775 0.525 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.435 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.430 ;
        RECT  2.920 -0.115 3.230 0.115 ;
        RECT  2.840 -0.115 2.920 0.275 ;
        RECT  2.520 -0.115 2.840 0.115 ;
        RECT  2.440 -0.115 2.520 0.275 ;
        RECT  2.120 -0.115 2.440 0.115 ;
        RECT  2.040 -0.115 2.120 0.275 ;
        RECT  1.745 -0.115 2.040 0.115 ;
        RECT  1.675 -0.115 1.745 0.270 ;
        RECT  0.000 -0.115 1.675 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 1.145 3.360 1.375 ;
        RECT  3.020 0.890 3.140 1.375 ;
        RECT  2.740 1.145 3.020 1.375 ;
        RECT  2.620 1.115 2.740 1.375 ;
        RECT  0.000 1.145 2.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 0.205 3.140 0.415 ;
        RECT  2.740 0.345 3.020 0.415 ;
        RECT  2.620 0.205 2.740 0.415 ;
        RECT  2.545 0.345 2.620 0.415 ;
        RECT  2.415 0.345 2.545 0.905 ;
        RECT  0.805 0.775 2.415 0.905 ;
        RECT  0.210 0.350 0.455 0.420 ;
        RECT  0.125 0.775 0.455 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        RECT  3.230 0.750 3.310 1.030 ;
        RECT  2.920 0.750 3.230 0.820 ;
        RECT  2.845 0.750 2.920 1.045 ;
        RECT  0.210 0.975 2.845 1.045 ;
        RECT  2.215 0.205 2.335 0.415 ;
        RECT  1.950 0.345 2.215 0.415 ;
        RECT  1.830 0.205 1.950 0.415 ;
        RECT  0.930 0.345 1.830 0.415 ;
        RECT  0.130 0.205 1.590 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI31D4BWP

MACRO AOI32D0BWP
    CLASS CORE ;
    FOREIGN AOI32D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0809 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.555 0.805 0.915 ;
        RECT  0.665 0.555 0.735 0.625 ;
        RECT  0.125 0.845 0.735 0.915 ;
        RECT  0.595 0.195 0.665 0.625 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.930 0.495 1.010 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.825 0.485 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.700 0.640 0.770 ;
        RECT  0.455 0.495 0.525 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.115 1.120 0.115 ;
        RECT  0.990 -0.115 1.070 0.300 ;
        RECT  0.130 -0.115 0.990 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.145 1.120 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.915 1.065 1.055 ;
        RECT  0.210 0.985 0.995 1.055 ;
    END
END AOI32D0BWP

MACRO AOI32D1BWP
    CLASS CORE ;
    FOREIGN AOI32D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1521 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.205 0.730 0.275 ;
        RECT  0.130 0.845 0.540 0.915 ;
        RECT  0.315 0.205 0.385 0.365 ;
        RECT  0.105 0.295 0.315 0.365 ;
        RECT  0.105 0.845 0.130 1.045 ;
        RECT  0.035 0.295 0.105 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.930 0.520 1.015 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.445 0.810 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.640 ;
        RECT  0.550 0.520 0.595 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.115 1.120 0.115 ;
        RECT  0.980 -0.115 1.080 0.270 ;
        RECT  0.170 -0.115 0.980 0.115 ;
        RECT  0.050 -0.115 0.170 0.215 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 1.145 1.120 1.375 ;
        RECT  0.815 0.985 0.885 1.375 ;
        RECT  0.000 1.145 0.815 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.845 1.065 1.005 ;
        RECT  0.720 0.845 0.995 0.915 ;
        RECT  0.650 0.845 0.720 1.055 ;
        RECT  0.210 0.985 0.650 1.055 ;
    END
END AOI32D1BWP

MACRO AOI32D2BWP
    CLASS CORE ;
    FOREIGN AOI32D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.205 1.690 0.275 ;
        RECT  1.270 0.205 1.505 0.345 ;
        RECT  1.200 0.205 1.270 0.920 ;
        RECT  0.570 0.205 1.200 0.275 ;
        RECT  0.210 0.850 1.200 0.920 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.770 ;
        RECT  1.505 0.700 1.855 0.770 ;
        RECT  1.435 0.495 1.505 0.770 ;
        RECT  1.340 0.495 1.435 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.630 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 0.495 1.130 0.780 ;
        RECT  0.245 0.710 1.060 0.780 ;
        RECT  0.170 0.495 0.245 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.965 0.640 ;
        RECT  0.415 0.345 0.875 0.415 ;
        RECT  0.315 0.345 0.415 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.420 ;
        RECT  1.300 -0.115 1.970 0.115 ;
        RECT  1.180 -0.115 1.300 0.135 ;
        RECT  0.130 -0.115 1.180 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.145 2.100 1.375 ;
        RECT  1.760 1.015 1.880 1.375 ;
        RECT  1.500 1.145 1.760 1.375 ;
        RECT  1.380 1.130 1.500 1.375 ;
        RECT  0.000 1.145 1.380 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 0.840 2.050 1.055 ;
        RECT  1.665 0.840 1.970 0.910 ;
        RECT  1.595 0.840 1.665 1.075 ;
        RECT  1.475 0.840 1.595 0.910 ;
        RECT  1.405 0.840 1.475 1.060 ;
        RECT  0.130 0.990 1.405 1.060 ;
        RECT  0.050 0.875 0.130 1.060 ;
    END
END AOI32D2BWP

MACRO AOI32D4BWP
    CLASS CORE ;
    FOREIGN AOI32D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.005 0.475 ;
        RECT  1.995 0.700 2.005 1.045 ;
        RECT  1.935 0.185 1.995 1.045 ;
        RECT  1.785 0.345 1.935 0.820 ;
        RECT  1.635 0.345 1.785 0.475 ;
        RECT  1.635 0.700 1.785 0.820 ;
        RECT  1.565 0.185 1.635 0.475 ;
        RECT  1.565 0.700 1.635 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.690 0.520 0.735 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.475 ;
        RECT  1.850 -0.115 2.110 0.115 ;
        RECT  1.730 -0.115 1.850 0.270 ;
        RECT  1.450 -0.115 1.730 0.115 ;
        RECT  1.370 -0.115 1.450 0.325 ;
        RECT  1.090 -0.115 1.370 0.115 ;
        RECT  1.020 -0.115 1.090 0.260 ;
        RECT  0.130 -0.115 1.020 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.675 2.190 1.375 ;
        RECT  1.850 1.145 2.110 1.375 ;
        RECT  1.730 0.890 1.850 1.375 ;
        RECT  1.470 1.145 1.730 1.375 ;
        RECT  1.350 0.890 1.470 1.375 ;
        RECT  0.900 1.145 1.350 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.635 0.345 1.715 0.475 ;
        RECT  1.635 0.700 1.715 0.820 ;
        RECT  1.565 0.185 1.635 0.475 ;
        RECT  1.565 0.700 1.635 1.045 ;
        RECT  1.495 0.545 1.610 0.615 ;
        RECT  1.425 0.395 1.495 0.820 ;
        RECT  1.265 0.395 1.425 0.465 ;
        RECT  1.265 0.750 1.425 0.820 ;
        RECT  1.125 0.545 1.355 0.615 ;
        RECT  1.195 0.185 1.265 0.465 ;
        RECT  1.195 0.750 1.265 1.045 ;
        RECT  1.055 0.345 1.125 0.915 ;
        RECT  0.210 0.985 1.090 1.055 ;
        RECT  0.950 0.345 1.055 0.415 ;
        RECT  0.130 0.845 1.055 0.915 ;
        RECT  0.880 0.205 0.950 0.415 ;
        RECT  0.580 0.205 0.880 0.275 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END AOI32D4BWP

MACRO AOI32XD4BWP
    CLASS CORE ;
    FOREIGN AOI32XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5898 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.715 4.145 1.005 ;
        RECT  1.575 0.715 4.075 0.785 ;
        RECT  1.960 0.345 2.370 0.415 ;
        RECT  1.890 0.345 1.960 0.485 ;
        RECT  1.575 0.415 1.890 0.485 ;
        RECT  1.365 0.345 1.575 0.785 ;
        RECT  0.990 0.345 1.365 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.665 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.255 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 4.035 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.495 3.045 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.345 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.965 -0.115 4.200 0.115 ;
        RECT  3.895 -0.115 3.965 0.275 ;
        RECT  3.605 -0.115 3.895 0.115 ;
        RECT  3.535 -0.115 3.605 0.275 ;
        RECT  0.685 -0.115 3.535 0.115 ;
        RECT  0.615 -0.115 0.685 0.275 ;
        RECT  0.315 -0.115 0.615 0.115 ;
        RECT  0.245 -0.115 0.315 0.275 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.145 4.200 1.375 ;
        RECT  1.530 1.005 1.650 1.375 ;
        RECT  1.280 1.145 1.530 1.375 ;
        RECT  1.160 1.005 1.280 1.375 ;
        RECT  0.880 1.145 1.160 1.375 ;
        RECT  0.800 0.860 0.880 1.375 ;
        RECT  0.500 1.145 0.800 1.375 ;
        RECT  0.420 0.860 0.500 1.375 ;
        RECT  0.125 1.145 0.420 1.375 ;
        RECT  0.055 0.770 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.075 0.715 4.145 1.005 ;
        RECT  1.645 0.715 4.075 0.785 ;
        RECT  1.960 0.345 2.370 0.415 ;
        RECT  1.890 0.345 1.960 0.485 ;
        RECT  1.645 0.415 1.890 0.485 ;
        RECT  0.990 0.345 1.295 0.415 ;
        RECT  4.075 0.270 4.145 0.415 ;
        RECT  3.810 0.345 4.075 0.415 ;
        RECT  3.870 0.865 3.990 1.075 ;
        RECT  3.630 0.865 3.870 0.935 ;
        RECT  3.690 0.205 3.810 0.415 ;
        RECT  3.425 0.345 3.690 0.415 ;
        RECT  3.510 0.865 3.630 1.075 ;
        RECT  3.090 0.865 3.510 0.935 ;
        RECT  3.355 0.185 3.425 0.415 ;
        RECT  2.610 0.345 3.355 0.415 ;
        RECT  2.525 0.205 3.270 0.275 ;
        RECT  2.970 0.865 3.090 1.075 ;
        RECT  2.730 0.865 2.970 0.935 ;
        RECT  2.610 0.865 2.730 1.075 ;
        RECT  2.370 0.865 2.610 0.935 ;
        RECT  2.455 0.205 2.525 0.440 ;
        RECT  1.805 0.205 2.455 0.275 ;
        RECT  2.250 0.865 2.370 1.075 ;
        RECT  2.010 0.865 2.250 0.935 ;
        RECT  1.890 0.865 2.010 1.075 ;
        RECT  1.065 0.865 1.890 0.935 ;
        RECT  1.735 0.205 1.805 0.325 ;
        RECT  0.875 0.205 1.650 0.275 ;
        RECT  0.995 0.720 1.065 1.000 ;
        RECT  0.685 0.720 0.995 0.790 ;
        RECT  0.805 0.205 0.875 0.415 ;
        RECT  0.505 0.345 0.805 0.415 ;
        RECT  0.615 0.720 0.685 1.000 ;
        RECT  0.305 0.720 0.615 0.790 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.125 0.345 0.435 0.415 ;
        RECT  0.235 0.720 0.305 1.000 ;
        RECT  0.055 0.245 0.125 0.415 ;
    END
END AOI32XD4BWP

MACRO AOI33D0BWP
    CLASS CORE ;
    FOREIGN AOI33D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0872 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.215 0.760 0.285 ;
        RECT  0.525 0.855 0.550 0.925 ;
        RECT  0.455 0.215 0.525 0.925 ;
        RECT  0.130 0.855 0.455 0.925 ;
        RECT  0.035 0.855 0.130 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.210 0.495 1.295 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.105 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.945 0.765 ;
        RECT  0.760 0.690 0.870 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.320 ;
        RECT  0.130 -0.115 1.270 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.270 0.920 1.350 1.375 ;
        RECT  0.970 1.145 1.270 1.375 ;
        RECT  0.850 0.985 0.970 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.845 1.155 1.050 ;
        RECT  0.770 0.845 1.085 0.915 ;
        RECT  0.700 0.845 0.770 1.065 ;
        RECT  0.220 0.995 0.700 1.065 ;
    END
END AOI33D0BWP

MACRO AOI33D1BWP
    CLASS CORE ;
    FOREIGN AOI33D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1727 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.215 0.740 0.345 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.035 0.845 0.130 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.210 0.495 1.295 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.105 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.815 0.495 0.875 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.355 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.400 ;
        RECT  0.130 -0.115 1.270 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.850 1.360 1.375 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.880 0.985 0.960 1.375 ;
        RECT  0.000 1.145 0.880 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.845 1.180 0.915 ;
        RECT  0.665 0.845 0.735 1.055 ;
        RECT  0.220 0.985 0.665 1.055 ;
    END
END AOI33D1BWP

MACRO AOI33D2BWP
    CLASS CORE ;
    FOREIGN AOI33D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2713 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.340 2.345 0.795 ;
        RECT  2.160 0.340 2.275 0.410 ;
        RECT  2.190 0.725 2.275 0.795 ;
        RECT  2.120 0.725 2.190 0.925 ;
        RECT  2.090 0.200 2.160 0.410 ;
        RECT  1.295 0.855 2.120 0.925 ;
        RECT  0.570 0.200 2.090 0.270 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.065 0.350 1.135 0.640 ;
        RECT  0.245 0.350 1.065 0.420 ;
        RECT  0.175 0.350 0.245 0.765 ;
        RECT  0.130 0.520 0.175 0.645 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.775 ;
        RECT  0.405 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.405 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.480 2.205 0.645 ;
        RECT  2.020 0.480 2.135 0.550 ;
        RECT  1.950 0.340 2.020 0.550 ;
        RECT  1.365 0.340 1.950 0.410 ;
        RECT  1.295 0.340 1.365 0.765 ;
        RECT  1.250 0.520 1.295 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0556 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.620 2.040 0.775 ;
        RECT  1.505 0.705 1.920 0.775 ;
        RECT  1.435 0.495 1.505 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0556 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.795 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 -0.115 2.380 0.115 ;
        RECT  2.240 -0.115 2.340 0.270 ;
        RECT  1.240 -0.115 2.240 0.115 ;
        RECT  1.120 -0.115 1.240 0.130 ;
        RECT  0.130 -0.115 1.120 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 2.380 1.375 ;
        RECT  0.930 0.985 1.050 1.375 ;
        RECT  0.690 1.145 0.930 1.375 ;
        RECT  0.570 0.985 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 0.915 2.330 1.065 ;
        RECT  1.205 0.995 2.260 1.065 ;
        RECT  1.135 0.755 1.205 1.065 ;
        RECT  0.845 0.845 1.135 0.915 ;
        RECT  0.775 0.845 0.845 1.075 ;
        RECT  0.485 0.845 0.775 0.915 ;
        RECT  0.415 0.845 0.485 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AOI33D2BWP

MACRO AOI33D4BWP
    CLASS CORE ;
    FOREIGN AOI33D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.350 1.830 0.475 ;
        RECT  1.730 0.860 1.810 1.045 ;
        RECT  1.575 0.860 1.730 0.960 ;
        RECT  1.445 0.350 1.575 0.960 ;
        RECT  1.365 0.350 1.445 1.045 ;
        RECT  1.355 0.350 1.365 0.475 ;
        RECT  1.355 0.750 1.365 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.130 0.640 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.675 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.660 0.495 0.735 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 -0.115 2.240 0.115 ;
        RECT  1.900 -0.115 2.020 0.135 ;
        RECT  1.640 -0.115 1.900 0.115 ;
        RECT  1.520 -0.115 1.640 0.135 ;
        RECT  1.240 -0.115 1.520 0.115 ;
        RECT  1.120 -0.115 1.240 0.135 ;
        RECT  0.130 -0.115 1.120 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 1.145 2.240 1.375 ;
        RECT  1.900 0.885 2.020 1.375 ;
        RECT  1.650 1.145 1.900 1.375 ;
        RECT  1.530 1.030 1.650 1.375 ;
        RECT  1.250 1.145 1.530 1.375 ;
        RECT  1.150 0.990 1.250 1.375 ;
        RECT  0.880 1.145 1.150 1.375 ;
        RECT  0.760 1.125 0.880 1.375 ;
        RECT  0.000 1.145 0.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.350 1.830 0.475 ;
        RECT  1.730 0.860 1.810 1.045 ;
        RECT  1.645 0.860 1.730 0.960 ;
        RECT  2.120 0.195 2.190 1.075 ;
        RECT  2.115 0.720 2.120 1.075 ;
        RECT  1.910 0.720 2.115 0.790 ;
        RECT  1.980 0.205 2.050 0.640 ;
        RECT  1.275 0.205 1.980 0.275 ;
        RECT  1.840 0.545 1.910 0.790 ;
        RECT  1.675 0.545 1.840 0.615 ;
        RECT  1.205 0.205 1.275 0.915 ;
        RECT  0.570 0.205 1.205 0.275 ;
        RECT  0.130 0.845 1.205 0.915 ;
        RECT  0.210 0.985 1.070 1.055 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END AOI33D4BWP

MACRO AOI33XD4BWP
    CLASS CORE ;
    FOREIGN AOI33XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5836 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.915 0.715 4.985 1.025 ;
        RECT  2.415 0.715 4.915 0.785 ;
        RECT  2.800 0.345 3.210 0.415 ;
        RECT  2.730 0.345 2.800 0.485 ;
        RECT  2.485 0.415 2.730 0.485 ;
        RECT  2.415 0.345 2.485 0.485 ;
        RECT  2.205 0.345 2.415 0.785 ;
        RECT  1.830 0.345 2.205 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.665 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.505 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 2.095 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.495 4.875 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 4.025 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.495 3.185 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.805 -0.115 5.040 0.115 ;
        RECT  4.735 -0.115 4.805 0.275 ;
        RECT  4.445 -0.115 4.735 0.115 ;
        RECT  4.375 -0.115 4.445 0.275 ;
        RECT  0.665 -0.115 4.375 0.115 ;
        RECT  0.595 -0.115 0.665 0.275 ;
        RECT  0.305 -0.115 0.595 0.115 ;
        RECT  0.235 -0.115 0.305 0.275 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.145 5.040 1.375 ;
        RECT  2.370 1.005 2.490 1.375 ;
        RECT  2.130 1.145 2.370 1.375 ;
        RECT  2.010 1.005 2.130 1.375 ;
        RECT  1.745 1.145 2.010 1.375 ;
        RECT  1.675 0.860 1.745 1.375 ;
        RECT  1.385 1.145 1.675 1.375 ;
        RECT  1.315 0.860 1.385 1.375 ;
        RECT  1.025 1.145 1.315 1.375 ;
        RECT  0.955 0.925 1.025 1.375 ;
        RECT  0.845 1.145 0.955 1.375 ;
        RECT  0.775 0.925 0.845 1.375 ;
        RECT  0.485 1.145 0.775 1.375 ;
        RECT  0.415 0.860 0.485 1.375 ;
        RECT  0.125 1.145 0.415 1.375 ;
        RECT  0.055 0.695 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.915 0.715 4.985 1.025 ;
        RECT  2.485 0.715 4.915 0.785 ;
        RECT  2.800 0.345 3.210 0.415 ;
        RECT  2.730 0.345 2.800 0.485 ;
        RECT  2.485 0.415 2.730 0.485 ;
        RECT  1.830 0.345 2.135 0.415 ;
        RECT  4.915 0.270 4.985 0.415 ;
        RECT  4.650 0.345 4.915 0.415 ;
        RECT  4.710 0.865 4.830 1.075 ;
        RECT  4.470 0.865 4.710 0.935 ;
        RECT  4.530 0.205 4.650 0.415 ;
        RECT  4.265 0.345 4.530 0.415 ;
        RECT  4.350 0.865 4.470 1.075 ;
        RECT  3.930 0.865 4.350 0.935 ;
        RECT  4.195 0.185 4.265 0.415 ;
        RECT  3.450 0.345 4.195 0.415 ;
        RECT  3.365 0.205 4.110 0.275 ;
        RECT  3.810 0.865 3.930 1.075 ;
        RECT  3.570 0.865 3.810 0.935 ;
        RECT  3.450 0.865 3.570 1.075 ;
        RECT  3.210 0.865 3.450 0.935 ;
        RECT  3.295 0.205 3.365 0.440 ;
        RECT  2.645 0.205 3.295 0.275 ;
        RECT  3.090 0.865 3.210 1.075 ;
        RECT  2.850 0.865 3.090 0.935 ;
        RECT  2.730 0.865 2.850 1.075 ;
        RECT  1.925 0.865 2.730 0.935 ;
        RECT  2.575 0.205 2.645 0.325 ;
        RECT  1.745 0.205 2.490 0.275 ;
        RECT  1.855 0.720 1.925 1.055 ;
        RECT  1.565 0.720 1.855 0.790 ;
        RECT  1.675 0.205 1.745 0.435 ;
        RECT  0.930 0.205 1.675 0.275 ;
        RECT  0.845 0.345 1.590 0.415 ;
        RECT  1.495 0.720 1.565 1.055 ;
        RECT  1.205 0.720 1.495 0.790 ;
        RECT  1.135 0.720 1.205 1.055 ;
        RECT  0.665 0.720 1.135 0.790 ;
        RECT  0.775 0.185 0.845 0.415 ;
        RECT  0.485 0.345 0.775 0.415 ;
        RECT  0.595 0.720 0.665 1.055 ;
        RECT  0.305 0.720 0.595 0.790 ;
        RECT  0.415 0.185 0.485 0.415 ;
        RECT  0.125 0.345 0.415 0.415 ;
        RECT  0.235 0.720 0.305 1.055 ;
        RECT  0.055 0.275 0.125 0.415 ;
    END
END AOI33XD4BWP

MACRO BENCD1BWP
    CLASS CORE ;
    FOREIGN BENCD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.740 0.125 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.1254 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.355 3.010 0.425 ;
        RECT  2.625 0.690 2.750 0.780 ;
        RECT  2.555 0.355 2.625 0.780 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.485 0.630 ;
        RECT  2.375 0.530 2.415 0.630 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.640 ;
        RECT  1.680 0.495 1.715 0.575 ;
        RECT  1.610 0.355 1.680 0.575 ;
        RECT  1.460 0.355 1.610 0.425 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0444 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 0.495 1.540 0.630 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.345 2.065 0.780 ;
        RECT  1.750 0.345 1.995 0.415 ;
        RECT  1.890 0.710 1.995 0.780 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.595 -0.115 3.220 0.115 ;
        RECT  2.525 -0.115 2.595 0.280 ;
        RECT  2.205 -0.115 2.525 0.115 ;
        RECT  2.135 -0.115 2.205 0.280 ;
        RECT  1.460 -0.115 2.135 0.115 ;
        RECT  1.360 -0.115 1.460 0.285 ;
        RECT  1.085 -0.115 1.360 0.115 ;
        RECT  1.015 -0.115 1.085 0.270 ;
        RECT  0.305 -0.115 1.015 0.115 ;
        RECT  0.235 -0.115 0.305 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.100 0.765 3.170 1.375 ;
        RECT  2.560 1.145 3.100 1.375 ;
        RECT  2.440 1.130 2.560 1.375 ;
        RECT  2.200 1.145 2.440 1.375 ;
        RECT  2.080 1.130 2.200 1.375 ;
        RECT  1.445 1.145 2.080 1.375 ;
        RECT  1.335 0.990 1.445 1.375 ;
        RECT  1.090 1.145 1.335 1.375 ;
        RECT  0.970 0.990 1.090 1.375 ;
        RECT  0.340 1.145 0.970 1.375 ;
        RECT  0.220 1.025 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.095 0.195 3.165 0.455 ;
        RECT  3.030 0.545 3.100 0.615 ;
        RECT  2.710 0.195 3.095 0.265 ;
        RECT  2.960 0.545 3.030 1.060 ;
        RECT  1.650 0.990 2.960 1.060 ;
        RECT  2.820 0.510 2.890 0.920 ;
        RECT  1.800 0.850 2.820 0.920 ;
        RECT  2.345 0.195 2.410 0.265 ;
        RECT  2.205 0.710 2.370 0.780 ;
        RECT  2.275 0.195 2.345 0.430 ;
        RECT  2.205 0.360 2.275 0.430 ;
        RECT  2.135 0.360 2.205 0.780 ;
        RECT  1.570 0.195 2.050 0.265 ;
        RECT  1.730 0.710 1.800 0.920 ;
        RECT  1.005 0.710 1.730 0.780 ;
        RECT  1.580 0.850 1.650 1.060 ;
        RECT  0.865 0.850 1.580 0.920 ;
        RECT  1.195 0.250 1.265 0.420 ;
        RECT  1.005 0.350 1.195 0.420 ;
        RECT  0.935 0.350 1.005 0.780 ;
        RECT  0.670 0.595 0.935 0.665 ;
        RECT  0.795 0.280 0.865 0.515 ;
        RECT  0.795 0.735 0.865 0.920 ;
        RECT  0.585 0.445 0.795 0.515 ;
        RECT  0.585 0.735 0.795 0.805 ;
        RECT  0.445 0.195 0.710 0.265 ;
        RECT  0.270 0.885 0.710 0.955 ;
        RECT  0.515 0.445 0.585 0.805 ;
        RECT  0.340 0.545 0.515 0.615 ;
        RECT  0.375 0.195 0.445 0.420 ;
        RECT  0.270 0.350 0.375 0.420 ;
        RECT  0.200 0.350 0.270 0.955 ;
        RECT  0.180 0.520 0.200 0.640 ;
    END
END BENCD1BWP

MACRO BENCD2BWP
    CLASS CORE ;
    FOREIGN BENCD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.185 0.305 0.465 ;
        RECT  0.245 0.740 0.305 1.040 ;
        RECT  0.235 0.185 0.245 1.040 ;
        RECT  0.175 0.355 0.235 0.905 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.345 4.690 0.415 ;
        RECT  4.375 0.345 4.445 0.780 ;
        RECT  4.210 0.345 4.375 0.415 ;
        RECT  3.725 0.710 4.375 0.780 ;
        RECT  3.655 0.710 3.725 0.910 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.185 0.545 3.300 0.625 ;
        RECT  2.975 0.495 3.185 0.625 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.0988 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.495 2.345 0.625 ;
        RECT  1.880 0.555 2.130 0.625 ;
        RECT  1.810 0.360 1.880 0.625 ;
        RECT  1.640 0.360 1.810 0.430 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0732 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.545 1.730 0.630 ;
        RECT  1.255 0.495 1.505 0.630 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.2710 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 0.710 3.150 0.780 ;
        RECT  2.650 0.555 2.720 0.780 ;
        RECT  2.625 0.555 2.650 0.625 ;
        RECT  2.555 0.345 2.625 0.625 ;
        RECT  2.025 0.345 2.555 0.415 ;
        RECT  1.955 0.345 2.025 0.465 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.915 -0.115 4.900 0.115 ;
        RECT  3.845 -0.115 3.915 0.300 ;
        RECT  3.325 -0.115 3.845 0.115 ;
        RECT  3.255 -0.115 3.325 0.280 ;
        RECT  3.125 -0.115 3.255 0.115 ;
        RECT  3.055 -0.115 3.125 0.280 ;
        RECT  2.785 -0.115 3.055 0.115 ;
        RECT  2.665 -0.115 2.785 0.135 ;
        RECT  1.625 -0.115 2.665 0.115 ;
        RECT  1.555 -0.115 1.625 0.290 ;
        RECT  1.245 -0.115 1.555 0.115 ;
        RECT  1.175 -0.115 1.245 0.280 ;
        RECT  0.485 -0.115 1.175 0.115 ;
        RECT  0.415 -0.115 0.485 0.270 ;
        RECT  0.125 -0.115 0.415 0.115 ;
        RECT  0.055 -0.115 0.125 0.290 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.145 4.900 1.375 ;
        RECT  4.560 1.130 4.680 1.375 ;
        RECT  3.945 1.145 4.560 1.375 ;
        RECT  3.825 1.130 3.945 1.375 ;
        RECT  3.560 1.145 3.825 1.375 ;
        RECT  3.440 1.130 3.560 1.375 ;
        RECT  2.960 1.145 3.440 1.375 ;
        RECT  2.840 1.130 2.960 1.375 ;
        RECT  1.270 1.145 2.840 1.375 ;
        RECT  1.150 0.990 1.270 1.375 ;
        RECT  0.520 1.145 1.150 1.375 ;
        RECT  0.400 1.025 0.520 1.375 ;
        RECT  0.125 1.145 0.400 1.375 ;
        RECT  0.055 0.970 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.775 0.195 4.845 0.475 ;
        RECT  4.775 0.745 4.845 1.060 ;
        RECT  4.125 0.195 4.775 0.265 ;
        RECT  4.010 0.990 4.775 1.060 ;
        RECT  4.595 0.520 4.665 0.920 ;
        RECT  3.875 0.850 4.595 0.920 ;
        RECT  3.585 0.545 4.295 0.615 ;
        RECT  4.055 0.195 4.125 0.465 ;
        RECT  3.705 0.395 4.055 0.465 ;
        RECT  3.805 0.850 3.875 1.060 ;
        RECT  1.410 0.990 3.805 1.060 ;
        RECT  3.635 0.185 3.705 0.465 ;
        RECT  3.515 0.545 3.585 0.920 ;
        RECT  1.560 0.850 3.515 0.920 ;
        RECT  3.445 0.185 3.505 0.465 ;
        RECT  3.435 0.185 3.445 0.780 ;
        RECT  3.375 0.350 3.435 0.780 ;
        RECT  2.895 0.350 3.375 0.420 ;
        RECT  3.250 0.710 3.375 0.780 ;
        RECT  1.870 0.205 2.970 0.275 ;
        RECT  2.825 0.350 2.895 0.640 ;
        RECT  1.710 0.710 2.570 0.780 ;
        RECT  1.750 0.195 1.870 0.275 ;
        RECT  1.490 0.710 1.560 0.920 ;
        RECT  1.185 0.710 1.490 0.780 ;
        RECT  1.185 0.350 1.470 0.420 ;
        RECT  1.340 0.850 1.410 1.060 ;
        RECT  1.045 0.850 1.340 0.920 ;
        RECT  1.115 0.350 1.185 0.780 ;
        RECT  0.850 0.595 1.115 0.665 ;
        RECT  0.975 0.735 1.045 0.920 ;
        RECT  0.955 0.280 1.025 0.515 ;
        RECT  0.765 0.735 0.975 0.805 ;
        RECT  0.765 0.445 0.955 0.515 ;
        RECT  0.450 0.885 0.890 0.955 ;
        RECT  0.625 0.195 0.870 0.265 ;
        RECT  0.695 0.445 0.765 0.805 ;
        RECT  0.530 0.520 0.695 0.640 ;
        RECT  0.555 0.195 0.625 0.420 ;
        RECT  0.450 0.350 0.555 0.420 ;
        RECT  0.380 0.350 0.450 0.955 ;
        RECT  0.320 0.545 0.380 0.615 ;
    END
END BENCD2BWP

MACRO BENCD4BWP
    CLASS CORE ;
    FOREIGN BENCD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.745 0.665 1.075 ;
        RECT  0.455 0.355 0.595 0.465 ;
        RECT  0.455 0.745 0.595 0.905 ;
        RECT  0.305 0.355 0.455 0.905 ;
        RECT  0.245 0.185 0.305 1.075 ;
        RECT  0.235 0.185 0.245 0.465 ;
        RECT  0.235 0.745 0.245 1.075 ;
        END
    END X2
    PIN S
        ANTENNADIFFAREA 0.4094 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.175 0.345 7.770 0.415 ;
        RECT  6.965 0.345 7.175 0.780 ;
        RECT  6.550 0.345 6.965 0.415 ;
        RECT  5.630 0.710 6.965 0.780 ;
        END
    END S
    PIN M2
        ANTENNAGATEAREA 0.1728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.495 5.145 0.765 ;
        RECT  5.050 0.495 5.075 0.625 ;
        END
    END M2
    PIN M1
        ANTENNAGATEAREA 0.1456 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.485 3.885 0.625 ;
        RECT  2.570 0.485 3.395 0.555 ;
        RECT  2.500 0.355 2.570 0.555 ;
        RECT  2.360 0.355 2.500 0.425 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.1520 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.430 0.640 ;
        END
    END M0
    PIN A
        ANTENNADIFFAREA 0.4766 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.710 4.990 0.780 ;
        RECT  4.165 0.345 4.375 0.780 ;
        RECT  2.650 0.345 4.165 0.415 ;
        RECT  4.110 0.710 4.165 0.780 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.260 -0.115 7.980 0.115 ;
        RECT  6.180 -0.115 6.260 0.305 ;
        RECT  5.840 -0.115 6.180 0.115 ;
        RECT  5.760 -0.115 5.840 0.305 ;
        RECT  5.445 -0.115 5.760 0.115 ;
        RECT  5.375 -0.115 5.445 0.280 ;
        RECT  5.085 -0.115 5.375 0.115 ;
        RECT  5.015 -0.115 5.085 0.280 ;
        RECT  4.660 -0.115 5.015 0.115 ;
        RECT  4.540 -0.115 4.660 0.135 ;
        RECT  4.240 -0.115 4.540 0.115 ;
        RECT  4.120 -0.115 4.240 0.135 ;
        RECT  2.370 -0.115 4.120 0.115 ;
        RECT  2.250 -0.115 2.370 0.270 ;
        RECT  1.960 -0.115 2.250 0.115 ;
        RECT  1.890 -0.115 1.960 0.270 ;
        RECT  1.570 -0.115 1.890 0.115 ;
        RECT  1.500 -0.115 1.570 0.270 ;
        RECT  0.850 -0.115 1.500 0.115 ;
        RECT  0.770 -0.115 0.850 0.280 ;
        RECT  0.510 -0.115 0.770 0.115 ;
        RECT  0.390 -0.115 0.510 0.280 ;
        RECT  0.125 -0.115 0.390 0.115 ;
        RECT  0.055 -0.115 0.125 0.465 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.750 1.145 7.980 1.375 ;
        RECT  7.670 0.860 7.750 1.375 ;
        RECT  7.400 1.145 7.670 1.375 ;
        RECT  7.280 1.130 7.400 1.375 ;
        RECT  6.290 1.145 7.280 1.375 ;
        RECT  6.170 1.005 6.290 1.375 ;
        RECT  5.930 1.145 6.170 1.375 ;
        RECT  5.810 1.005 5.930 1.375 ;
        RECT  5.560 1.145 5.810 1.375 ;
        RECT  5.440 1.130 5.560 1.375 ;
        RECT  5.175 1.145 5.440 1.375 ;
        RECT  5.055 1.130 5.175 1.375 ;
        RECT  4.800 1.145 5.055 1.375 ;
        RECT  4.680 1.130 4.800 1.375 ;
        RECT  4.420 1.145 4.680 1.375 ;
        RECT  4.300 1.130 4.420 1.375 ;
        RECT  1.940 1.145 4.300 1.375 ;
        RECT  1.870 1.000 1.940 1.375 ;
        RECT  1.580 1.145 1.870 1.375 ;
        RECT  1.480 0.840 1.580 1.375 ;
        RECT  0.850 1.145 1.480 1.375 ;
        RECT  0.770 0.925 0.850 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.125 1.145 0.390 1.375 ;
        RECT  0.055 0.695 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.245 0.345 7.770 0.415 ;
        RECT  6.550 0.345 6.895 0.415 ;
        RECT  5.630 0.710 6.895 0.780 ;
        RECT  4.445 0.710 4.990 0.780 ;
        RECT  2.650 0.345 4.095 0.415 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.745 0.665 1.075 ;
        RECT  0.525 0.355 0.595 0.465 ;
        RECT  0.525 0.745 0.595 0.905 ;
        RECT  7.855 0.195 7.925 0.475 ;
        RECT  7.855 0.720 7.925 1.045 ;
        RECT  6.465 0.195 7.855 0.265 ;
        RECT  7.565 0.720 7.855 0.790 ;
        RECT  7.385 0.540 7.775 0.615 ;
        RECT  7.495 0.720 7.565 1.060 ;
        RECT  6.370 0.990 7.495 1.060 ;
        RECT  7.305 0.540 7.385 0.920 ;
        RECT  5.720 0.850 7.305 0.920 ;
        RECT  5.540 0.545 6.865 0.615 ;
        RECT  6.395 0.195 6.465 0.465 ;
        RECT  6.045 0.390 6.395 0.465 ;
        RECT  5.975 0.185 6.045 0.465 ;
        RECT  5.625 0.390 5.975 0.465 ;
        RECT  5.650 0.850 5.720 1.060 ;
        RECT  2.085 0.990 5.650 1.060 ;
        RECT  5.555 0.185 5.625 0.465 ;
        RECT  5.470 0.545 5.540 0.920 ;
        RECT  2.270 0.850 5.470 0.920 ;
        RECT  5.320 0.350 5.390 0.780 ;
        RECT  5.290 0.350 5.320 0.420 ;
        RECT  5.240 0.710 5.320 0.780 ;
        RECT  5.170 0.210 5.290 0.420 ;
        RECT  4.810 0.350 5.170 0.420 ;
        RECT  3.120 0.205 4.870 0.275 ;
        RECT  4.740 0.350 4.810 0.615 ;
        RECT  4.495 0.545 4.740 0.615 ;
        RECT  2.410 0.710 4.030 0.780 ;
        RECT  3.050 0.195 3.120 0.275 ;
        RECT  2.470 0.195 3.050 0.265 ;
        RECT  2.200 0.710 2.270 0.920 ;
        RECT  1.920 0.710 2.200 0.780 ;
        RECT  1.920 0.350 2.190 0.420 ;
        RECT  2.015 0.850 2.085 1.060 ;
        RECT  1.745 0.850 2.015 0.920 ;
        RECT  1.850 0.350 1.920 0.780 ;
        RECT  1.350 0.545 1.850 0.615 ;
        RECT  1.695 0.355 1.765 0.475 ;
        RECT  1.675 0.700 1.745 0.920 ;
        RECT  1.385 0.355 1.695 0.425 ;
        RECT  1.385 0.700 1.675 0.770 ;
        RECT  1.315 0.205 1.385 0.425 ;
        RECT  1.315 0.700 1.385 0.860 ;
        RECT  1.200 0.355 1.315 0.425 ;
        RECT  1.200 0.700 1.315 0.770 ;
        RECT  1.010 0.205 1.230 0.275 ;
        RECT  1.010 0.865 1.230 0.935 ;
        RECT  1.130 0.355 1.200 0.770 ;
        RECT  0.890 0.515 1.130 0.640 ;
        RECT  0.935 0.205 1.010 0.445 ;
        RECT  0.935 0.725 1.010 0.935 ;
        RECT  0.820 0.370 0.935 0.445 ;
        RECT  0.820 0.725 0.935 0.795 ;
        RECT  0.750 0.370 0.820 0.795 ;
        RECT  0.555 0.545 0.750 0.615 ;
    END
END BENCD4BWP

MACRO BHDBWP
    CLASS CORE ;
    FOREIGN BHDBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNAGATEAREA 0.0288 ;
        ANTENNADIFFAREA 0.0264 ;
        DIRECTION INOUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 0.905 ;
        RECT  0.410 0.185 0.455 0.300 ;
        RECT  0.430 0.745 0.455 0.905 ;
        RECT  0.195 0.745 0.430 0.815 ;
        RECT  0.125 0.520 0.195 0.815 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.310 -0.115 0.560 0.115 ;
        RECT  0.230 -0.115 0.310 0.300 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.560 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.975 0.470 1.045 ;
        RECT  0.300 0.370 0.370 0.640 ;
        RECT  0.125 0.370 0.300 0.440 ;
        RECT  0.050 0.895 0.130 1.045 ;
        RECT  0.055 0.255 0.125 0.440 ;
    END
END BHDBWP

MACRO BMLD1BWP
    CLASS CORE ;
    FOREIGN BMLD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0496 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.635 3.325 0.905 ;
        RECT  3.255 0.520 3.290 0.905 ;
        RECT  3.220 0.520 3.255 0.705 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.355 1.225 0.640 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.060 ;
        RECT  3.500 0.185 3.535 0.290 ;
        RECT  3.515 0.770 3.535 1.060 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.405 0.520 0.420 0.640 ;
        RECT  0.315 0.520 0.405 0.905 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.355 2.345 0.640 ;
        RECT  2.210 0.520 2.255 0.640 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.495 1.430 0.640 ;
        RECT  1.295 0.495 1.385 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 -0.115 3.640 0.115 ;
        RECT  3.280 -0.115 3.400 0.135 ;
        RECT  2.355 -0.115 3.280 0.115 ;
        RECT  2.285 -0.115 2.355 0.270 ;
        RECT  1.340 -0.115 2.285 0.115 ;
        RECT  1.220 -0.115 1.340 0.135 ;
        RECT  0.340 -0.115 1.220 0.115 ;
        RECT  0.220 -0.115 0.340 0.130 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.145 3.640 1.375 ;
        RECT  3.280 1.000 3.400 1.375 ;
        RECT  2.380 1.145 3.280 1.375 ;
        RECT  2.260 1.130 2.380 1.375 ;
        RECT  1.380 1.145 2.260 1.375 ;
        RECT  1.260 1.130 1.380 1.375 ;
        RECT  0.360 1.145 1.260 1.375 ;
        RECT  0.240 1.125 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.405 0.365 3.465 0.640 ;
        RECT  3.395 0.205 3.405 0.640 ;
        RECT  3.335 0.205 3.395 0.435 ;
        RECT  2.805 0.205 3.335 0.275 ;
        RECT  3.150 0.345 3.165 0.470 ;
        RECT  3.150 0.770 3.165 1.050 ;
        RECT  3.095 0.345 3.150 1.050 ;
        RECT  3.080 0.345 3.095 0.840 ;
        RECT  3.025 0.520 3.080 0.640 ;
        RECT  2.945 0.990 3.010 1.060 ;
        RECT  2.945 0.345 3.000 0.445 ;
        RECT  2.875 0.345 2.945 1.060 ;
        RECT  0.510 0.990 2.875 1.060 ;
        RECT  2.735 0.205 2.805 0.905 ;
        RECT  2.560 0.230 2.630 0.905 ;
        RECT  2.470 0.230 2.560 0.300 ;
        RECT  2.415 0.520 2.485 0.920 ;
        RECT  1.725 0.850 2.415 0.920 ;
        RECT  2.140 0.710 2.170 0.780 ;
        RECT  2.070 0.195 2.140 0.780 ;
        RECT  2.050 0.520 2.070 0.780 ;
        RECT  2.010 0.520 2.050 0.640 ;
        RECT  1.940 0.710 1.970 0.780 ;
        RECT  1.870 0.205 1.940 0.780 ;
        RECT  1.065 0.205 1.870 0.275 ;
        RECT  1.850 0.710 1.870 0.780 ;
        RECT  1.725 0.345 1.790 0.415 ;
        RECT  1.655 0.345 1.725 0.920 ;
        RECT  1.500 0.345 1.570 0.920 ;
        RECT  1.410 0.345 1.500 0.415 ;
        RECT  0.750 0.850 1.500 0.920 ;
        RECT  1.065 0.710 1.190 0.780 ;
        RECT  0.995 0.205 1.065 0.780 ;
        RECT  0.855 0.200 0.925 0.780 ;
        RECT  0.265 0.200 0.855 0.270 ;
        RECT  0.820 0.680 0.855 0.780 ;
        RECT  0.680 0.340 0.750 0.920 ;
        RECT  0.650 0.340 0.680 0.460 ;
        RECT  0.655 0.785 0.680 0.920 ;
        RECT  0.560 0.520 0.610 0.640 ;
        RECT  0.490 0.370 0.560 0.905 ;
        RECT  0.440 0.985 0.510 1.060 ;
        RECT  0.410 0.370 0.490 0.440 ;
        RECT  0.475 0.785 0.490 0.905 ;
        RECT  0.120 0.985 0.440 1.055 ;
        RECT  0.245 0.200 0.265 0.445 ;
        RECT  0.195 0.200 0.245 0.640 ;
        RECT  0.175 0.375 0.195 0.640 ;
        RECT  0.105 0.185 0.125 0.305 ;
        RECT  0.105 0.755 0.120 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END BMLD1BWP

MACRO BMLD2BWP
    CLASS CORE ;
    FOREIGN BMLD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0500 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.635 3.325 0.905 ;
        RECT  3.255 0.520 3.290 0.905 ;
        RECT  3.220 0.520 3.255 0.705 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.355 1.225 0.640 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.380 3.745 0.845 ;
        RECT  3.590 0.380 3.675 0.450 ;
        RECT  3.545 0.775 3.675 0.845 ;
        RECT  3.520 0.215 3.590 0.450 ;
        RECT  3.475 0.775 3.545 1.065 ;
        RECT  3.450 0.215 3.520 0.285 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.405 0.520 0.420 0.640 ;
        RECT  0.315 0.520 0.405 0.905 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.355 2.345 0.640 ;
        RECT  2.210 0.520 2.255 0.640 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.495 1.430 0.640 ;
        RECT  1.295 0.495 1.385 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.660 -0.115 3.730 0.300 ;
        RECT  3.380 -0.115 3.660 0.115 ;
        RECT  3.260 -0.115 3.380 0.135 ;
        RECT  2.355 -0.115 3.260 0.115 ;
        RECT  2.285 -0.115 2.355 0.270 ;
        RECT  1.340 -0.115 2.285 0.115 ;
        RECT  1.220 -0.115 1.340 0.135 ;
        RECT  0.340 -0.115 1.220 0.115 ;
        RECT  0.220 -0.115 0.340 0.130 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.935 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.000 3.390 1.375 ;
        RECT  2.380 1.145 3.270 1.375 ;
        RECT  2.260 1.130 2.380 1.375 ;
        RECT  1.380 1.145 2.260 1.375 ;
        RECT  1.260 1.130 1.380 1.375 ;
        RECT  0.360 1.145 1.260 1.375 ;
        RECT  0.240 1.125 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.450 0.520 3.520 0.640 ;
        RECT  3.380 0.365 3.450 0.590 ;
        RECT  3.325 0.365 3.380 0.435 ;
        RECT  3.255 0.205 3.325 0.435 ;
        RECT  2.805 0.205 3.255 0.275 ;
        RECT  3.150 0.770 3.185 1.050 ;
        RECT  3.150 0.345 3.165 0.470 ;
        RECT  3.115 0.345 3.150 1.050 ;
        RECT  3.080 0.345 3.115 0.840 ;
        RECT  3.025 0.520 3.080 0.640 ;
        RECT  2.945 0.990 3.010 1.060 ;
        RECT  2.945 0.345 3.000 0.445 ;
        RECT  2.875 0.345 2.945 1.060 ;
        RECT  0.510 0.990 2.875 1.060 ;
        RECT  2.735 0.205 2.805 0.905 ;
        RECT  2.560 0.230 2.630 0.905 ;
        RECT  2.470 0.230 2.560 0.300 ;
        RECT  2.415 0.520 2.485 0.920 ;
        RECT  1.725 0.850 2.415 0.920 ;
        RECT  2.140 0.710 2.170 0.780 ;
        RECT  2.070 0.195 2.140 0.780 ;
        RECT  2.050 0.520 2.070 0.780 ;
        RECT  2.010 0.520 2.050 0.640 ;
        RECT  1.940 0.710 1.970 0.780 ;
        RECT  1.870 0.205 1.940 0.780 ;
        RECT  1.065 0.205 1.870 0.275 ;
        RECT  1.850 0.710 1.870 0.780 ;
        RECT  1.725 0.345 1.790 0.415 ;
        RECT  1.655 0.345 1.725 0.920 ;
        RECT  1.500 0.345 1.570 0.920 ;
        RECT  1.410 0.345 1.500 0.415 ;
        RECT  0.750 0.850 1.500 0.920 ;
        RECT  1.065 0.710 1.190 0.780 ;
        RECT  0.995 0.205 1.065 0.780 ;
        RECT  0.855 0.200 0.925 0.780 ;
        RECT  0.265 0.200 0.855 0.270 ;
        RECT  0.820 0.680 0.855 0.780 ;
        RECT  0.680 0.340 0.750 0.920 ;
        RECT  0.650 0.340 0.680 0.460 ;
        RECT  0.655 0.785 0.680 0.920 ;
        RECT  0.560 0.520 0.610 0.640 ;
        RECT  0.490 0.370 0.560 0.905 ;
        RECT  0.440 0.985 0.510 1.060 ;
        RECT  0.410 0.370 0.490 0.440 ;
        RECT  0.475 0.785 0.490 0.905 ;
        RECT  0.120 0.985 0.440 1.055 ;
        RECT  0.245 0.200 0.265 0.445 ;
        RECT  0.195 0.200 0.245 0.640 ;
        RECT  0.175 0.375 0.195 0.640 ;
        RECT  0.105 0.185 0.125 0.305 ;
        RECT  0.105 0.755 0.120 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END BMLD2BWP

MACRO BMLD4BWP
    CLASS CORE ;
    FOREIGN BMLD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN X2
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.370 0.495 4.460 0.765 ;
        END
    END X2
    PIN S
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.625 ;
        RECT  1.575 0.545 1.715 0.625 ;
        END
    END S
    PIN PP
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.200 5.085 0.485 ;
        RECT  5.075 0.785 5.085 1.075 ;
        RECT  5.015 0.200 5.075 1.075 ;
        RECT  4.865 0.200 5.015 0.905 ;
        RECT  4.610 0.200 4.865 0.280 ;
        RECT  4.725 0.785 4.865 0.905 ;
        RECT  4.655 0.785 4.725 1.075 ;
        END
    END PP
    PIN M1
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.520 0.590 0.640 ;
        RECT  0.475 0.520 0.545 0.905 ;
        RECT  0.455 0.775 0.475 0.905 ;
        END
    END M1
    PIN M0
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.355 3.185 0.640 ;
        RECT  3.070 0.520 3.115 0.640 ;
        END
    END M0
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.355 2.205 0.625 ;
        RECT  1.995 0.545 2.135 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 -0.115 5.320 0.115 ;
        RECT  5.195 -0.115 5.265 0.480 ;
        RECT  4.920 -0.115 5.195 0.115 ;
        RECT  4.800 -0.115 4.920 0.130 ;
        RECT  4.540 -0.115 4.800 0.115 ;
        RECT  4.420 -0.115 4.540 0.130 ;
        RECT  3.590 -0.115 4.420 0.115 ;
        RECT  3.510 -0.115 3.590 0.290 ;
        RECT  3.240 -0.115 3.510 0.115 ;
        RECT  3.120 -0.115 3.240 0.260 ;
        RECT  2.245 -0.115 3.120 0.115 ;
        RECT  2.125 -0.115 2.245 0.135 ;
        RECT  1.860 -0.115 2.125 0.115 ;
        RECT  1.740 -0.115 1.860 0.135 ;
        RECT  1.490 -0.115 1.740 0.115 ;
        RECT  1.370 -0.115 1.490 0.275 ;
        RECT  0.520 -0.115 1.370 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.120 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.120 0.465 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 1.145 5.320 1.375 ;
        RECT  5.195 0.735 5.265 1.375 ;
        RECT  4.930 1.145 5.195 1.375 ;
        RECT  4.810 0.985 4.930 1.375 ;
        RECT  4.545 1.145 4.810 1.375 ;
        RECT  4.475 0.905 4.545 1.375 ;
        RECT  3.625 1.145 4.475 1.375 ;
        RECT  3.505 1.130 3.625 1.375 ;
        RECT  3.240 1.145 3.505 1.375 ;
        RECT  3.120 1.130 3.240 1.375 ;
        RECT  1.900 1.145 3.120 1.375 ;
        RECT  1.780 1.130 1.900 1.375 ;
        RECT  1.515 1.145 1.780 1.375 ;
        RECT  1.395 1.130 1.515 1.375 ;
        RECT  0.520 1.145 1.395 1.375 ;
        RECT  0.400 1.130 0.520 1.375 ;
        RECT  0.120 1.145 0.400 1.375 ;
        RECT  0.050 0.765 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.610 0.200 4.795 0.280 ;
        RECT  4.725 0.785 4.795 0.905 ;
        RECT  4.655 0.785 4.725 1.075 ;
        RECT  4.650 0.350 4.730 0.640 ;
        RECT  4.525 0.350 4.650 0.420 ;
        RECT  4.455 0.200 4.525 0.420 ;
        RECT  3.960 0.200 4.455 0.270 ;
        RECT  4.300 0.845 4.390 0.915 ;
        RECT  4.300 0.355 4.350 0.425 ;
        RECT  4.230 0.355 4.300 0.915 ;
        RECT  4.185 0.520 4.230 0.640 ;
        RECT  4.105 0.990 4.195 1.060 ;
        RECT  4.105 0.340 4.160 0.440 ;
        RECT  4.035 0.340 4.105 1.060 ;
        RECT  0.305 0.990 4.035 1.060 ;
        RECT  3.890 0.200 3.960 0.910 ;
        RECT  3.715 0.205 3.785 0.920 ;
        RECT  3.695 0.205 3.715 0.450 ;
        RECT  3.310 0.850 3.715 0.920 ;
        RECT  3.405 0.380 3.695 0.450 ;
        RECT  3.335 0.190 3.405 0.450 ;
        RECT  3.335 0.520 3.405 0.780 ;
        RECT  3.210 0.710 3.335 0.780 ;
        RECT  3.140 0.710 3.210 0.920 ;
        RECT  2.615 0.850 3.140 0.920 ;
        RECT  3.000 0.710 3.050 0.780 ;
        RECT  3.000 0.240 3.020 0.380 ;
        RECT  2.930 0.240 3.000 0.780 ;
        RECT  2.920 0.545 2.930 0.780 ;
        RECT  2.850 0.545 2.920 0.615 ;
        RECT  2.790 0.325 2.845 0.445 ;
        RECT  2.780 0.710 2.840 0.780 ;
        RECT  2.780 0.205 2.790 0.445 ;
        RECT  2.710 0.205 2.780 0.780 ;
        RECT  1.645 0.205 2.710 0.275 ;
        RECT  2.615 0.355 2.640 0.485 ;
        RECT  2.545 0.355 2.615 0.920 ;
        RECT  2.380 0.345 2.450 0.920 ;
        RECT  2.320 0.345 2.380 0.415 ;
        RECT  1.925 0.850 2.380 0.920 ;
        RECT  1.925 0.345 2.050 0.415 ;
        RECT  1.855 0.345 1.925 0.920 ;
        RECT  0.910 0.850 1.855 0.920 ;
        RECT  1.285 0.710 1.710 0.780 ;
        RECT  1.575 0.205 1.645 0.420 ;
        RECT  1.285 0.350 1.575 0.420 ;
        RECT  1.210 0.225 1.285 0.780 ;
        RECT  1.070 0.205 1.140 0.775 ;
        RECT  0.515 0.205 1.070 0.275 ;
        RECT  0.980 0.685 1.070 0.775 ;
        RECT  0.840 0.345 0.910 0.920 ;
        RECT  0.800 0.775 0.840 0.920 ;
        RECT  0.730 0.520 0.770 0.640 ;
        RECT  0.660 0.355 0.730 0.915 ;
        RECT  0.590 0.355 0.660 0.425 ;
        RECT  0.620 0.795 0.660 0.915 ;
        RECT  0.445 0.205 0.515 0.420 ;
        RECT  0.400 0.350 0.445 0.420 ;
        RECT  0.330 0.350 0.400 0.640 ;
        RECT  0.260 0.210 0.330 0.280 ;
        RECT  0.260 0.760 0.305 1.060 ;
        RECT  0.235 0.210 0.260 1.060 ;
        RECT  0.190 0.210 0.235 0.830 ;
    END
END BMLD4BWP

MACRO BUFFD0BWP
    CLASS CORE ;
    FOREIGN BUFFD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.215 0.525 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.645 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.345 0.370 0.915 ;
        RECT  0.125 0.345 0.300 0.415 ;
        RECT  0.125 0.845 0.300 0.915 ;
        RECT  0.055 0.225 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END BUFFD0BWP

MACRO BUFFD12BWP
    CLASS CORE ;
    FOREIGN BUFFD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.6048 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.720 2.870 0.950 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.135 0.305 2.415 0.465 ;
        RECT  2.125 0.305 2.135 0.950 ;
        RECT  2.055 0.185 2.125 0.950 ;
        RECT  1.785 0.305 2.055 0.950 ;
        RECT  1.765 0.305 1.785 0.465 ;
        RECT  0.950 0.720 1.785 0.950 ;
        RECT  1.695 0.185 1.765 0.465 ;
        RECT  1.405 0.305 1.695 0.465 ;
        RECT  1.335 0.185 1.405 0.465 ;
        RECT  1.045 0.305 1.335 0.465 ;
        RECT  0.975 0.185 1.045 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.455 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.465 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.235 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.235 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.235 ;
        RECT  1.610 -0.115 1.850 0.115 ;
        RECT  1.490 -0.115 1.610 0.235 ;
        RECT  1.250 -0.115 1.490 0.115 ;
        RECT  1.130 -0.115 1.250 0.235 ;
        RECT  0.860 -0.115 1.130 0.115 ;
        RECT  0.780 -0.115 0.860 0.465 ;
        RECT  0.495 -0.115 0.780 0.115 ;
        RECT  0.405 -0.115 0.495 0.260 ;
        RECT  0.140 -0.115 0.405 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.680 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 1.020 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.020 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.020 1.970 1.375 ;
        RECT  1.610 1.145 1.850 1.375 ;
        RECT  1.490 1.020 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 1.020 1.250 1.375 ;
        RECT  0.860 1.145 1.130 1.375 ;
        RECT  0.780 0.720 0.860 1.375 ;
        RECT  0.490 1.145 0.780 1.375 ;
        RECT  0.410 0.995 0.490 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.720 2.870 0.950 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.205 0.305 2.415 0.465 ;
        RECT  1.695 0.185 1.715 0.465 ;
        RECT  0.950 0.720 1.715 0.950 ;
        RECT  1.405 0.305 1.695 0.465 ;
        RECT  1.335 0.185 1.405 0.465 ;
        RECT  1.045 0.305 1.335 0.465 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  2.235 0.545 2.855 0.615 ;
        RECT  0.690 0.545 1.695 0.615 ;
        RECT  0.580 0.195 0.690 1.050 ;
        RECT  0.330 0.335 0.580 0.415 ;
        RECT  0.305 0.845 0.580 0.925 ;
        RECT  0.210 0.205 0.330 0.415 ;
        RECT  0.235 0.845 0.305 0.985 ;
    END
END BUFFD12BWP

MACRO BUFFD16BWP
    CLASS CORE ;
    FOREIGN BUFFD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.8064 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.715 3.850 0.945 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.465 0.305 3.755 0.465 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.105 0.305 3.395 0.465 ;
        RECT  3.035 0.185 3.105 0.465 ;
        RECT  2.835 0.305 3.035 0.465 ;
        RECT  2.745 0.305 2.835 0.945 ;
        RECT  2.675 0.185 2.745 0.945 ;
        RECT  2.485 0.305 2.675 0.945 ;
        RECT  2.385 0.305 2.485 0.465 ;
        RECT  1.210 0.715 2.485 0.945 ;
        RECT  2.315 0.185 2.385 0.465 ;
        RECT  2.025 0.305 2.315 0.465 ;
        RECT  1.955 0.185 2.025 0.465 ;
        RECT  1.665 0.305 1.955 0.465 ;
        RECT  1.595 0.185 1.665 0.465 ;
        RECT  1.305 0.305 1.595 0.465 ;
        RECT  1.235 0.185 1.305 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.665 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.465 ;
        RECT  3.670 -0.115 3.930 0.115 ;
        RECT  3.550 -0.115 3.670 0.235 ;
        RECT  3.310 -0.115 3.550 0.115 ;
        RECT  3.190 -0.115 3.310 0.235 ;
        RECT  2.950 -0.115 3.190 0.115 ;
        RECT  2.830 -0.115 2.950 0.235 ;
        RECT  2.590 -0.115 2.830 0.115 ;
        RECT  2.470 -0.115 2.590 0.235 ;
        RECT  2.230 -0.115 2.470 0.115 ;
        RECT  2.110 -0.115 2.230 0.235 ;
        RECT  1.870 -0.115 2.110 0.115 ;
        RECT  1.750 -0.115 1.870 0.235 ;
        RECT  1.510 -0.115 1.750 0.115 ;
        RECT  1.390 -0.115 1.510 0.235 ;
        RECT  1.100 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.100 0.465 ;
        RECT  0.720 -0.115 1.020 0.115 ;
        RECT  0.600 -0.115 0.720 0.265 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.680 4.010 1.375 ;
        RECT  3.670 1.145 3.930 1.375 ;
        RECT  3.550 1.015 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 1.015 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 1.015 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 1.015 2.590 1.375 ;
        RECT  2.230 1.145 2.470 1.375 ;
        RECT  2.110 1.015 2.230 1.375 ;
        RECT  1.870 1.145 2.110 1.375 ;
        RECT  1.750 1.015 1.870 1.375 ;
        RECT  1.510 1.145 1.750 1.375 ;
        RECT  1.390 1.015 1.510 1.375 ;
        RECT  1.120 1.145 1.390 1.375 ;
        RECT  1.000 0.710 1.120 1.375 ;
        RECT  0.700 1.145 1.000 1.375 ;
        RECT  0.620 0.860 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 1.000 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.715 3.850 0.945 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.465 0.305 3.755 0.465 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.105 0.305 3.395 0.465 ;
        RECT  3.035 0.185 3.105 0.465 ;
        RECT  2.905 0.305 3.035 0.465 ;
        RECT  2.385 0.305 2.415 0.465 ;
        RECT  1.210 0.715 2.415 0.945 ;
        RECT  2.315 0.185 2.385 0.465 ;
        RECT  2.025 0.305 2.315 0.465 ;
        RECT  1.955 0.185 2.025 0.465 ;
        RECT  1.665 0.305 1.955 0.465 ;
        RECT  1.595 0.185 1.665 0.465 ;
        RECT  1.305 0.305 1.595 0.465 ;
        RECT  1.235 0.185 1.305 0.465 ;
        RECT  2.935 0.545 3.795 0.615 ;
        RECT  0.920 0.545 2.385 0.615 ;
        RECT  0.790 0.195 0.920 1.065 ;
        RECT  0.510 0.335 0.790 0.415 ;
        RECT  0.505 0.705 0.790 0.785 ;
        RECT  0.430 0.185 0.510 0.415 ;
        RECT  0.435 0.705 0.505 1.035 ;
        RECT  0.125 0.845 0.435 0.925 ;
        RECT  0.130 0.335 0.430 0.415 ;
        RECT  0.050 0.245 0.130 0.415 ;
        RECT  0.055 0.845 0.125 0.965 ;
    END
END BUFFD16BWP

MACRO BUFFD1BWP
    CLASS CORE ;
    FOREIGN BUFFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 1.045 ;
        RECT  0.435 0.185 0.455 0.465 ;
        RECT  0.435 0.735 0.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.355 0.520 0.385 0.640 ;
        RECT  0.285 0.335 0.355 0.925 ;
        RECT  0.130 0.335 0.285 0.405 ;
        RECT  0.130 0.855 0.285 0.925 ;
        RECT  0.050 0.205 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END BUFFD1BWP

MACRO BUFFD20BWP
    CLASS CORE ;
    FOREIGN BUFFD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.0080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.730 4.690 0.960 ;
        RECT  4.595 0.185 4.665 0.465 ;
        RECT  4.305 0.305 4.595 0.465 ;
        RECT  4.235 0.185 4.305 0.465 ;
        RECT  3.945 0.305 4.235 0.465 ;
        RECT  3.875 0.185 3.945 0.465 ;
        RECT  3.585 0.305 3.875 0.465 ;
        RECT  3.515 0.185 3.585 0.465 ;
        RECT  3.255 0.305 3.515 0.465 ;
        RECT  3.225 0.305 3.255 0.960 ;
        RECT  3.155 0.185 3.225 0.960 ;
        RECT  2.905 0.305 3.155 0.960 ;
        RECT  2.865 0.305 2.905 0.465 ;
        RECT  1.330 0.730 2.905 0.960 ;
        RECT  2.795 0.185 2.865 0.465 ;
        RECT  2.505 0.305 2.795 0.465 ;
        RECT  2.435 0.185 2.505 0.465 ;
        RECT  2.145 0.305 2.435 0.465 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.305 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.305 1.715 0.465 ;
        RECT  1.355 0.185 1.425 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.665 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.115 4.900 0.115 ;
        RECT  4.770 -0.115 4.850 0.465 ;
        RECT  4.510 -0.115 4.770 0.115 ;
        RECT  4.390 -0.115 4.510 0.235 ;
        RECT  4.150 -0.115 4.390 0.115 ;
        RECT  4.030 -0.115 4.150 0.235 ;
        RECT  3.790 -0.115 4.030 0.115 ;
        RECT  3.670 -0.115 3.790 0.235 ;
        RECT  3.430 -0.115 3.670 0.115 ;
        RECT  3.310 -0.115 3.430 0.235 ;
        RECT  3.070 -0.115 3.310 0.115 ;
        RECT  2.950 -0.115 3.070 0.235 ;
        RECT  2.710 -0.115 2.950 0.115 ;
        RECT  2.590 -0.115 2.710 0.235 ;
        RECT  2.350 -0.115 2.590 0.115 ;
        RECT  2.230 -0.115 2.350 0.235 ;
        RECT  1.990 -0.115 2.230 0.115 ;
        RECT  1.870 -0.115 1.990 0.235 ;
        RECT  1.630 -0.115 1.870 0.115 ;
        RECT  1.510 -0.115 1.630 0.235 ;
        RECT  1.245 -0.115 1.510 0.115 ;
        RECT  1.175 -0.115 1.245 0.465 ;
        RECT  0.875 -0.115 1.175 0.115 ;
        RECT  0.805 -0.115 0.875 0.255 ;
        RECT  0.495 -0.115 0.805 0.115 ;
        RECT  0.425 -0.115 0.495 0.255 ;
        RECT  0.130 -0.115 0.425 0.115 ;
        RECT  0.050 -0.115 0.130 0.410 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.145 4.900 1.375 ;
        RECT  4.770 0.680 4.850 1.375 ;
        RECT  4.510 1.145 4.770 1.375 ;
        RECT  4.390 1.030 4.510 1.375 ;
        RECT  4.150 1.145 4.390 1.375 ;
        RECT  4.030 1.030 4.150 1.375 ;
        RECT  3.790 1.145 4.030 1.375 ;
        RECT  3.670 1.030 3.790 1.375 ;
        RECT  3.430 1.145 3.670 1.375 ;
        RECT  3.310 1.030 3.430 1.375 ;
        RECT  3.070 1.145 3.310 1.375 ;
        RECT  2.950 1.030 3.070 1.375 ;
        RECT  2.710 1.145 2.950 1.375 ;
        RECT  2.590 1.030 2.710 1.375 ;
        RECT  2.350 1.145 2.590 1.375 ;
        RECT  2.230 1.030 2.350 1.375 ;
        RECT  1.990 1.145 2.230 1.375 ;
        RECT  1.870 1.030 1.990 1.375 ;
        RECT  1.630 1.145 1.870 1.375 ;
        RECT  1.510 1.030 1.630 1.375 ;
        RECT  1.245 1.145 1.510 1.375 ;
        RECT  1.175 0.720 1.245 1.375 ;
        RECT  0.875 1.145 1.175 1.375 ;
        RECT  0.805 0.860 0.875 1.375 ;
        RECT  0.510 1.145 0.805 1.375 ;
        RECT  0.410 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.325 0.730 4.690 0.960 ;
        RECT  4.595 0.185 4.665 0.465 ;
        RECT  4.305 0.305 4.595 0.465 ;
        RECT  4.235 0.185 4.305 0.465 ;
        RECT  3.945 0.305 4.235 0.465 ;
        RECT  3.875 0.185 3.945 0.465 ;
        RECT  3.585 0.305 3.875 0.465 ;
        RECT  3.515 0.185 3.585 0.465 ;
        RECT  3.325 0.305 3.515 0.465 ;
        RECT  2.795 0.185 2.835 0.465 ;
        RECT  1.330 0.730 2.835 0.960 ;
        RECT  2.505 0.305 2.795 0.465 ;
        RECT  2.435 0.185 2.505 0.465 ;
        RECT  2.145 0.305 2.435 0.465 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.305 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.305 1.715 0.465 ;
        RECT  1.355 0.185 1.425 0.465 ;
        RECT  3.355 0.545 4.575 0.615 ;
        RECT  1.105 0.545 2.805 0.615 ;
        RECT  0.945 0.185 1.105 1.065 ;
        RECT  0.685 0.335 0.945 0.415 ;
        RECT  0.710 0.700 0.945 0.780 ;
        RECT  0.590 0.700 0.710 1.065 ;
        RECT  0.615 0.185 0.685 0.415 ;
        RECT  0.330 0.335 0.615 0.415 ;
        RECT  0.305 0.845 0.590 0.925 ;
        RECT  0.210 0.205 0.330 0.415 ;
        RECT  0.235 0.845 0.305 0.985 ;
    END
END BUFFD20BWP

MACRO BUFFD24BWP
    CLASS CORE ;
    FOREIGN BUFFD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.2096 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.715 5.670 0.945 ;
        RECT  5.575 0.185 5.645 0.465 ;
        RECT  5.285 0.305 5.575 0.465 ;
        RECT  5.215 0.185 5.285 0.465 ;
        RECT  4.925 0.305 5.215 0.465 ;
        RECT  4.855 0.185 4.925 0.465 ;
        RECT  4.565 0.305 4.855 0.465 ;
        RECT  4.495 0.185 4.565 0.465 ;
        RECT  4.205 0.305 4.495 0.465 ;
        RECT  4.135 0.185 4.205 0.465 ;
        RECT  3.845 0.305 4.135 0.465 ;
        RECT  3.815 0.185 3.845 0.465 ;
        RECT  3.775 0.185 3.815 0.945 ;
        RECT  3.485 0.305 3.775 0.945 ;
        RECT  3.465 0.185 3.485 0.945 ;
        RECT  3.415 0.185 3.465 0.465 ;
        RECT  1.590 0.715 3.465 0.945 ;
        RECT  3.125 0.305 3.415 0.465 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  2.765 0.305 3.055 0.465 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.405 0.305 2.695 0.465 ;
        RECT  2.335 0.185 2.405 0.465 ;
        RECT  2.045 0.305 2.335 0.465 ;
        RECT  1.975 0.185 2.045 0.465 ;
        RECT  1.685 0.305 1.975 0.465 ;
        RECT  1.615 0.185 1.685 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2016 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.945 0.625 ;
        RECT  0.175 0.495 0.245 0.760 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 -0.115 5.880 0.115 ;
        RECT  5.750 -0.115 5.830 0.475 ;
        RECT  5.490 -0.115 5.750 0.115 ;
        RECT  5.370 -0.115 5.490 0.235 ;
        RECT  5.130 -0.115 5.370 0.115 ;
        RECT  5.010 -0.115 5.130 0.235 ;
        RECT  4.770 -0.115 5.010 0.115 ;
        RECT  4.650 -0.115 4.770 0.235 ;
        RECT  4.410 -0.115 4.650 0.115 ;
        RECT  4.290 -0.115 4.410 0.235 ;
        RECT  4.050 -0.115 4.290 0.115 ;
        RECT  3.930 -0.115 4.050 0.235 ;
        RECT  3.690 -0.115 3.930 0.115 ;
        RECT  3.570 -0.115 3.690 0.235 ;
        RECT  3.330 -0.115 3.570 0.115 ;
        RECT  3.210 -0.115 3.330 0.235 ;
        RECT  2.970 -0.115 3.210 0.115 ;
        RECT  2.850 -0.115 2.970 0.235 ;
        RECT  2.610 -0.115 2.850 0.115 ;
        RECT  2.490 -0.115 2.610 0.235 ;
        RECT  2.250 -0.115 2.490 0.115 ;
        RECT  2.130 -0.115 2.250 0.235 ;
        RECT  1.890 -0.115 2.130 0.115 ;
        RECT  1.770 -0.115 1.890 0.235 ;
        RECT  1.480 -0.115 1.770 0.115 ;
        RECT  1.400 -0.115 1.480 0.465 ;
        RECT  1.075 -0.115 1.400 0.115 ;
        RECT  1.005 -0.115 1.075 0.245 ;
        RECT  0.695 -0.115 1.005 0.115 ;
        RECT  0.625 -0.115 0.695 0.245 ;
        RECT  0.315 -0.115 0.625 0.115 ;
        RECT  0.245 -0.115 0.315 0.245 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.145 5.880 1.375 ;
        RECT  5.750 0.680 5.830 1.375 ;
        RECT  5.490 1.145 5.750 1.375 ;
        RECT  5.370 1.015 5.490 1.375 ;
        RECT  5.130 1.145 5.370 1.375 ;
        RECT  5.010 1.015 5.130 1.375 ;
        RECT  4.770 1.145 5.010 1.375 ;
        RECT  4.650 1.015 4.770 1.375 ;
        RECT  4.410 1.145 4.650 1.375 ;
        RECT  4.290 1.015 4.410 1.375 ;
        RECT  4.050 1.145 4.290 1.375 ;
        RECT  3.930 1.015 4.050 1.375 ;
        RECT  3.690 1.145 3.930 1.375 ;
        RECT  3.570 1.015 3.690 1.375 ;
        RECT  3.330 1.145 3.570 1.375 ;
        RECT  3.210 1.015 3.330 1.375 ;
        RECT  2.970 1.145 3.210 1.375 ;
        RECT  2.850 1.015 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.015 2.610 1.375 ;
        RECT  2.250 1.145 2.490 1.375 ;
        RECT  2.130 1.015 2.250 1.375 ;
        RECT  1.890 1.145 2.130 1.375 ;
        RECT  1.770 1.015 1.890 1.375 ;
        RECT  1.475 1.145 1.770 1.375 ;
        RECT  1.405 0.740 1.475 1.375 ;
        RECT  1.075 1.145 1.405 1.375 ;
        RECT  1.005 0.880 1.075 1.375 ;
        RECT  0.700 1.145 1.005 1.375 ;
        RECT  0.620 0.880 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 1.020 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.715 5.670 0.945 ;
        RECT  5.575 0.185 5.645 0.465 ;
        RECT  5.285 0.305 5.575 0.465 ;
        RECT  5.215 0.185 5.285 0.465 ;
        RECT  4.925 0.305 5.215 0.465 ;
        RECT  4.855 0.185 4.925 0.465 ;
        RECT  4.565 0.305 4.855 0.465 ;
        RECT  4.495 0.185 4.565 0.465 ;
        RECT  4.205 0.305 4.495 0.465 ;
        RECT  4.135 0.185 4.205 0.465 ;
        RECT  3.885 0.305 4.135 0.465 ;
        RECT  3.125 0.305 3.395 0.465 ;
        RECT  1.590 0.715 3.395 0.945 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  2.765 0.305 3.055 0.465 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.405 0.305 2.695 0.465 ;
        RECT  2.335 0.185 2.405 0.465 ;
        RECT  2.045 0.305 2.335 0.465 ;
        RECT  1.975 0.185 2.045 0.465 ;
        RECT  1.685 0.305 1.975 0.465 ;
        RECT  1.615 0.185 1.685 0.465 ;
        RECT  3.915 0.545 5.675 0.615 ;
        RECT  1.325 0.545 3.365 0.615 ;
        RECT  1.145 0.195 1.325 1.070 ;
        RECT  0.890 0.325 1.145 0.415 ;
        RECT  0.910 0.705 1.145 0.795 ;
        RECT  0.790 0.705 0.910 1.070 ;
        RECT  0.810 0.185 0.890 0.415 ;
        RECT  0.510 0.325 0.810 0.415 ;
        RECT  0.530 0.705 0.790 0.795 ;
        RECT  0.410 0.705 0.530 1.065 ;
        RECT  0.430 0.185 0.510 0.415 ;
        RECT  0.130 0.325 0.430 0.415 ;
        RECT  0.125 0.845 0.410 0.915 ;
        RECT  0.050 0.275 0.130 0.415 ;
        RECT  0.055 0.845 0.125 0.965 ;
    END
END BUFFD24BWP

MACRO BUFFD2BWP
    CLASS CORE ;
    FOREIGN BUFFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.765 ;
        RECT  0.585 0.355 0.595 0.465 ;
        RECT  0.585 0.665 0.595 0.765 ;
        RECT  0.515 0.185 0.585 0.465 ;
        RECT  0.515 0.665 0.585 1.075 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.115 0.840 0.115 ;
        RECT  0.690 -0.115 0.770 0.280 ;
        RECT  0.370 -0.115 0.690 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.145 0.840 1.375 ;
        RECT  0.690 0.840 0.770 1.375 ;
        RECT  0.360 1.145 0.690 1.375 ;
        RECT  0.280 1.000 0.360 1.375 ;
        RECT  0.000 1.145 0.280 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.345 0.435 0.930 ;
        RECT  0.150 0.345 0.365 0.415 ;
        RECT  0.150 0.860 0.365 0.930 ;
        RECT  0.070 0.245 0.150 0.415 ;
        RECT  0.070 0.860 0.150 1.035 ;
    END
END BUFFD2BWP

MACRO BUFFD3BWP
    CLASS CORE ;
    FOREIGN BUFFD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.185 0.945 0.490 ;
        RECT  0.875 0.700 0.945 1.045 ;
        RECT  0.855 0.185 0.875 1.045 ;
        RECT  0.665 0.355 0.855 0.820 ;
        RECT  0.545 0.355 0.665 0.475 ;
        RECT  0.545 0.700 0.665 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.280 ;
        RECT  0.360 -0.115 0.640 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 0.890 0.760 1.375 ;
        RECT  0.360 1.145 0.640 1.375 ;
        RECT  0.240 0.995 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.545 0.355 0.595 0.475 ;
        RECT  0.545 0.700 0.595 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        RECT  0.375 0.545 0.575 0.615 ;
        RECT  0.305 0.345 0.375 0.925 ;
        RECT  0.130 0.345 0.305 0.415 ;
        RECT  0.130 0.855 0.305 0.925 ;
        RECT  0.050 0.245 0.130 0.415 ;
        RECT  0.050 0.855 0.130 1.025 ;
    END
END BUFFD3BWP

MACRO BUFFD4BWP
    CLASS CORE ;
    FOREIGN BUFFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.025 0.465 ;
        RECT  1.015 0.700 1.025 1.045 ;
        RECT  0.955 0.185 1.015 1.045 ;
        RECT  0.805 0.355 0.955 0.820 ;
        RECT  0.665 0.355 0.805 0.465 ;
        RECT  0.665 0.700 0.805 0.820 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.700 0.665 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.475 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.280 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.275 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.680 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.890 0.870 1.375 ;
        RECT  0.500 1.145 0.750 1.375 ;
        RECT  0.400 0.975 0.500 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.465 ;
        RECT  0.665 0.700 0.735 0.820 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.700 0.665 1.045 ;
        RECT  0.525 0.545 0.705 0.615 ;
        RECT  0.450 0.345 0.525 0.905 ;
        RECT  0.305 0.345 0.450 0.415 ;
        RECT  0.305 0.835 0.450 0.905 ;
        RECT  0.235 0.245 0.305 0.415 ;
        RECT  0.235 0.835 0.305 0.995 ;
    END
END BUFFD4BWP

MACRO BUFFD6BWP
    CLASS CORE ;
    FOREIGN BUFFD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3024 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.700 1.445 1.045 ;
        RECT  1.155 0.355 1.375 0.465 ;
        RECT  1.155 0.700 1.375 0.820 ;
        RECT  1.085 0.355 1.155 0.820 ;
        RECT  1.065 0.355 1.085 1.045 ;
        RECT  0.995 0.185 1.065 1.045 ;
        RECT  0.945 0.355 0.995 0.820 ;
        RECT  0.685 0.355 0.945 0.465 ;
        RECT  0.685 0.700 0.945 0.820 ;
        RECT  0.615 0.185 0.685 0.465 ;
        RECT  0.615 0.700 0.685 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.465 ;
        RECT  1.280 -0.115 1.550 0.115 ;
        RECT  1.160 -0.115 1.280 0.280 ;
        RECT  0.900 -0.115 1.160 0.115 ;
        RECT  0.780 -0.115 0.900 0.280 ;
        RECT  0.500 -0.115 0.780 0.115 ;
        RECT  0.420 -0.115 0.500 0.270 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.735 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 0.890 1.280 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.780 0.890 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 1.000 0.520 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.700 1.445 1.045 ;
        RECT  1.225 0.355 1.375 0.465 ;
        RECT  1.225 0.700 1.375 0.820 ;
        RECT  0.685 0.355 0.875 0.465 ;
        RECT  0.685 0.700 0.875 0.820 ;
        RECT  0.615 0.185 0.685 0.465 ;
        RECT  0.615 0.700 0.685 1.045 ;
        RECT  1.245 0.540 1.535 0.620 ;
        RECT  0.525 0.545 0.855 0.615 ;
        RECT  0.445 0.345 0.525 0.915 ;
        RECT  0.305 0.345 0.445 0.415 ;
        RECT  0.305 0.845 0.445 0.915 ;
        RECT  0.235 0.245 0.305 0.415 ;
        RECT  0.235 0.845 0.305 0.995 ;
    END
END BUFFD6BWP

MACRO BUFFD8BWP
    CLASS CORE ;
    FOREIGN BUFFD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.720 2.035 0.950 ;
        RECT  1.935 0.185 2.005 0.465 ;
        RECT  1.645 0.305 1.935 0.465 ;
        RECT  1.575 0.185 1.645 0.465 ;
        RECT  1.555 0.185 1.575 0.950 ;
        RECT  1.245 0.305 1.555 0.950 ;
        RECT  1.225 0.185 1.245 0.950 ;
        RECT  1.155 0.185 1.225 0.465 ;
        RECT  0.765 0.720 1.225 0.950 ;
        RECT  0.865 0.305 1.155 0.465 ;
        RECT  0.795 0.185 0.865 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.260 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.465 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.720 -0.115 1.840 0.235 ;
        RECT  1.460 -0.115 1.720 0.115 ;
        RECT  1.340 -0.115 1.460 0.235 ;
        RECT  1.080 -0.115 1.340 0.115 ;
        RECT  0.960 -0.115 1.080 0.235 ;
        RECT  0.690 -0.115 0.960 0.115 ;
        RECT  0.610 -0.115 0.690 0.465 ;
        RECT  0.340 -0.115 0.610 0.115 ;
        RECT  0.220 -0.115 0.340 0.255 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.680 2.190 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.720 1.020 1.840 1.375 ;
        RECT  1.460 1.145 1.720 1.375 ;
        RECT  1.340 1.020 1.460 1.375 ;
        RECT  1.080 1.145 1.340 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.690 1.145 0.960 1.375 ;
        RECT  0.610 0.700 0.690 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.015 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.720 2.035 0.950 ;
        RECT  1.935 0.185 2.005 0.465 ;
        RECT  1.645 0.305 1.935 0.465 ;
        RECT  0.865 0.305 1.155 0.465 ;
        RECT  0.765 0.720 1.155 0.950 ;
        RECT  0.795 0.185 0.865 0.465 ;
        RECT  1.685 0.540 1.985 0.620 ;
        RECT  0.515 0.545 1.135 0.615 ;
        RECT  0.425 0.185 0.515 1.055 ;
        RECT  0.125 0.335 0.425 0.415 ;
        RECT  0.125 0.850 0.425 0.930 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.850 0.125 1.035 ;
    END
END BUFFD8BWP

MACRO BUFTD0BWP
    CLASS CORE ;
    FOREIGN BUFTD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.215 1.505 1.045 ;
        RECT  1.420 0.215 1.435 0.370 ;
        RECT  1.410 0.895 1.435 1.045 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.490 1.050 0.775 ;
        RECT  0.880 0.705 0.980 0.775 ;
        RECT  0.810 0.705 0.880 1.045 ;
        RECT  0.385 0.975 0.810 1.045 ;
        RECT  0.315 0.710 0.385 1.045 ;
        RECT  0.265 0.710 0.315 0.780 ;
        RECT  0.175 0.520 0.265 0.780 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.670 0.540 0.735 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.115 1.540 0.115 ;
        RECT  1.170 -0.115 1.290 0.125 ;
        RECT  0.750 -0.115 1.170 0.115 ;
        RECT  0.630 -0.115 0.750 0.130 ;
        RECT  0.315 -0.115 0.630 0.115 ;
        RECT  0.245 -0.115 0.315 0.305 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 1.005 1.300 1.375 ;
        RECT  0.870 1.145 1.180 1.375 ;
        RECT  0.750 1.130 0.870 1.375 ;
        RECT  0.360 1.145 0.750 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.685 1.355 0.805 ;
        RECT  1.280 0.205 1.350 0.605 ;
        RECT  0.585 0.205 1.280 0.275 ;
        RECT  1.130 0.350 1.200 0.925 ;
        RECT  1.030 0.350 1.130 0.420 ;
        RECT  1.070 0.850 1.130 0.925 ;
        RECT  0.990 0.850 1.070 1.055 ;
        RECT  0.585 0.805 0.710 0.875 ;
        RECT  0.515 0.205 0.585 0.875 ;
        RECT  0.410 0.205 0.515 0.275 ;
        RECT  0.365 0.380 0.435 0.640 ;
        RECT  0.125 0.380 0.365 0.450 ;
        RECT  0.105 0.850 0.130 0.970 ;
        RECT  0.105 0.210 0.125 0.450 ;
        RECT  0.035 0.210 0.105 0.970 ;
        RECT  1.350 0.485 1.365 0.605 ;
    END
END BUFTD0BWP

MACRO BUFTD12BWP
    CLASS CORE ;
    FOREIGN BUFTD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5516 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.185 3.825 0.485 ;
        RECT  3.755 0.775 3.825 1.070 ;
        RECT  3.465 0.335 3.755 0.485 ;
        RECT  3.465 0.775 3.755 0.925 ;
        RECT  3.395 0.185 3.465 0.485 ;
        RECT  3.395 0.775 3.465 1.070 ;
        RECT  3.105 0.335 3.395 0.485 ;
        RECT  3.105 0.775 3.395 0.925 ;
        RECT  3.035 0.185 3.105 0.485 ;
        RECT  3.035 0.775 3.105 1.070 ;
        RECT  2.975 0.335 3.035 0.485 ;
        RECT  2.975 0.775 3.035 0.925 ;
        RECT  2.765 0.335 2.975 0.925 ;
        RECT  2.745 0.335 2.765 0.485 ;
        RECT  2.745 0.775 2.765 0.925 ;
        RECT  2.675 0.185 2.745 0.485 ;
        RECT  2.675 0.775 2.745 1.070 ;
        RECT  2.390 0.335 2.675 0.485 ;
        RECT  2.385 0.775 2.675 0.925 ;
        RECT  2.270 0.215 2.390 0.485 ;
        RECT  2.315 0.775 2.385 1.070 ;
        RECT  2.025 0.775 2.315 0.925 ;
        RECT  1.915 0.215 2.270 0.345 ;
        RECT  1.955 0.775 2.025 1.070 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.520 1.505 0.780 ;
        RECT  1.085 0.710 1.425 0.780 ;
        RECT  1.015 0.710 1.085 0.940 ;
        RECT  0.390 0.870 1.015 0.940 ;
        RECT  0.315 0.495 0.390 0.940 ;
        RECT  0.175 0.495 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1064 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.170 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.430 ;
        RECT  3.670 -0.115 3.935 0.115 ;
        RECT  3.550 -0.115 3.670 0.250 ;
        RECT  3.310 -0.115 3.550 0.115 ;
        RECT  3.190 -0.115 3.310 0.250 ;
        RECT  2.950 -0.115 3.190 0.115 ;
        RECT  2.830 -0.115 2.950 0.250 ;
        RECT  2.580 -0.115 2.830 0.115 ;
        RECT  2.460 -0.115 2.580 0.250 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.145 ;
        RECT  1.820 -0.115 2.080 0.115 ;
        RECT  1.700 -0.115 1.820 0.140 ;
        RECT  1.090 -0.115 1.700 0.115 ;
        RECT  0.970 -0.115 1.090 0.250 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.330 -0.115 0.600 0.115 ;
        RECT  0.230 -0.115 0.330 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.145 4.060 1.375 ;
        RECT  3.935 0.720 4.005 1.375 ;
        RECT  3.670 1.145 3.935 1.375 ;
        RECT  3.550 0.995 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 0.995 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 0.995 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 0.995 2.590 1.375 ;
        RECT  2.230 1.145 2.470 1.375 ;
        RECT  2.110 0.995 2.230 1.375 ;
        RECT  1.845 1.145 2.110 1.375 ;
        RECT  1.775 0.790 1.845 1.375 ;
        RECT  1.480 1.145 1.775 1.375 ;
        RECT  1.360 0.990 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.010 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.755 0.185 3.825 0.485 ;
        RECT  3.755 0.775 3.825 1.070 ;
        RECT  3.465 0.335 3.755 0.485 ;
        RECT  3.465 0.775 3.755 0.925 ;
        RECT  3.395 0.185 3.465 0.485 ;
        RECT  3.395 0.775 3.465 1.070 ;
        RECT  3.105 0.335 3.395 0.485 ;
        RECT  3.105 0.775 3.395 0.925 ;
        RECT  3.045 0.185 3.105 0.485 ;
        RECT  3.045 0.775 3.105 1.070 ;
        RECT  2.675 0.185 2.695 0.485 ;
        RECT  2.675 0.775 2.695 1.070 ;
        RECT  2.390 0.335 2.675 0.485 ;
        RECT  2.385 0.775 2.675 0.925 ;
        RECT  2.270 0.215 2.390 0.485 ;
        RECT  2.315 0.775 2.385 1.070 ;
        RECT  2.025 0.775 2.315 0.925 ;
        RECT  1.915 0.215 2.270 0.345 ;
        RECT  1.955 0.775 2.025 1.070 ;
        RECT  1.645 0.635 2.000 0.705 ;
        RECT  1.815 0.455 1.990 0.525 ;
        RECT  1.745 0.225 1.815 0.525 ;
        RECT  1.250 0.225 1.745 0.295 ;
        RECT  1.575 0.365 1.645 1.070 ;
        RECT  1.330 0.365 1.575 0.435 ;
        RECT  1.170 0.850 1.575 0.920 ;
        RECT  1.180 0.225 1.250 0.390 ;
        RECT  0.885 0.320 1.180 0.390 ;
        RECT  0.805 0.210 0.885 0.390 ;
        RECT  0.735 0.210 0.805 0.800 ;
        RECT  0.410 0.210 0.735 0.280 ;
        RECT  0.610 0.730 0.735 0.800 ;
        RECT  0.585 0.350 0.665 0.640 ;
        RECT  0.130 0.350 0.585 0.420 ;
        RECT  0.105 0.250 0.130 0.420 ;
        RECT  0.105 0.735 0.125 1.040 ;
        RECT  0.035 0.250 0.105 1.040 ;
    END
END BUFTD12BWP

MACRO BUFTD16BWP
    CLASS CORE ;
    FOREIGN BUFTD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7420 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.455 0.185 4.525 0.485 ;
        RECT  4.455 0.775 4.525 1.070 ;
        RECT  4.165 0.335 4.455 0.485 ;
        RECT  4.165 0.775 4.455 0.925 ;
        RECT  4.095 0.185 4.165 0.485 ;
        RECT  4.095 0.775 4.165 1.070 ;
        RECT  3.805 0.335 4.095 0.485 ;
        RECT  3.805 0.775 4.095 0.925 ;
        RECT  3.735 0.185 3.805 0.485 ;
        RECT  3.735 0.775 3.805 1.070 ;
        RECT  3.445 0.335 3.735 0.485 ;
        RECT  3.445 0.775 3.735 0.925 ;
        RECT  3.375 0.185 3.445 0.485 ;
        RECT  3.375 0.775 3.445 1.070 ;
        RECT  3.255 0.335 3.375 0.485 ;
        RECT  3.255 0.775 3.375 0.925 ;
        RECT  3.085 0.335 3.255 0.925 ;
        RECT  3.045 0.185 3.085 1.070 ;
        RECT  3.015 0.185 3.045 0.485 ;
        RECT  3.015 0.775 3.045 1.070 ;
        RECT  2.725 0.335 3.015 0.485 ;
        RECT  2.725 0.775 3.015 0.925 ;
        RECT  2.655 0.185 2.725 0.485 ;
        RECT  2.655 0.775 2.725 1.070 ;
        RECT  2.390 0.335 2.655 0.485 ;
        RECT  2.365 0.775 2.655 0.925 ;
        RECT  2.270 0.215 2.390 0.485 ;
        RECT  2.295 0.775 2.365 1.070 ;
        RECT  2.005 0.775 2.295 0.925 ;
        RECT  1.915 0.215 2.270 0.345 ;
        RECT  1.935 0.775 2.005 1.070 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.520 1.505 0.780 ;
        RECT  1.085 0.710 1.425 0.780 ;
        RECT  1.015 0.710 1.085 0.935 ;
        RECT  0.390 0.865 1.015 0.935 ;
        RECT  0.315 0.495 0.390 0.935 ;
        RECT  0.175 0.495 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1064 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.495 1.170 0.625 ;
        RECT  0.840 0.495 0.910 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 -0.115 4.760 0.115 ;
        RECT  4.635 -0.115 4.705 0.420 ;
        RECT  4.370 -0.115 4.635 0.115 ;
        RECT  4.250 -0.115 4.370 0.255 ;
        RECT  4.010 -0.115 4.250 0.115 ;
        RECT  3.890 -0.115 4.010 0.255 ;
        RECT  3.650 -0.115 3.890 0.115 ;
        RECT  3.530 -0.115 3.650 0.255 ;
        RECT  3.290 -0.115 3.530 0.115 ;
        RECT  3.170 -0.115 3.290 0.255 ;
        RECT  2.930 -0.115 3.170 0.115 ;
        RECT  2.810 -0.115 2.930 0.255 ;
        RECT  2.560 -0.115 2.810 0.115 ;
        RECT  2.460 -0.115 2.560 0.260 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.145 ;
        RECT  1.820 -0.115 2.080 0.115 ;
        RECT  1.700 -0.115 1.820 0.140 ;
        RECT  1.090 -0.115 1.700 0.115 ;
        RECT  0.970 -0.115 1.090 0.250 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.315 -0.115 0.600 0.115 ;
        RECT  0.245 -0.115 0.315 0.280 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 1.145 4.760 1.375 ;
        RECT  4.635 0.720 4.705 1.375 ;
        RECT  4.370 1.145 4.635 1.375 ;
        RECT  4.250 0.995 4.370 1.375 ;
        RECT  4.010 1.145 4.250 1.375 ;
        RECT  3.890 0.995 4.010 1.375 ;
        RECT  3.650 1.145 3.890 1.375 ;
        RECT  3.530 0.995 3.650 1.375 ;
        RECT  3.290 1.145 3.530 1.375 ;
        RECT  3.170 0.995 3.290 1.375 ;
        RECT  2.930 1.145 3.170 1.375 ;
        RECT  2.810 0.995 2.930 1.375 ;
        RECT  2.570 1.145 2.810 1.375 ;
        RECT  2.450 0.995 2.570 1.375 ;
        RECT  2.210 1.145 2.450 1.375 ;
        RECT  2.090 0.995 2.210 1.375 ;
        RECT  1.825 1.145 2.090 1.375 ;
        RECT  1.755 0.790 1.825 1.375 ;
        RECT  1.480 1.145 1.755 1.375 ;
        RECT  1.360 0.990 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.010 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 1.005 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.455 0.185 4.525 0.485 ;
        RECT  4.455 0.775 4.525 1.070 ;
        RECT  4.165 0.335 4.455 0.485 ;
        RECT  4.165 0.775 4.455 0.925 ;
        RECT  4.095 0.185 4.165 0.485 ;
        RECT  4.095 0.775 4.165 1.070 ;
        RECT  3.805 0.335 4.095 0.485 ;
        RECT  3.805 0.775 4.095 0.925 ;
        RECT  3.735 0.185 3.805 0.485 ;
        RECT  3.735 0.775 3.805 1.070 ;
        RECT  3.445 0.335 3.735 0.485 ;
        RECT  3.445 0.775 3.735 0.925 ;
        RECT  3.375 0.185 3.445 0.485 ;
        RECT  3.375 0.775 3.445 1.070 ;
        RECT  3.325 0.335 3.375 0.485 ;
        RECT  3.325 0.775 3.375 0.925 ;
        RECT  2.725 0.335 2.975 0.485 ;
        RECT  2.725 0.775 2.975 0.925 ;
        RECT  2.655 0.185 2.725 0.485 ;
        RECT  2.655 0.775 2.725 1.070 ;
        RECT  2.390 0.335 2.655 0.485 ;
        RECT  2.365 0.775 2.655 0.925 ;
        RECT  2.270 0.215 2.390 0.485 ;
        RECT  2.295 0.775 2.365 1.070 ;
        RECT  2.005 0.775 2.295 0.925 ;
        RECT  1.915 0.215 2.270 0.345 ;
        RECT  1.935 0.775 2.005 1.070 ;
        RECT  1.815 0.455 2.000 0.525 ;
        RECT  1.645 0.635 2.000 0.705 ;
        RECT  1.745 0.225 1.815 0.525 ;
        RECT  1.250 0.225 1.745 0.295 ;
        RECT  1.575 0.365 1.645 1.070 ;
        RECT  1.330 0.365 1.575 0.435 ;
        RECT  1.170 0.850 1.575 0.920 ;
        RECT  1.180 0.225 1.250 0.390 ;
        RECT  0.885 0.320 1.180 0.390 ;
        RECT  0.770 0.210 0.885 0.390 ;
        RECT  0.700 0.210 0.770 0.795 ;
        RECT  0.400 0.210 0.700 0.280 ;
        RECT  0.610 0.725 0.700 0.795 ;
        RECT  0.550 0.350 0.630 0.640 ;
        RECT  0.130 0.350 0.550 0.420 ;
        RECT  0.105 0.250 0.130 0.420 ;
        RECT  0.105 0.735 0.125 1.040 ;
        RECT  0.035 0.250 0.105 1.040 ;
    END
END BUFTD16BWP

MACRO BUFTD1BWP
    CLASS CORE ;
    FOREIGN BUFTD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0702 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.215 1.505 1.045 ;
        RECT  1.420 0.215 1.435 0.370 ;
        RECT  1.390 0.900 1.435 1.045 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0528 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.490 0.995 0.610 ;
        RECT  0.875 0.490 0.945 0.940 ;
        RECT  0.505 0.870 0.875 0.940 ;
        RECT  0.435 0.710 0.505 0.940 ;
        RECT  0.265 0.710 0.435 0.780 ;
        RECT  0.175 0.520 0.265 0.780 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0528 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.355 0.805 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.540 0.115 ;
        RECT  1.190 -0.115 1.310 0.130 ;
        RECT  0.740 -0.115 1.190 0.115 ;
        RECT  0.620 -0.115 0.740 0.130 ;
        RECT  0.315 -0.115 0.620 0.115 ;
        RECT  0.245 -0.115 0.315 0.305 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 1.005 1.300 1.375 ;
        RECT  0.930 1.145 1.180 1.375 ;
        RECT  0.810 1.010 0.930 1.375 ;
        RECT  0.330 1.145 0.810 1.375 ;
        RECT  0.250 0.860 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.460 1.365 0.580 ;
        RECT  1.180 0.650 1.355 0.770 ;
        RECT  1.260 0.200 1.330 0.580 ;
        RECT  0.645 0.200 1.260 0.270 ;
        RECT  1.110 0.350 1.180 0.925 ;
        RECT  1.010 0.350 1.110 0.420 ;
        RECT  1.090 0.850 1.110 0.925 ;
        RECT  1.020 0.850 1.090 1.040 ;
        RECT  0.645 0.720 0.710 0.790 ;
        RECT  0.575 0.200 0.645 0.790 ;
        RECT  0.410 0.200 0.575 0.270 ;
        RECT  0.365 0.380 0.435 0.640 ;
        RECT  0.125 0.380 0.365 0.450 ;
        RECT  0.105 0.850 0.130 0.970 ;
        RECT  0.105 0.245 0.125 0.450 ;
        RECT  0.035 0.245 0.105 0.970 ;
    END
END BUFTD1BWP

MACRO BUFTD20BWP
    CLASS CORE ;
    FOREIGN BUFTD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.9438 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.275 0.185 6.345 0.465 ;
        RECT  6.275 0.720 6.345 1.070 ;
        RECT  5.985 0.345 6.275 0.465 ;
        RECT  5.985 0.720 6.275 0.840 ;
        RECT  5.915 0.185 5.985 0.465 ;
        RECT  5.915 0.720 5.985 1.070 ;
        RECT  5.625 0.345 5.915 0.465 ;
        RECT  5.625 0.720 5.915 0.840 ;
        RECT  5.555 0.185 5.625 0.465 ;
        RECT  5.555 0.720 5.625 1.070 ;
        RECT  5.265 0.345 5.555 0.465 ;
        RECT  5.265 0.720 5.555 0.840 ;
        RECT  5.195 0.185 5.265 0.465 ;
        RECT  5.195 0.720 5.265 1.070 ;
        RECT  4.905 0.345 5.195 0.465 ;
        RECT  4.905 0.720 5.195 0.840 ;
        RECT  4.835 0.185 4.905 0.465 ;
        RECT  4.835 0.720 4.905 1.070 ;
        RECT  4.545 0.345 4.835 0.465 ;
        RECT  4.545 0.720 4.835 0.840 ;
        RECT  4.515 0.185 4.545 0.465 ;
        RECT  4.515 0.720 4.545 1.070 ;
        RECT  4.475 0.185 4.515 1.070 ;
        RECT  4.305 0.345 4.475 0.840 ;
        RECT  4.185 0.345 4.305 0.465 ;
        RECT  4.185 0.720 4.305 0.840 ;
        RECT  4.115 0.185 4.185 0.465 ;
        RECT  4.115 0.720 4.185 1.070 ;
        RECT  3.825 0.345 4.115 0.465 ;
        RECT  3.825 0.720 4.115 0.840 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.755 0.720 3.825 1.070 ;
        RECT  3.465 0.345 3.755 0.465 ;
        RECT  3.465 0.720 3.755 0.840 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.720 3.465 1.070 ;
        RECT  3.090 0.345 3.395 0.465 ;
        RECT  3.105 0.720 3.395 0.840 ;
        RECT  3.035 0.720 3.105 1.070 ;
        RECT  3.010 0.210 3.090 0.465 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.495 2.630 0.915 ;
        RECT  1.930 0.845 2.550 0.915 ;
        RECT  1.850 0.495 1.930 0.915 ;
        RECT  1.630 0.845 1.850 0.915 ;
        RECT  1.560 0.845 1.630 1.050 ;
        RECT  0.390 0.980 1.560 1.050 ;
        RECT  0.315 0.495 0.390 1.050 ;
        RECT  0.175 0.495 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1640 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.345 0.625 ;
        RECT  2.135 0.495 2.215 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 -0.115 6.580 0.115 ;
        RECT  6.455 -0.115 6.525 0.420 ;
        RECT  6.190 -0.115 6.455 0.115 ;
        RECT  6.070 -0.115 6.190 0.255 ;
        RECT  5.830 -0.115 6.070 0.115 ;
        RECT  5.710 -0.115 5.830 0.255 ;
        RECT  5.470 -0.115 5.710 0.115 ;
        RECT  5.350 -0.115 5.470 0.255 ;
        RECT  5.110 -0.115 5.350 0.115 ;
        RECT  4.990 -0.115 5.110 0.255 ;
        RECT  4.750 -0.115 4.990 0.115 ;
        RECT  4.630 -0.115 4.750 0.255 ;
        RECT  4.390 -0.115 4.630 0.115 ;
        RECT  4.270 -0.115 4.390 0.255 ;
        RECT  4.030 -0.115 4.270 0.115 ;
        RECT  3.910 -0.115 4.030 0.255 ;
        RECT  3.670 -0.115 3.910 0.115 ;
        RECT  3.550 -0.115 3.670 0.255 ;
        RECT  3.300 -0.115 3.550 0.115 ;
        RECT  3.180 -0.115 3.300 0.255 ;
        RECT  2.915 -0.115 3.180 0.115 ;
        RECT  2.795 -0.115 2.915 0.140 ;
        RECT  2.360 -0.115 2.795 0.115 ;
        RECT  2.240 -0.115 2.360 0.140 ;
        RECT  1.520 -0.115 2.240 0.115 ;
        RECT  1.400 -0.115 1.520 0.280 ;
        RECT  1.100 -0.115 1.400 0.115 ;
        RECT  0.980 -0.115 1.100 0.140 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.330 -0.115 0.600 0.115 ;
        RECT  0.230 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.580 1.375 ;
        RECT  6.450 0.720 6.530 1.375 ;
        RECT  6.190 1.145 6.450 1.375 ;
        RECT  6.070 0.910 6.190 1.375 ;
        RECT  5.830 1.145 6.070 1.375 ;
        RECT  5.710 0.910 5.830 1.375 ;
        RECT  5.470 1.145 5.710 1.375 ;
        RECT  5.350 0.910 5.470 1.375 ;
        RECT  5.110 1.145 5.350 1.375 ;
        RECT  4.990 0.910 5.110 1.375 ;
        RECT  4.750 1.145 4.990 1.375 ;
        RECT  4.630 0.910 4.750 1.375 ;
        RECT  4.390 1.145 4.630 1.375 ;
        RECT  4.270 0.910 4.390 1.375 ;
        RECT  4.030 1.145 4.270 1.375 ;
        RECT  3.910 0.910 4.030 1.375 ;
        RECT  3.670 1.145 3.910 1.375 ;
        RECT  3.550 0.910 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 0.910 3.310 1.375 ;
        RECT  2.925 1.145 3.190 1.375 ;
        RECT  2.855 0.790 2.925 1.375 ;
        RECT  1.080 1.145 2.855 1.375 ;
        RECT  0.960 1.120 1.080 1.375 ;
        RECT  0.340 1.145 0.960 1.375 ;
        RECT  0.220 1.120 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.275 0.185 6.345 0.465 ;
        RECT  6.275 0.720 6.345 1.070 ;
        RECT  5.985 0.345 6.275 0.465 ;
        RECT  5.985 0.720 6.275 0.840 ;
        RECT  5.915 0.185 5.985 0.465 ;
        RECT  5.915 0.720 5.985 1.070 ;
        RECT  5.625 0.345 5.915 0.465 ;
        RECT  5.625 0.720 5.915 0.840 ;
        RECT  5.555 0.185 5.625 0.465 ;
        RECT  5.555 0.720 5.625 1.070 ;
        RECT  5.265 0.345 5.555 0.465 ;
        RECT  5.265 0.720 5.555 0.840 ;
        RECT  5.195 0.185 5.265 0.465 ;
        RECT  5.195 0.720 5.265 1.070 ;
        RECT  4.905 0.345 5.195 0.465 ;
        RECT  4.905 0.720 5.195 0.840 ;
        RECT  4.835 0.185 4.905 0.465 ;
        RECT  4.835 0.720 4.905 1.070 ;
        RECT  4.585 0.345 4.835 0.465 ;
        RECT  4.585 0.720 4.835 0.840 ;
        RECT  4.185 0.345 4.235 0.465 ;
        RECT  4.185 0.720 4.235 0.840 ;
        RECT  4.115 0.185 4.185 0.465 ;
        RECT  4.115 0.720 4.185 1.070 ;
        RECT  3.825 0.345 4.115 0.465 ;
        RECT  3.825 0.720 4.115 0.840 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.755 0.720 3.825 1.070 ;
        RECT  1.420 0.350 1.490 0.910 ;
        RECT  1.300 0.350 1.420 0.420 ;
        RECT  0.590 0.840 1.420 0.910 ;
        RECT  1.280 0.520 1.350 0.770 ;
        RECT  1.180 0.210 1.300 0.420 ;
        RECT  0.670 0.700 1.280 0.770 ;
        RECT  0.410 0.210 1.180 0.280 ;
        RECT  1.000 0.355 1.100 0.630 ;
        RECT  0.140 0.355 1.000 0.425 ;
        RECT  0.590 0.520 0.670 0.770 ;
        RECT  0.105 0.185 0.140 0.425 ;
        RECT  0.105 0.765 0.130 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        RECT  3.465 0.345 3.755 0.465 ;
        RECT  3.465 0.720 3.755 0.840 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.720 3.465 1.070 ;
        RECT  3.090 0.345 3.395 0.465 ;
        RECT  3.105 0.720 3.395 0.840 ;
        RECT  3.035 0.720 3.105 1.070 ;
        RECT  3.010 0.210 3.090 0.465 ;
        RECT  2.780 0.635 2.950 0.705 ;
        RECT  2.850 0.210 2.920 0.550 ;
        RECT  1.725 0.210 2.850 0.280 ;
        RECT  2.710 0.355 2.780 1.065 ;
        RECT  1.850 0.355 2.710 0.425 ;
        RECT  1.710 0.995 2.710 1.065 ;
        RECT  1.655 0.210 1.725 0.420 ;
        RECT  1.490 0.350 1.655 0.420 ;
    END
END BUFTD20BWP

MACRO BUFTD24BWP
    CLASS CORE ;
    FOREIGN BUFTD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.1342 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.975 0.185 7.045 0.465 ;
        RECT  6.975 0.710 7.045 1.070 ;
        RECT  6.685 0.345 6.975 0.465 ;
        RECT  6.685 0.710 6.975 0.840 ;
        RECT  6.615 0.185 6.685 0.465 ;
        RECT  6.615 0.710 6.685 1.070 ;
        RECT  6.325 0.345 6.615 0.465 ;
        RECT  6.325 0.710 6.615 0.840 ;
        RECT  6.255 0.185 6.325 0.465 ;
        RECT  6.255 0.710 6.325 1.070 ;
        RECT  5.965 0.345 6.255 0.465 ;
        RECT  5.965 0.710 6.255 0.840 ;
        RECT  5.895 0.185 5.965 0.465 ;
        RECT  5.895 0.710 5.965 1.070 ;
        RECT  5.605 0.345 5.895 0.465 ;
        RECT  5.605 0.710 5.895 0.840 ;
        RECT  5.535 0.185 5.605 0.465 ;
        RECT  5.535 0.710 5.605 1.070 ;
        RECT  5.245 0.345 5.535 0.465 ;
        RECT  5.245 0.710 5.535 0.840 ;
        RECT  5.175 0.185 5.245 0.465 ;
        RECT  5.175 0.710 5.245 1.070 ;
        RECT  4.885 0.345 5.175 0.465 ;
        RECT  4.885 0.710 5.175 0.840 ;
        RECT  4.815 0.185 4.885 0.465 ;
        RECT  4.815 0.710 4.885 1.070 ;
        RECT  4.525 0.345 4.815 0.465 ;
        RECT  4.525 0.710 4.815 0.840 ;
        RECT  4.515 0.185 4.525 0.465 ;
        RECT  4.515 0.710 4.525 1.070 ;
        RECT  4.455 0.185 4.515 1.070 ;
        RECT  4.305 0.345 4.455 0.840 ;
        RECT  4.165 0.345 4.305 0.465 ;
        RECT  4.165 0.720 4.305 0.840 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.720 4.165 1.070 ;
        RECT  3.805 0.345 4.095 0.465 ;
        RECT  3.805 0.720 4.095 0.840 ;
        RECT  3.735 0.185 3.805 0.465 ;
        RECT  3.735 0.720 3.805 1.070 ;
        RECT  3.445 0.345 3.735 0.465 ;
        RECT  3.445 0.720 3.735 0.840 ;
        RECT  3.375 0.185 3.445 0.465 ;
        RECT  3.375 0.720 3.445 1.070 ;
        RECT  3.100 0.345 3.375 0.465 ;
        RECT  3.085 0.720 3.375 0.840 ;
        RECT  3.000 0.220 3.100 0.465 ;
        RECT  3.015 0.720 3.085 1.070 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.1048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.520 2.615 0.915 ;
        RECT  1.930 0.845 2.545 0.915 ;
        RECT  1.855 0.495 1.930 0.915 ;
        RECT  1.630 0.845 1.855 0.915 ;
        RECT  1.560 0.845 1.630 1.050 ;
        RECT  0.390 0.980 1.560 1.050 ;
        RECT  0.315 0.520 0.390 1.050 ;
        RECT  0.175 0.520 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1640 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.345 0.625 ;
        RECT  2.135 0.495 2.215 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.225 -0.115 7.280 0.115 ;
        RECT  7.155 -0.115 7.225 0.430 ;
        RECT  6.890 -0.115 7.155 0.115 ;
        RECT  6.770 -0.115 6.890 0.255 ;
        RECT  6.530 -0.115 6.770 0.115 ;
        RECT  6.410 -0.115 6.530 0.255 ;
        RECT  6.170 -0.115 6.410 0.115 ;
        RECT  6.050 -0.115 6.170 0.255 ;
        RECT  5.810 -0.115 6.050 0.115 ;
        RECT  5.690 -0.115 5.810 0.255 ;
        RECT  5.450 -0.115 5.690 0.115 ;
        RECT  5.330 -0.115 5.450 0.255 ;
        RECT  5.090 -0.115 5.330 0.115 ;
        RECT  4.970 -0.115 5.090 0.255 ;
        RECT  4.730 -0.115 4.970 0.115 ;
        RECT  4.610 -0.115 4.730 0.255 ;
        RECT  4.370 -0.115 4.610 0.115 ;
        RECT  4.250 -0.115 4.370 0.255 ;
        RECT  4.010 -0.115 4.250 0.115 ;
        RECT  3.890 -0.115 4.010 0.255 ;
        RECT  3.650 -0.115 3.890 0.115 ;
        RECT  3.530 -0.115 3.650 0.255 ;
        RECT  3.290 -0.115 3.530 0.115 ;
        RECT  3.170 -0.115 3.290 0.255 ;
        RECT  2.915 -0.115 3.170 0.115 ;
        RECT  2.795 -0.115 2.915 0.140 ;
        RECT  2.360 -0.115 2.795 0.115 ;
        RECT  2.240 -0.115 2.360 0.140 ;
        RECT  1.520 -0.115 2.240 0.115 ;
        RECT  1.400 -0.115 1.520 0.270 ;
        RECT  1.100 -0.115 1.400 0.115 ;
        RECT  0.980 -0.115 1.100 0.140 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.315 -0.115 0.600 0.115 ;
        RECT  0.245 -0.115 0.315 0.300 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.230 1.145 7.280 1.375 ;
        RECT  7.150 0.720 7.230 1.375 ;
        RECT  6.890 1.145 7.150 1.375 ;
        RECT  6.770 0.910 6.890 1.375 ;
        RECT  6.530 1.145 6.770 1.375 ;
        RECT  6.410 0.910 6.530 1.375 ;
        RECT  6.170 1.145 6.410 1.375 ;
        RECT  6.050 0.910 6.170 1.375 ;
        RECT  5.810 1.145 6.050 1.375 ;
        RECT  5.690 0.910 5.810 1.375 ;
        RECT  5.450 1.145 5.690 1.375 ;
        RECT  5.330 0.910 5.450 1.375 ;
        RECT  5.090 1.145 5.330 1.375 ;
        RECT  4.970 0.910 5.090 1.375 ;
        RECT  4.730 1.145 4.970 1.375 ;
        RECT  4.610 0.910 4.730 1.375 ;
        RECT  4.370 1.145 4.610 1.375 ;
        RECT  4.250 0.910 4.370 1.375 ;
        RECT  4.010 1.145 4.250 1.375 ;
        RECT  3.890 0.910 4.010 1.375 ;
        RECT  3.650 1.145 3.890 1.375 ;
        RECT  3.530 0.910 3.650 1.375 ;
        RECT  3.290 1.145 3.530 1.375 ;
        RECT  3.170 0.910 3.290 1.375 ;
        RECT  2.905 1.145 3.170 1.375 ;
        RECT  2.835 0.790 2.905 1.375 ;
        RECT  1.080 1.145 2.835 1.375 ;
        RECT  0.960 1.120 1.080 1.375 ;
        RECT  0.340 1.145 0.960 1.375 ;
        RECT  0.220 1.120 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.975 0.185 7.045 0.465 ;
        RECT  6.975 0.710 7.045 1.070 ;
        RECT  6.685 0.345 6.975 0.465 ;
        RECT  6.685 0.710 6.975 0.840 ;
        RECT  6.615 0.185 6.685 0.465 ;
        RECT  6.615 0.710 6.685 1.070 ;
        RECT  6.325 0.345 6.615 0.465 ;
        RECT  6.325 0.710 6.615 0.840 ;
        RECT  6.255 0.185 6.325 0.465 ;
        RECT  6.255 0.710 6.325 1.070 ;
        RECT  5.965 0.345 6.255 0.465 ;
        RECT  5.965 0.710 6.255 0.840 ;
        RECT  5.895 0.185 5.965 0.465 ;
        RECT  5.895 0.710 5.965 1.070 ;
        RECT  5.605 0.345 5.895 0.465 ;
        RECT  5.605 0.710 5.895 0.840 ;
        RECT  5.535 0.185 5.605 0.465 ;
        RECT  5.535 0.710 5.605 1.070 ;
        RECT  5.245 0.345 5.535 0.465 ;
        RECT  5.245 0.710 5.535 0.840 ;
        RECT  5.175 0.185 5.245 0.465 ;
        RECT  5.175 0.710 5.245 1.070 ;
        RECT  4.885 0.345 5.175 0.465 ;
        RECT  4.885 0.710 5.175 0.840 ;
        RECT  4.815 0.185 4.885 0.465 ;
        RECT  4.815 0.710 4.885 1.070 ;
        RECT  4.585 0.345 4.815 0.465 ;
        RECT  4.585 0.710 4.815 0.840 ;
        RECT  4.165 0.345 4.235 0.465 ;
        RECT  4.165 0.720 4.235 0.840 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.720 4.165 1.070 ;
        RECT  3.805 0.345 4.095 0.465 ;
        RECT  3.805 0.720 4.095 0.840 ;
        RECT  3.735 0.185 3.805 0.465 ;
        RECT  3.735 0.720 3.805 1.070 ;
        RECT  3.445 0.345 3.735 0.465 ;
        RECT  3.445 0.720 3.735 0.840 ;
        RECT  3.375 0.185 3.445 0.465 ;
        RECT  3.375 0.720 3.445 1.070 ;
        RECT  3.100 0.345 3.375 0.465 ;
        RECT  3.085 0.720 3.375 0.840 ;
        RECT  3.000 0.220 3.100 0.465 ;
        RECT  3.015 0.720 3.085 1.070 ;
        RECT  1.180 0.210 1.300 0.420 ;
        RECT  0.670 0.700 1.280 0.770 ;
        RECT  0.410 0.210 1.180 0.280 ;
        RECT  1.000 0.370 1.100 0.630 ;
        RECT  0.125 0.370 1.000 0.440 ;
        RECT  0.590 0.520 0.670 0.770 ;
        RECT  0.105 0.765 0.130 1.045 ;
        RECT  0.105 0.250 0.125 0.440 ;
        RECT  0.035 0.250 0.105 1.045 ;
        RECT  2.755 0.635 2.930 0.705 ;
        RECT  2.825 0.210 2.895 0.550 ;
        RECT  1.735 0.210 2.825 0.280 ;
        RECT  2.685 0.355 2.755 1.065 ;
        RECT  1.850 0.355 2.685 0.425 ;
        RECT  1.710 0.995 2.685 1.065 ;
        RECT  1.665 0.210 1.735 0.420 ;
        RECT  1.490 0.350 1.665 0.420 ;
        RECT  1.420 0.350 1.490 0.910 ;
        RECT  1.300 0.350 1.420 0.420 ;
        RECT  0.590 0.840 1.420 0.910 ;
        RECT  1.280 0.520 1.350 0.770 ;
    END
END BUFTD24BWP

MACRO BUFTD2BWP
    CLASS CORE ;
    FOREIGN BUFTD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0798 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.370 1.645 0.905 ;
        RECT  1.470 0.370 1.575 0.440 ;
        RECT  1.445 0.835 1.575 0.905 ;
        RECT  1.400 0.245 1.470 0.440 ;
        RECT  1.375 0.835 1.445 1.015 ;
        RECT  1.380 0.245 1.400 0.365 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.520 1.020 0.780 ;
        RECT  0.945 0.710 0.950 0.780 ;
        RECT  0.875 0.710 0.945 0.930 ;
        RECT  0.505 0.860 0.875 0.930 ;
        RECT  0.435 0.710 0.505 0.930 ;
        RECT  0.265 0.710 0.435 0.780 ;
        RECT  0.175 0.495 0.265 0.780 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.645 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 -0.115 1.680 0.115 ;
        RECT  1.540 -0.115 1.640 0.300 ;
        RECT  1.275 -0.115 1.540 0.115 ;
        RECT  1.155 -0.115 1.275 0.135 ;
        RECT  0.720 -0.115 1.155 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.285 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.145 1.680 1.375 ;
        RECT  1.540 0.990 1.640 1.375 ;
        RECT  1.270 1.145 1.540 1.375 ;
        RECT  1.190 1.000 1.270 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 1.010 0.930 1.375 ;
        RECT  0.320 1.145 0.810 1.375 ;
        RECT  0.240 0.860 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.090 0.360 1.160 0.930 ;
        RECT  0.960 0.360 1.090 0.430 ;
        RECT  1.085 0.860 1.090 0.930 ;
        RECT  1.015 0.860 1.085 1.060 ;
        RECT  0.645 0.720 0.710 0.790 ;
        RECT  0.575 0.205 0.645 0.790 ;
        RECT  0.410 0.205 0.575 0.275 ;
        RECT  0.365 0.355 0.435 0.640 ;
        RECT  0.125 0.355 0.365 0.425 ;
        RECT  0.105 0.850 0.130 0.970 ;
        RECT  0.105 0.245 0.125 0.425 ;
        RECT  0.035 0.245 0.105 0.970 ;
        RECT  1.160 0.665 1.420 0.735 ;
        RECT  1.310 0.460 1.330 0.580 ;
        RECT  1.240 0.205 1.310 0.580 ;
        RECT  0.645 0.205 1.240 0.275 ;
    END
END BUFTD2BWP

MACRO BUFTD3BWP
    CLASS CORE ;
    FOREIGN BUFTD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1513 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.215 1.905 0.345 ;
        RECT  1.835 0.775 1.905 1.065 ;
        RECT  1.715 0.775 1.835 0.925 ;
        RECT  1.505 0.215 1.715 0.925 ;
        RECT  1.415 0.215 1.505 0.345 ;
        RECT  1.485 0.785 1.505 0.925 ;
        RECT  1.415 0.785 1.485 1.065 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.520 1.020 0.780 ;
        RECT  0.945 0.710 0.950 0.780 ;
        RECT  0.875 0.710 0.945 0.930 ;
        RECT  0.490 0.860 0.875 0.930 ;
        RECT  0.420 0.710 0.490 0.930 ;
        RECT  0.265 0.710 0.420 0.780 ;
        RECT  0.175 0.495 0.265 0.780 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.645 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.115 1.960 0.115 ;
        RECT  1.600 -0.115 1.720 0.145 ;
        RECT  1.315 -0.115 1.600 0.115 ;
        RECT  1.195 -0.115 1.315 0.135 ;
        RECT  0.740 -0.115 1.195 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.315 -0.115 0.620 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.145 1.960 1.375 ;
        RECT  1.600 1.010 1.720 1.375 ;
        RECT  1.310 1.145 1.600 1.375 ;
        RECT  1.240 0.805 1.310 1.375 ;
        RECT  0.930 1.145 1.240 1.375 ;
        RECT  0.810 1.010 0.930 1.375 ;
        RECT  0.320 1.145 0.810 1.375 ;
        RECT  0.240 0.860 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.215 1.905 0.345 ;
        RECT  1.835 0.775 1.905 1.065 ;
        RECT  1.785 0.775 1.835 0.925 ;
        RECT  1.415 0.215 1.435 0.345 ;
        RECT  1.415 0.785 1.435 1.065 ;
        RECT  1.320 0.465 1.410 0.535 ;
        RECT  1.090 0.355 1.095 1.060 ;
        RECT  0.990 0.355 1.090 0.425 ;
        RECT  1.025 0.860 1.090 1.060 ;
        RECT  0.645 0.720 0.710 0.790 ;
        RECT  0.575 0.205 0.645 0.790 ;
        RECT  0.410 0.205 0.575 0.275 ;
        RECT  0.365 0.355 0.435 0.640 ;
        RECT  0.125 0.355 0.365 0.425 ;
        RECT  0.105 0.850 0.130 0.970 ;
        RECT  0.105 0.245 0.125 0.425 ;
        RECT  0.035 0.245 0.105 0.970 ;
        RECT  1.160 0.645 1.410 0.715 ;
        RECT  1.250 0.205 1.320 0.535 ;
        RECT  0.645 0.205 1.250 0.275 ;
        RECT  1.095 0.355 1.160 0.930 ;
    END
END BUFTD3BWP

MACRO BUFTD4BWP
    CLASS CORE ;
    FOREIGN BUFTD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1708 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.215 1.870 0.345 ;
        RECT  1.795 0.775 1.865 1.065 ;
        RECT  1.715 0.775 1.795 0.925 ;
        RECT  1.505 0.215 1.715 0.925 ;
        RECT  1.410 0.215 1.505 0.345 ;
        RECT  1.485 0.785 1.505 0.925 ;
        RECT  1.415 0.785 1.485 1.065 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.520 1.020 0.780 ;
        RECT  0.945 0.710 0.950 0.780 ;
        RECT  0.875 0.710 0.945 0.930 ;
        RECT  0.490 0.860 0.875 0.930 ;
        RECT  0.420 0.710 0.490 0.930 ;
        RECT  0.265 0.710 0.420 0.780 ;
        RECT  0.175 0.495 0.265 0.780 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.645 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.420 ;
        RECT  1.700 -0.115 1.970 0.115 ;
        RECT  1.580 -0.115 1.700 0.145 ;
        RECT  1.315 -0.115 1.580 0.115 ;
        RECT  1.195 -0.115 1.315 0.135 ;
        RECT  0.740 -0.115 1.195 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.315 -0.115 0.620 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.145 2.100 1.375 ;
        RECT  1.975 0.775 2.045 1.375 ;
        RECT  1.700 1.145 1.975 1.375 ;
        RECT  1.580 1.015 1.700 1.375 ;
        RECT  1.310 1.145 1.580 1.375 ;
        RECT  1.240 0.805 1.310 1.375 ;
        RECT  0.930 1.145 1.240 1.375 ;
        RECT  0.810 1.010 0.930 1.375 ;
        RECT  0.320 1.145 0.810 1.375 ;
        RECT  0.240 0.860 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.215 1.870 0.345 ;
        RECT  1.795 0.775 1.865 1.065 ;
        RECT  1.785 0.775 1.795 0.925 ;
        RECT  1.410 0.215 1.435 0.345 ;
        RECT  1.415 0.785 1.435 1.065 ;
        RECT  1.310 0.465 1.410 0.535 ;
        RECT  1.160 0.645 1.410 0.715 ;
        RECT  1.240 0.205 1.310 0.535 ;
        RECT  1.025 0.860 1.090 1.065 ;
        RECT  0.645 0.720 0.710 0.790 ;
        RECT  0.575 0.205 0.645 0.790 ;
        RECT  0.410 0.205 0.575 0.275 ;
        RECT  0.365 0.355 0.435 0.640 ;
        RECT  0.125 0.355 0.365 0.425 ;
        RECT  0.105 0.850 0.130 0.970 ;
        RECT  0.105 0.245 0.125 0.425 ;
        RECT  0.035 0.245 0.105 0.970 ;
        RECT  0.645 0.205 1.240 0.275 ;
        RECT  1.095 0.355 1.160 0.930 ;
        RECT  1.090 0.355 1.095 1.065 ;
        RECT  1.000 0.355 1.090 0.425 ;
    END
END BUFTD4BWP

MACRO BUFTD6BWP
    CLASS CORE ;
    FOREIGN BUFTD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2618 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.195 2.710 0.485 ;
        RECT  2.635 0.775 2.705 1.070 ;
        RECT  2.415 0.300 2.635 0.485 ;
        RECT  2.415 0.775 2.635 0.925 ;
        RECT  2.345 0.300 2.415 0.925 ;
        RECT  2.275 0.195 2.345 1.070 ;
        RECT  2.205 0.300 2.275 0.925 ;
        RECT  1.985 0.300 2.205 0.390 ;
        RECT  1.985 0.775 2.205 0.925 ;
        RECT  1.915 0.215 1.985 0.390 ;
        RECT  1.915 0.775 1.985 1.070 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 0.520 1.380 0.780 ;
        RECT  1.085 0.710 1.300 0.780 ;
        RECT  1.015 0.710 1.085 0.930 ;
        RECT  0.385 0.860 1.015 0.930 ;
        RECT  0.315 0.495 0.385 0.930 ;
        RECT  0.175 0.495 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.055 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.115 2.940 0.115 ;
        RECT  2.815 -0.115 2.885 0.450 ;
        RECT  2.550 -0.115 2.815 0.115 ;
        RECT  2.430 -0.115 2.550 0.230 ;
        RECT  2.190 -0.115 2.430 0.115 ;
        RECT  2.070 -0.115 2.190 0.230 ;
        RECT  1.820 -0.115 2.070 0.115 ;
        RECT  1.700 -0.115 1.820 0.140 ;
        RECT  1.090 -0.115 1.700 0.115 ;
        RECT  0.970 -0.115 1.090 0.250 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.315 -0.115 0.600 0.115 ;
        RECT  0.245 -0.115 0.315 0.280 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.145 2.940 1.375 ;
        RECT  2.815 0.720 2.885 1.375 ;
        RECT  2.550 1.145 2.815 1.375 ;
        RECT  2.430 1.005 2.550 1.375 ;
        RECT  2.190 1.145 2.430 1.375 ;
        RECT  2.070 1.005 2.190 1.375 ;
        RECT  1.785 1.145 2.070 1.375 ;
        RECT  1.715 0.790 1.785 1.375 ;
        RECT  1.450 1.145 1.715 1.375 ;
        RECT  1.330 0.990 1.450 1.375 ;
        RECT  1.090 1.145 1.330 1.375 ;
        RECT  0.970 1.000 1.090 1.375 ;
        RECT  0.330 1.145 0.970 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.635 0.195 2.710 0.485 ;
        RECT  2.635 0.775 2.705 1.070 ;
        RECT  2.485 0.300 2.635 0.485 ;
        RECT  2.485 0.775 2.635 0.925 ;
        RECT  1.985 0.300 2.135 0.390 ;
        RECT  1.985 0.775 2.135 0.925 ;
        RECT  1.915 0.215 1.985 0.390 ;
        RECT  1.915 0.775 1.985 1.070 ;
        RECT  1.800 0.460 2.105 0.530 ;
        RECT  1.605 0.635 1.960 0.705 ;
        RECT  1.730 0.225 1.800 0.530 ;
        RECT  1.240 0.225 1.730 0.295 ;
        RECT  1.535 0.365 1.605 1.070 ;
        RECT  1.330 0.365 1.535 0.435 ;
        RECT  1.260 0.850 1.535 0.920 ;
        RECT  1.160 0.850 1.260 0.950 ;
        RECT  1.170 0.225 1.240 0.390 ;
        RECT  0.805 0.320 1.170 0.390 ;
        RECT  0.735 0.215 0.805 0.790 ;
        RECT  0.410 0.215 0.735 0.285 ;
        RECT  0.580 0.720 0.735 0.790 ;
        RECT  0.565 0.355 0.635 0.640 ;
        RECT  0.130 0.355 0.565 0.425 ;
        RECT  0.035 0.250 0.105 1.045 ;
        RECT  0.105 0.250 0.130 0.425 ;
        RECT  0.105 0.770 0.130 1.045 ;
    END
END BUFTD6BWP

MACRO BUFTD8BWP
    CLASS CORE ;
    FOREIGN BUFTD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3528 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.030 0.220 3.150 0.430 ;
        RECT  3.055 0.775 3.125 1.070 ;
        RECT  2.765 0.775 3.055 0.925 ;
        RECT  2.770 0.290 3.030 0.430 ;
        RECT  2.695 0.220 2.770 0.430 ;
        RECT  2.695 0.775 2.765 1.070 ;
        RECT  2.650 0.220 2.695 0.925 ;
        RECT  2.485 0.290 2.650 0.925 ;
        RECT  2.390 0.290 2.485 0.430 ;
        RECT  2.405 0.775 2.485 0.925 ;
        RECT  2.335 0.775 2.405 1.070 ;
        RECT  2.270 0.220 2.390 0.430 ;
        RECT  2.025 0.775 2.335 0.925 ;
        RECT  1.915 0.220 2.270 0.360 ;
        RECT  1.955 0.775 2.025 1.070 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.0760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.520 1.505 0.775 ;
        RECT  1.090 0.705 1.425 0.775 ;
        RECT  1.020 0.705 1.090 0.935 ;
        RECT  0.390 0.865 1.020 0.935 ;
        RECT  0.315 0.495 0.390 0.935 ;
        RECT  0.175 0.495 0.315 0.640 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.1064 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.170 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.115 3.360 0.115 ;
        RECT  3.235 -0.115 3.305 0.420 ;
        RECT  2.935 -0.115 3.235 0.115 ;
        RECT  2.865 -0.115 2.935 0.180 ;
        RECT  2.555 -0.115 2.865 0.115 ;
        RECT  2.485 -0.115 2.555 0.180 ;
        RECT  2.200 -0.115 2.485 0.115 ;
        RECT  2.080 -0.115 2.200 0.145 ;
        RECT  1.820 -0.115 2.080 0.115 ;
        RECT  1.700 -0.115 1.820 0.140 ;
        RECT  1.090 -0.115 1.700 0.115 ;
        RECT  0.970 -0.115 1.090 0.250 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.315 -0.115 0.600 0.115 ;
        RECT  0.245 -0.115 0.315 0.280 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.145 3.360 1.375 ;
        RECT  3.235 0.720 3.305 1.375 ;
        RECT  2.970 1.145 3.235 1.375 ;
        RECT  2.850 1.005 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.005 2.610 1.375 ;
        RECT  2.240 1.145 2.490 1.375 ;
        RECT  2.120 1.005 2.240 1.375 ;
        RECT  1.835 1.145 2.120 1.375 ;
        RECT  1.765 0.790 1.835 1.375 ;
        RECT  1.480 1.145 1.765 1.375 ;
        RECT  1.360 0.990 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.010 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 1.005 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.030 0.220 3.150 0.430 ;
        RECT  3.055 0.775 3.125 1.070 ;
        RECT  2.765 0.775 3.055 0.925 ;
        RECT  2.770 0.290 3.030 0.430 ;
        RECT  2.765 0.220 2.770 0.430 ;
        RECT  2.390 0.290 2.415 0.430 ;
        RECT  2.405 0.775 2.415 0.925 ;
        RECT  2.335 0.775 2.405 1.070 ;
        RECT  2.270 0.220 2.390 0.430 ;
        RECT  2.025 0.775 2.335 0.925 ;
        RECT  1.915 0.220 2.270 0.360 ;
        RECT  1.955 0.775 2.025 1.070 ;
        RECT  1.645 0.635 2.000 0.705 ;
        RECT  1.815 0.455 1.990 0.525 ;
        RECT  1.745 0.225 1.815 0.525 ;
        RECT  1.250 0.225 1.745 0.295 ;
        RECT  1.575 0.365 1.645 1.070 ;
        RECT  1.330 0.365 1.575 0.435 ;
        RECT  1.170 0.850 1.575 0.920 ;
        RECT  1.180 0.225 1.250 0.390 ;
        RECT  0.885 0.320 1.180 0.390 ;
        RECT  0.805 0.210 0.885 0.390 ;
        RECT  0.735 0.210 0.805 0.795 ;
        RECT  0.400 0.210 0.735 0.280 ;
        RECT  0.610 0.725 0.735 0.795 ;
        RECT  0.590 0.350 0.665 0.640 ;
        RECT  0.130 0.350 0.590 0.420 ;
        RECT  0.105 0.250 0.130 0.420 ;
        RECT  0.105 0.735 0.125 1.040 ;
        RECT  0.035 0.250 0.105 1.040 ;
    END
END BUFTD8BWP

MACRO CKAN2D0BWP
    CLASS CORE ;
    FOREIGN CKAN2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0423 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 1.050 ;
        RECT  0.680 0.215 0.735 0.340 ;
        RECT  0.695 0.910 0.735 1.050 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.990 0.580 1.375 ;
        RECT  0.150 1.145 0.460 1.375 ;
        RECT  0.070 0.950 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.660 0.640 ;
        RECT  0.515 0.205 0.585 0.915 ;
        RECT  0.050 0.205 0.515 0.275 ;
        RECT  0.340 0.845 0.515 0.915 ;
        RECT  0.260 0.845 0.340 1.070 ;
    END
END CKAN2D0BWP

MACRO CKAN2D1BWP
    CLASS CORE ;
    FOREIGN CKAN2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0845 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.200 0.805 1.050 ;
        RECT  0.700 0.200 0.735 0.350 ;
        RECT  0.700 0.750 0.735 1.050 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.355 0.400 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.990 0.580 1.375 ;
        RECT  0.150 1.145 0.460 1.375 ;
        RECT  0.070 0.960 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.645 0.640 ;
        RECT  0.515 0.205 0.585 0.915 ;
        RECT  0.050 0.205 0.515 0.275 ;
        RECT  0.340 0.845 0.515 0.915 ;
        RECT  0.260 0.845 0.340 1.070 ;
    END
END CKAN2D1BWP

MACRO CKAN2D2BWP
    CLASS CORE ;
    FOREIGN CKAN2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0910 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.905 ;
        RECT  0.725 0.355 0.735 0.425 ;
        RECT  0.725 0.780 0.735 0.905 ;
        RECT  0.655 0.245 0.725 0.425 ;
        RECT  0.655 0.780 0.725 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.280 ;
        RECT  0.000 -0.115 0.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.990 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.950 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.545 0.650 0.615 ;
        RECT  0.490 0.205 0.560 0.915 ;
        RECT  0.130 0.205 0.490 0.275 ;
        RECT  0.310 0.845 0.490 0.915 ;
        RECT  0.230 0.845 0.310 1.070 ;
        RECT  0.050 0.205 0.130 0.345 ;
    END
END CKAN2D2BWP

MACRO CKAN2D4BWP
    CLASS CORE ;
    FOREIGN CKAN2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1820 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.245 1.025 0.495 ;
        RECT  1.015 0.720 1.025 1.050 ;
        RECT  0.955 0.245 1.015 1.050 ;
        RECT  0.805 0.355 0.955 0.840 ;
        RECT  0.665 0.355 0.805 0.475 ;
        RECT  0.665 0.720 0.805 0.840 ;
        RECT  0.595 0.245 0.665 0.475 ;
        RECT  0.595 0.720 0.665 1.050 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.375 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.675 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.910 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.990 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.950 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.475 ;
        RECT  0.665 0.720 0.735 0.840 ;
        RECT  0.595 0.245 0.665 0.475 ;
        RECT  0.595 0.720 0.665 1.050 ;
        RECT  0.525 0.545 0.705 0.615 ;
        RECT  0.455 0.345 0.525 0.915 ;
        RECT  0.130 0.345 0.455 0.415 ;
        RECT  0.310 0.845 0.455 0.915 ;
        RECT  0.230 0.845 0.310 1.075 ;
        RECT  0.050 0.205 0.130 0.415 ;
    END
END CKAN2D4BWP

MACRO CKAN2D8BWP
    CLASS CORE ;
    FOREIGN CKAN2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.720 1.890 0.950 ;
        RECT  1.790 0.210 1.870 0.455 ;
        RECT  1.490 0.335 1.790 0.455 ;
        RECT  1.410 0.215 1.490 0.455 ;
        RECT  1.295 0.335 1.410 0.455 ;
        RECT  1.110 0.335 1.295 0.950 ;
        RECT  1.085 0.215 1.110 0.950 ;
        RECT  1.030 0.215 1.085 0.455 ;
        RECT  0.630 0.720 1.085 0.950 ;
        RECT  0.730 0.335 1.030 0.455 ;
        RECT  0.650 0.215 0.730 0.455 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.350 ;
        RECT  1.700 -0.115 1.970 0.115 ;
        RECT  1.580 -0.115 1.700 0.255 ;
        RECT  1.320 -0.115 1.580 0.115 ;
        RECT  1.200 -0.115 1.320 0.255 ;
        RECT  0.940 -0.115 1.200 0.115 ;
        RECT  0.820 -0.115 0.940 0.255 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.675 2.050 1.375 ;
        RECT  0.540 1.145 1.970 1.375 ;
        RECT  0.420 0.990 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.720 1.890 0.950 ;
        RECT  1.790 0.210 1.870 0.455 ;
        RECT  1.490 0.335 1.790 0.455 ;
        RECT  1.410 0.215 1.490 0.455 ;
        RECT  1.365 0.335 1.410 0.455 ;
        RECT  0.730 0.335 1.015 0.455 ;
        RECT  0.630 0.720 1.015 0.950 ;
        RECT  0.650 0.215 0.730 0.455 ;
        RECT  1.395 0.545 1.920 0.615 ;
        RECT  0.540 0.545 0.985 0.615 ;
        RECT  0.470 0.205 0.540 0.915 ;
        RECT  0.125 0.205 0.470 0.275 ;
        RECT  0.305 0.845 0.470 0.915 ;
        RECT  0.235 0.845 0.305 1.050 ;
        RECT  0.055 0.205 0.125 0.355 ;
    END
END CKAN2D8BWP

MACRO CKBD0BWP
    CLASS CORE ;
    FOREIGN CKBD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0374 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.200 0.525 1.050 ;
        RECT  0.435 0.200 0.455 0.320 ;
        RECT  0.435 0.910 0.455 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0136 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.355 0.520 0.385 0.640 ;
        RECT  0.285 0.340 0.355 0.925 ;
        RECT  0.130 0.340 0.285 0.410 ;
        RECT  0.130 0.855 0.285 0.925 ;
        RECT  0.050 0.200 0.130 0.410 ;
        RECT  0.050 0.855 0.130 1.050 ;
    END
END CKBD0BWP

MACRO CKBD12BWP
    CLASS CORE ;
    FOREIGN CKBD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5987 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 0.195 2.890 0.450 ;
        RECT  2.135 0.725 2.885 0.955 ;
        RECT  2.510 0.290 2.810 0.450 ;
        RECT  2.430 0.190 2.510 0.450 ;
        RECT  2.150 0.290 2.430 0.450 ;
        RECT  2.135 0.190 2.150 0.450 ;
        RECT  2.070 0.190 2.135 0.955 ;
        RECT  1.790 0.290 2.070 0.955 ;
        RECT  1.785 0.190 1.790 0.955 ;
        RECT  1.710 0.190 1.785 0.450 ;
        RECT  0.970 0.725 1.785 0.955 ;
        RECT  1.430 0.290 1.710 0.450 ;
        RECT  1.350 0.190 1.430 0.450 ;
        RECT  1.070 0.290 1.350 0.450 ;
        RECT  0.990 0.190 1.070 0.450 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1088 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.455 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 2.940 0.115 ;
        RECT  0.800 -0.115 0.880 0.450 ;
        RECT  0.130 -0.115 0.800 0.115 ;
        RECT  0.050 -0.115 0.130 0.335 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 2.940 1.375 ;
        RECT  2.600 1.025 2.720 1.375 ;
        RECT  2.350 1.145 2.600 1.375 ;
        RECT  2.230 1.025 2.350 1.375 ;
        RECT  1.995 1.145 2.230 1.375 ;
        RECT  1.865 1.025 1.995 1.375 ;
        RECT  1.630 1.145 1.865 1.375 ;
        RECT  1.510 1.025 1.630 1.375 ;
        RECT  1.270 1.145 1.510 1.375 ;
        RECT  1.150 1.025 1.270 1.375 ;
        RECT  0.880 1.145 1.150 1.375 ;
        RECT  0.800 0.735 0.880 1.375 ;
        RECT  0.520 1.145 0.800 1.375 ;
        RECT  0.400 0.885 0.520 1.375 ;
        RECT  0.130 1.145 0.400 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.810 0.195 2.890 0.450 ;
        RECT  2.205 0.725 2.885 0.955 ;
        RECT  2.510 0.290 2.810 0.450 ;
        RECT  2.430 0.190 2.510 0.450 ;
        RECT  2.205 0.290 2.430 0.450 ;
        RECT  1.710 0.190 1.715 0.450 ;
        RECT  0.970 0.725 1.715 0.955 ;
        RECT  1.430 0.290 1.710 0.450 ;
        RECT  1.350 0.190 1.430 0.450 ;
        RECT  1.070 0.290 1.350 0.450 ;
        RECT  0.990 0.190 1.070 0.450 ;
        RECT  2.235 0.535 2.890 0.605 ;
        RECT  0.710 0.535 1.685 0.605 ;
        RECT  0.700 0.305 0.710 0.605 ;
        RECT  0.600 0.305 0.700 1.035 ;
        RECT  0.210 0.305 0.600 0.405 ;
        RECT  0.320 0.715 0.600 0.815 ;
        RECT  0.220 0.715 0.320 1.035 ;
    END
END CKBD12BWP

MACRO CKBD16BWP
    CLASS CORE ;
    FOREIGN CKBD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.195 3.730 0.455 ;
        RECT  2.695 0.725 3.725 0.955 ;
        RECT  3.370 0.295 3.650 0.455 ;
        RECT  3.290 0.195 3.370 0.455 ;
        RECT  3.010 0.295 3.290 0.455 ;
        RECT  2.930 0.195 3.010 0.455 ;
        RECT  2.695 0.295 2.930 0.455 ;
        RECT  2.650 0.295 2.695 0.955 ;
        RECT  2.555 0.195 2.650 0.955 ;
        RECT  2.345 0.295 2.555 0.955 ;
        RECT  2.290 0.295 2.345 0.455 ;
        RECT  1.110 0.725 2.345 0.955 ;
        RECT  2.210 0.195 2.290 0.455 ;
        RECT  1.930 0.295 2.210 0.455 ;
        RECT  1.850 0.195 1.930 0.455 ;
        RECT  1.570 0.295 1.850 0.455 ;
        RECT  1.490 0.195 1.570 0.455 ;
        RECT  1.210 0.295 1.490 0.455 ;
        RECT  1.130 0.195 1.210 0.455 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1360 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.625 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.115 3.780 0.115 ;
        RECT  0.950 -0.115 1.030 0.455 ;
        RECT  0.000 -0.115 0.950 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.145 3.780 1.375 ;
        RECT  3.450 1.025 3.570 1.375 ;
        RECT  3.210 1.145 3.450 1.375 ;
        RECT  3.090 1.025 3.210 1.375 ;
        RECT  2.850 1.145 3.090 1.375 ;
        RECT  2.730 1.025 2.850 1.375 ;
        RECT  2.490 1.145 2.730 1.375 ;
        RECT  2.370 1.025 2.490 1.375 ;
        RECT  2.130 1.145 2.370 1.375 ;
        RECT  2.010 1.025 2.130 1.375 ;
        RECT  1.770 1.145 2.010 1.375 ;
        RECT  1.650 1.025 1.770 1.375 ;
        RECT  1.410 1.145 1.650 1.375 ;
        RECT  1.290 1.025 1.410 1.375 ;
        RECT  1.030 1.145 1.290 1.375 ;
        RECT  0.950 0.695 1.030 1.375 ;
        RECT  0.690 1.145 0.950 1.375 ;
        RECT  0.570 0.890 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.195 3.730 0.455 ;
        RECT  2.765 0.725 3.725 0.955 ;
        RECT  3.370 0.295 3.650 0.455 ;
        RECT  3.290 0.195 3.370 0.455 ;
        RECT  3.010 0.295 3.290 0.455 ;
        RECT  2.930 0.195 3.010 0.455 ;
        RECT  2.765 0.295 2.930 0.455 ;
        RECT  2.210 0.195 2.275 0.455 ;
        RECT  1.110 0.725 2.275 0.955 ;
        RECT  1.930 0.295 2.210 0.455 ;
        RECT  1.850 0.195 1.930 0.455 ;
        RECT  1.570 0.295 1.850 0.455 ;
        RECT  1.490 0.195 1.570 0.455 ;
        RECT  1.210 0.295 1.490 0.455 ;
        RECT  1.130 0.195 1.210 0.455 ;
        RECT  2.810 0.535 3.540 0.605 ;
        RECT  0.870 0.535 2.210 0.605 ;
        RECT  0.860 0.305 0.870 0.605 ;
        RECT  0.760 0.305 0.860 1.030 ;
        RECT  0.130 0.305 0.760 0.395 ;
        RECT  0.500 0.720 0.760 0.820 ;
        RECT  0.400 0.720 0.500 1.030 ;
        RECT  0.140 0.720 0.400 0.820 ;
        RECT  0.050 0.720 0.140 1.030 ;
        RECT  0.050 0.225 0.130 0.395 ;
    END
END CKBD16BWP

MACRO CKBD1BWP
    CLASS CORE ;
    FOREIGN CKBD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0748 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.200 0.525 1.050 ;
        RECT  0.435 0.200 0.455 0.330 ;
        RECT  0.435 0.735 0.455 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.355 0.520 0.385 0.640 ;
        RECT  0.285 0.335 0.355 0.925 ;
        RECT  0.130 0.335 0.285 0.405 ;
        RECT  0.130 0.855 0.285 0.925 ;
        RECT  0.050 0.245 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.050 ;
    END
END CKBD1BWP

MACRO CKBD20BWP
    CLASS CORE ;
    FOREIGN CKBD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.710 4.330 0.940 ;
        RECT  4.220 0.190 4.300 0.450 ;
        RECT  3.910 0.310 4.220 0.450 ;
        RECT  3.830 0.190 3.910 0.450 ;
        RECT  3.550 0.310 3.830 0.450 ;
        RECT  3.470 0.190 3.550 0.450 ;
        RECT  3.190 0.310 3.470 0.450 ;
        RECT  3.115 0.190 3.190 0.450 ;
        RECT  3.110 0.190 3.115 0.940 ;
        RECT  2.830 0.310 3.110 0.940 ;
        RECT  2.765 0.190 2.830 0.940 ;
        RECT  2.750 0.190 2.765 0.450 ;
        RECT  1.290 0.710 2.765 0.940 ;
        RECT  2.470 0.310 2.750 0.450 ;
        RECT  2.390 0.190 2.470 0.450 ;
        RECT  2.110 0.310 2.390 0.450 ;
        RECT  2.030 0.190 2.110 0.450 ;
        RECT  1.750 0.310 2.030 0.450 ;
        RECT  1.670 0.190 1.750 0.450 ;
        RECT  1.390 0.310 1.670 0.450 ;
        RECT  1.310 0.190 1.390 0.450 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1632 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.785 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.490 -0.115 4.620 0.115 ;
        RECT  4.410 -0.115 4.490 0.450 ;
        RECT  4.120 -0.115 4.410 0.115 ;
        RECT  4.000 -0.115 4.120 0.240 ;
        RECT  3.750 -0.115 4.000 0.115 ;
        RECT  3.630 -0.115 3.750 0.240 ;
        RECT  3.390 -0.115 3.630 0.115 ;
        RECT  3.270 -0.115 3.390 0.240 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.240 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.240 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.240 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.240 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.240 ;
        RECT  1.210 -0.115 1.470 0.115 ;
        RECT  1.130 -0.115 1.210 0.450 ;
        RECT  0.130 -0.115 1.130 0.115 ;
        RECT  0.050 -0.115 0.130 0.350 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.485 1.145 4.620 1.375 ;
        RECT  4.415 0.750 4.485 1.375 ;
        RECT  4.120 1.145 4.415 1.375 ;
        RECT  4.000 1.010 4.120 1.375 ;
        RECT  3.750 1.145 4.000 1.375 ;
        RECT  3.630 1.010 3.750 1.375 ;
        RECT  3.390 1.145 3.630 1.375 ;
        RECT  3.270 1.010 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 1.010 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.010 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.010 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 1.010 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 1.010 1.590 1.375 ;
        RECT  1.210 1.145 1.470 1.375 ;
        RECT  1.130 0.695 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.910 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.910 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.705 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.710 4.330 0.940 ;
        RECT  4.220 0.190 4.300 0.450 ;
        RECT  3.910 0.310 4.220 0.450 ;
        RECT  3.830 0.190 3.910 0.450 ;
        RECT  3.550 0.310 3.830 0.450 ;
        RECT  3.470 0.190 3.550 0.450 ;
        RECT  3.190 0.310 3.470 0.450 ;
        RECT  3.185 0.190 3.190 0.450 ;
        RECT  2.470 0.310 2.695 0.450 ;
        RECT  1.290 0.710 2.695 0.940 ;
        RECT  2.390 0.190 2.470 0.450 ;
        RECT  2.110 0.310 2.390 0.450 ;
        RECT  2.030 0.190 2.110 0.450 ;
        RECT  1.750 0.310 2.030 0.450 ;
        RECT  1.670 0.190 1.750 0.450 ;
        RECT  1.390 0.310 1.670 0.450 ;
        RECT  1.310 0.190 1.390 0.450 ;
        RECT  3.245 0.525 4.295 0.595 ;
        RECT  1.050 0.525 2.635 0.595 ;
        RECT  0.940 0.290 1.050 1.035 ;
        RECT  0.210 0.290 0.940 0.390 ;
        RECT  0.680 0.740 0.940 0.840 ;
        RECT  0.580 0.740 0.680 1.035 ;
        RECT  0.320 0.740 0.580 0.840 ;
        RECT  0.220 0.740 0.320 1.035 ;
    END
END CKBD20BWP

MACRO CKBD24BWP
    CLASS CORE ;
    FOREIGN CKBD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.1424 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 0.190 5.190 0.450 ;
        RECT  3.815 0.710 5.185 0.940 ;
        RECT  4.830 0.310 5.110 0.450 ;
        RECT  4.750 0.190 4.830 0.450 ;
        RECT  4.470 0.310 4.750 0.450 ;
        RECT  4.390 0.190 4.470 0.450 ;
        RECT  4.110 0.310 4.390 0.450 ;
        RECT  4.030 0.190 4.110 0.450 ;
        RECT  3.815 0.310 4.030 0.450 ;
        RECT  3.750 0.310 3.815 0.940 ;
        RECT  3.670 0.190 3.750 0.940 ;
        RECT  3.465 0.310 3.670 0.940 ;
        RECT  3.390 0.310 3.465 0.450 ;
        RECT  1.490 0.710 3.465 0.940 ;
        RECT  3.310 0.190 3.390 0.450 ;
        RECT  3.030 0.310 3.310 0.450 ;
        RECT  2.950 0.190 3.030 0.450 ;
        RECT  2.670 0.310 2.950 0.450 ;
        RECT  2.590 0.190 2.670 0.450 ;
        RECT  2.310 0.310 2.590 0.450 ;
        RECT  2.230 0.190 2.310 0.450 ;
        RECT  1.950 0.310 2.230 0.450 ;
        RECT  1.870 0.190 1.950 0.450 ;
        RECT  1.590 0.310 1.870 0.450 ;
        RECT  1.510 0.190 1.590 0.450 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.945 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 -0.115 5.460 0.115 ;
        RECT  5.295 -0.115 5.365 0.310 ;
        RECT  5.030 -0.115 5.295 0.115 ;
        RECT  4.910 -0.115 5.030 0.240 ;
        RECT  4.670 -0.115 4.910 0.115 ;
        RECT  4.550 -0.115 4.670 0.240 ;
        RECT  4.310 -0.115 4.550 0.115 ;
        RECT  4.190 -0.115 4.310 0.240 ;
        RECT  3.950 -0.115 4.190 0.115 ;
        RECT  3.830 -0.115 3.950 0.240 ;
        RECT  3.590 -0.115 3.830 0.115 ;
        RECT  3.470 -0.115 3.590 0.240 ;
        RECT  3.230 -0.115 3.470 0.115 ;
        RECT  3.110 -0.115 3.230 0.240 ;
        RECT  2.870 -0.115 3.110 0.115 ;
        RECT  2.750 -0.115 2.870 0.240 ;
        RECT  2.510 -0.115 2.750 0.115 ;
        RECT  2.390 -0.115 2.510 0.240 ;
        RECT  2.150 -0.115 2.390 0.115 ;
        RECT  2.030 -0.115 2.150 0.240 ;
        RECT  1.790 -0.115 2.030 0.115 ;
        RECT  1.670 -0.115 1.790 0.240 ;
        RECT  1.410 -0.115 1.670 0.115 ;
        RECT  1.330 -0.115 1.410 0.450 ;
        RECT  0.000 -0.115 1.330 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 1.145 5.460 1.375 ;
        RECT  5.295 0.790 5.365 1.375 ;
        RECT  5.030 1.145 5.295 1.375 ;
        RECT  4.910 1.010 5.030 1.375 ;
        RECT  4.670 1.145 4.910 1.375 ;
        RECT  4.550 1.010 4.670 1.375 ;
        RECT  4.310 1.145 4.550 1.375 ;
        RECT  4.190 1.010 4.310 1.375 ;
        RECT  3.950 1.145 4.190 1.375 ;
        RECT  3.830 1.010 3.950 1.375 ;
        RECT  3.590 1.145 3.830 1.375 ;
        RECT  3.470 1.010 3.590 1.375 ;
        RECT  3.230 1.145 3.470 1.375 ;
        RECT  3.110 1.010 3.230 1.375 ;
        RECT  2.870 1.145 3.110 1.375 ;
        RECT  2.750 1.010 2.870 1.375 ;
        RECT  2.510 1.145 2.750 1.375 ;
        RECT  2.390 1.010 2.510 1.375 ;
        RECT  2.150 1.145 2.390 1.375 ;
        RECT  2.030 1.010 2.150 1.375 ;
        RECT  1.790 1.145 2.030 1.375 ;
        RECT  1.670 1.010 1.790 1.375 ;
        RECT  1.410 1.145 1.670 1.375 ;
        RECT  1.330 0.695 1.410 1.375 ;
        RECT  1.070 1.145 1.330 1.375 ;
        RECT  0.950 0.890 1.070 1.375 ;
        RECT  0.710 1.145 0.950 1.375 ;
        RECT  0.590 0.890 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 0.890 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.110 0.190 5.190 0.450 ;
        RECT  3.885 0.710 5.185 0.940 ;
        RECT  4.830 0.310 5.110 0.450 ;
        RECT  4.750 0.190 4.830 0.450 ;
        RECT  4.470 0.310 4.750 0.450 ;
        RECT  4.390 0.190 4.470 0.450 ;
        RECT  4.110 0.310 4.390 0.450 ;
        RECT  4.030 0.190 4.110 0.450 ;
        RECT  3.885 0.310 4.030 0.450 ;
        RECT  3.390 0.310 3.395 0.450 ;
        RECT  1.490 0.710 3.395 0.940 ;
        RECT  3.310 0.190 3.390 0.450 ;
        RECT  3.030 0.310 3.310 0.450 ;
        RECT  2.950 0.190 3.030 0.450 ;
        RECT  2.670 0.310 2.950 0.450 ;
        RECT  2.590 0.190 2.670 0.450 ;
        RECT  2.310 0.310 2.590 0.450 ;
        RECT  2.230 0.190 2.310 0.450 ;
        RECT  1.950 0.310 2.230 0.450 ;
        RECT  1.870 0.190 1.950 0.450 ;
        RECT  1.590 0.310 1.870 0.450 ;
        RECT  1.510 0.190 1.590 0.450 ;
        RECT  3.915 0.525 5.115 0.595 ;
        RECT  1.240 0.525 3.365 0.595 ;
        RECT  1.140 0.190 1.240 1.035 ;
        RECT  0.870 0.305 1.140 0.415 ;
        RECT  0.880 0.710 1.140 0.820 ;
        RECT  0.780 0.710 0.880 1.035 ;
        RECT  0.790 0.210 0.870 0.415 ;
        RECT  0.510 0.305 0.790 0.415 ;
        RECT  0.520 0.710 0.780 0.820 ;
        RECT  0.420 0.710 0.520 1.035 ;
        RECT  0.430 0.210 0.510 0.415 ;
        RECT  0.130 0.305 0.430 0.415 ;
        RECT  0.140 0.710 0.420 0.820 ;
        RECT  0.050 0.710 0.140 1.035 ;
        RECT  0.050 0.210 0.130 0.415 ;
    END
END CKBD24BWP

MACRO CKBD2BWP
    CLASS CORE ;
    FOREIGN CKBD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.405 0.665 0.840 ;
        RECT  0.575 0.405 0.595 0.475 ;
        RECT  0.575 0.755 0.595 0.840 ;
        RECT  0.505 0.245 0.575 0.475 ;
        RECT  0.505 0.755 0.575 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.115 0.840 0.115 ;
        RECT  0.690 -0.115 0.770 0.320 ;
        RECT  0.380 -0.115 0.690 0.115 ;
        RECT  0.260 -0.115 0.380 0.265 ;
        RECT  0.000 -0.115 0.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.145 0.840 1.375 ;
        RECT  0.690 0.920 0.770 1.375 ;
        RECT  0.380 1.145 0.690 1.375 ;
        RECT  0.260 0.995 0.380 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.420 0.545 0.510 0.615 ;
        RECT  0.350 0.335 0.420 0.925 ;
        RECT  0.150 0.335 0.350 0.405 ;
        RECT  0.150 0.855 0.350 0.925 ;
        RECT  0.070 0.245 0.150 0.405 ;
        RECT  0.070 0.855 0.150 1.050 ;
    END
END CKBD2BWP

MACRO CKBD3BWP
    CLASS CORE ;
    FOREIGN CKBD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.215 0.945 0.475 ;
        RECT  0.875 0.700 0.945 1.050 ;
        RECT  0.855 0.215 0.875 1.050 ;
        RECT  0.665 0.355 0.855 0.820 ;
        RECT  0.545 0.355 0.665 0.475 ;
        RECT  0.545 0.700 0.665 0.820 ;
        RECT  0.475 0.245 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.275 ;
        RECT  0.360 -0.115 0.640 0.115 ;
        RECT  0.240 -0.115 0.360 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 0.890 0.760 1.375 ;
        RECT  0.360 1.145 0.640 1.375 ;
        RECT  0.240 0.995 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.545 0.355 0.595 0.475 ;
        RECT  0.545 0.700 0.595 0.820 ;
        RECT  0.475 0.245 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.050 ;
        RECT  0.395 0.545 0.565 0.615 ;
        RECT  0.325 0.335 0.395 0.915 ;
        RECT  0.130 0.335 0.325 0.405 ;
        RECT  0.130 0.845 0.325 0.915 ;
        RECT  0.050 0.245 0.130 0.405 ;
        RECT  0.050 0.845 0.130 0.985 ;
    END
END CKBD3BWP

MACRO CKBD4BWP
    CLASS CORE ;
    FOREIGN CKBD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1904 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.235 1.025 0.495 ;
        RECT  1.015 0.700 1.025 1.050 ;
        RECT  0.955 0.235 1.015 1.050 ;
        RECT  0.805 0.355 0.955 0.820 ;
        RECT  0.665 0.355 0.805 0.475 ;
        RECT  0.665 0.700 0.805 0.820 ;
        RECT  0.595 0.235 0.665 0.475 ;
        RECT  0.595 0.700 0.665 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.440 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.280 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.365 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.675 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.890 0.870 1.375 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.910 0.490 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.475 ;
        RECT  0.665 0.700 0.735 0.820 ;
        RECT  0.595 0.235 0.665 0.475 ;
        RECT  0.595 0.700 0.665 1.050 ;
        RECT  0.380 0.545 0.650 0.615 ;
        RECT  0.310 0.350 0.380 0.820 ;
        RECT  0.305 0.350 0.310 0.420 ;
        RECT  0.305 0.750 0.310 0.820 ;
        RECT  0.235 0.245 0.305 0.420 ;
        RECT  0.235 0.750 0.305 1.045 ;
    END
END CKBD4BWP

MACRO CKBD6BWP
    CLASS CORE ;
    FOREIGN CKBD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2856 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.235 1.445 0.475 ;
        RECT  1.375 0.700 1.445 1.015 ;
        RECT  1.155 0.355 1.375 0.475 ;
        RECT  1.155 0.700 1.375 0.820 ;
        RECT  1.085 0.355 1.155 0.820 ;
        RECT  1.065 0.355 1.085 1.045 ;
        RECT  0.995 0.235 1.065 1.045 ;
        RECT  0.945 0.355 0.995 0.820 ;
        RECT  0.685 0.355 0.945 0.475 ;
        RECT  0.685 0.700 0.945 0.820 ;
        RECT  0.615 0.235 0.685 0.475 ;
        RECT  0.615 0.700 0.685 1.015 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.375 ;
        RECT  1.280 -0.115 1.550 0.115 ;
        RECT  1.160 -0.115 1.280 0.275 ;
        RECT  0.900 -0.115 1.160 0.115 ;
        RECT  0.780 -0.115 0.900 0.275 ;
        RECT  0.500 -0.115 0.780 0.115 ;
        RECT  0.420 -0.115 0.500 0.280 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.365 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.685 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 0.890 1.280 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.780 0.890 0.900 1.375 ;
        RECT  0.500 1.145 0.780 1.375 ;
        RECT  0.420 0.895 0.500 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.235 1.445 0.475 ;
        RECT  1.375 0.700 1.445 1.015 ;
        RECT  1.225 0.355 1.375 0.475 ;
        RECT  1.225 0.700 1.375 0.820 ;
        RECT  0.685 0.355 0.875 0.475 ;
        RECT  0.685 0.700 0.875 0.820 ;
        RECT  0.615 0.235 0.685 0.475 ;
        RECT  0.615 0.700 0.685 1.015 ;
        RECT  1.255 0.545 1.605 0.615 ;
        RECT  0.380 0.545 0.845 0.615 ;
        RECT  0.310 0.350 0.380 0.805 ;
        RECT  0.305 0.350 0.310 0.420 ;
        RECT  0.305 0.735 0.310 0.805 ;
        RECT  0.235 0.260 0.305 0.420 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END CKBD6BWP

MACRO CKBD8BWP
    CLASS CORE ;
    FOREIGN CKBD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3808 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.720 2.030 0.950 ;
        RECT  1.930 0.255 2.010 0.455 ;
        RECT  1.630 0.350 1.930 0.455 ;
        RECT  1.575 0.255 1.630 0.455 ;
        RECT  1.550 0.255 1.575 0.950 ;
        RECT  1.250 0.345 1.550 0.950 ;
        RECT  1.225 0.215 1.250 0.950 ;
        RECT  1.170 0.215 1.225 0.455 ;
        RECT  0.770 0.720 1.225 0.950 ;
        RECT  0.870 0.345 1.170 0.455 ;
        RECT  0.790 0.255 0.870 0.455 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0816 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.290 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.395 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.720 -0.115 1.840 0.275 ;
        RECT  1.460 -0.115 1.720 0.115 ;
        RECT  1.340 -0.115 1.460 0.275 ;
        RECT  1.080 -0.115 1.340 0.115 ;
        RECT  0.960 -0.115 1.080 0.275 ;
        RECT  0.690 -0.115 0.960 0.115 ;
        RECT  0.610 -0.115 0.690 0.460 ;
        RECT  0.340 -0.115 0.610 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.675 2.190 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.720 1.020 1.840 1.375 ;
        RECT  1.460 1.145 1.720 1.375 ;
        RECT  1.340 1.020 1.460 1.375 ;
        RECT  1.080 1.145 1.340 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.690 1.145 0.960 1.375 ;
        RECT  0.610 0.735 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.920 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.720 2.030 0.950 ;
        RECT  1.930 0.255 2.010 0.455 ;
        RECT  1.645 0.350 1.930 0.455 ;
        RECT  0.870 0.345 1.155 0.455 ;
        RECT  0.770 0.720 1.155 0.950 ;
        RECT  0.790 0.255 0.870 0.455 ;
        RECT  1.675 0.545 2.060 0.615 ;
        RECT  0.520 0.545 1.125 0.615 ;
        RECT  0.420 0.255 0.520 1.035 ;
        RECT  0.125 0.345 0.420 0.425 ;
        RECT  0.125 0.740 0.420 0.840 ;
        RECT  0.055 0.265 0.125 0.425 ;
        RECT  0.055 0.740 0.125 1.035 ;
    END
END CKBD8BWP

MACRO CKLHQD12BWP
    CLASS CORE ;
    FOREIGN CKLHQD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.6048 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.435 0.185 5.505 0.465 ;
        RECT  5.435 0.700 5.505 1.035 ;
        RECT  5.125 0.345 5.435 0.465 ;
        RECT  5.145 0.700 5.435 0.820 ;
        RECT  5.075 0.700 5.145 1.035 ;
        RECT  5.055 0.185 5.125 0.465 ;
        RECT  4.785 0.700 5.075 0.820 ;
        RECT  4.745 0.345 5.055 0.465 ;
        RECT  4.715 0.700 4.785 1.035 ;
        RECT  4.675 0.185 4.745 0.465 ;
        RECT  4.655 0.700 4.715 0.820 ;
        RECT  4.655 0.345 4.675 0.465 ;
        RECT  4.425 0.345 4.655 0.820 ;
        RECT  4.365 0.345 4.425 1.035 ;
        RECT  4.355 0.185 4.365 1.035 ;
        RECT  4.305 0.185 4.355 0.820 ;
        RECT  4.295 0.185 4.305 0.465 ;
        RECT  4.065 0.700 4.305 0.820 ;
        RECT  3.985 0.345 4.295 0.465 ;
        RECT  3.995 0.700 4.065 1.035 ;
        RECT  3.705 0.700 3.995 0.820 ;
        RECT  3.915 0.185 3.985 0.465 ;
        RECT  3.625 0.345 3.915 0.465 ;
        RECT  3.635 0.700 3.705 1.035 ;
        RECT  3.555 0.185 3.625 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0822 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.205 0.520 3.275 0.795 ;
        RECT  2.630 0.725 3.205 0.795 ;
        RECT  2.510 0.545 2.630 0.795 ;
        RECT  2.485 0.725 2.510 0.795 ;
        RECT  2.415 0.725 2.485 0.925 ;
        RECT  1.785 0.855 2.415 0.925 ;
        RECT  1.700 0.635 1.785 0.925 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 -0.115 5.740 0.115 ;
        RECT  5.615 -0.115 5.685 0.465 ;
        RECT  5.340 -0.115 5.615 0.115 ;
        RECT  5.220 -0.115 5.340 0.275 ;
        RECT  4.960 -0.115 5.220 0.115 ;
        RECT  4.840 -0.115 4.960 0.275 ;
        RECT  4.580 -0.115 4.840 0.115 ;
        RECT  4.460 -0.115 4.580 0.275 ;
        RECT  4.200 -0.115 4.460 0.115 ;
        RECT  4.080 -0.115 4.200 0.275 ;
        RECT  3.830 -0.115 4.080 0.115 ;
        RECT  3.710 -0.115 3.830 0.270 ;
        RECT  3.420 -0.115 3.710 0.115 ;
        RECT  3.340 -0.115 3.420 0.275 ;
        RECT  2.265 -0.115 3.340 0.115 ;
        RECT  2.195 -0.115 2.265 0.305 ;
        RECT  1.045 -0.115 2.195 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.145 5.740 1.375 ;
        RECT  5.615 0.680 5.685 1.375 ;
        RECT  5.350 1.145 5.615 1.375 ;
        RECT  5.230 0.890 5.350 1.375 ;
        RECT  4.990 1.145 5.230 1.375 ;
        RECT  4.870 0.890 4.990 1.375 ;
        RECT  4.630 1.145 4.870 1.375 ;
        RECT  4.510 0.890 4.630 1.375 ;
        RECT  4.270 1.145 4.510 1.375 ;
        RECT  4.150 0.890 4.270 1.375 ;
        RECT  3.910 1.145 4.150 1.375 ;
        RECT  3.790 0.890 3.910 1.375 ;
        RECT  3.550 1.145 3.790 1.375 ;
        RECT  3.430 1.005 3.550 1.375 ;
        RECT  3.010 1.145 3.430 1.375 ;
        RECT  2.890 1.005 3.010 1.375 ;
        RECT  1.080 1.145 2.890 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.435 0.185 5.505 0.465 ;
        RECT  5.435 0.700 5.505 1.035 ;
        RECT  5.125 0.345 5.435 0.465 ;
        RECT  5.145 0.700 5.435 0.820 ;
        RECT  5.075 0.700 5.145 1.035 ;
        RECT  5.055 0.185 5.125 0.465 ;
        RECT  4.785 0.700 5.075 0.820 ;
        RECT  4.745 0.345 5.055 0.465 ;
        RECT  4.725 0.700 4.785 1.035 ;
        RECT  4.725 0.185 4.745 0.465 ;
        RECT  3.985 0.345 4.235 0.465 ;
        RECT  4.065 0.700 4.235 0.820 ;
        RECT  3.995 0.700 4.065 1.035 ;
        RECT  3.705 0.700 3.995 0.820 ;
        RECT  3.915 0.185 3.985 0.465 ;
        RECT  3.625 0.345 3.915 0.465 ;
        RECT  3.635 0.700 3.705 1.035 ;
        RECT  3.555 0.185 3.625 0.465 ;
        RECT  4.755 0.545 5.435 0.615 ;
        RECT  3.445 0.545 4.205 0.615 ;
        RECT  3.375 0.355 3.445 0.935 ;
        RECT  3.240 0.355 3.375 0.425 ;
        RECT  2.625 0.865 3.375 0.935 ;
        RECT  3.170 0.215 3.240 0.425 ;
        RECT  2.350 0.215 3.170 0.285 ;
        RECT  2.900 0.375 2.980 0.640 ;
        RECT  2.335 0.375 2.900 0.445 ;
        RECT  2.555 0.865 2.625 1.035 ;
        RECT  2.265 0.375 2.335 0.785 ;
        RECT  2.085 0.375 2.265 0.445 ;
        RECT  1.970 0.715 2.265 0.785 ;
        RECT  1.935 0.540 2.180 0.610 ;
        RECT  2.015 0.185 2.085 0.445 ;
        RECT  1.865 0.210 1.935 0.610 ;
        RECT  1.590 0.995 1.870 1.065 ;
        RECT  1.260 0.210 1.865 0.280 ;
        RECT  1.715 0.360 1.785 0.480 ;
        RECT  1.590 0.410 1.715 0.480 ;
        RECT  1.520 0.410 1.590 1.065 ;
        RECT  1.470 0.520 1.520 0.640 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.360 1.400 1.050 ;
        RECT  1.330 0.360 1.355 0.950 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.190 0.210 1.260 0.800 ;
        RECT  1.130 0.210 1.190 0.280 ;
        RECT  1.175 0.680 1.190 0.800 ;
        RECT  0.955 0.680 1.175 0.750 ;
        RECT  1.050 0.370 1.120 0.550 ;
        RECT  0.770 0.370 1.050 0.440 ;
        RECT  0.885 0.610 0.955 0.750 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.185 0.770 0.800 ;
        RECT  0.590 0.185 0.700 0.255 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.335 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD12BWP

MACRO CKLHQD16BWP
    CLASS CORE ;
    FOREIGN CKLHQD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.8064 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.415 0.185 6.485 0.465 ;
        RECT  6.415 0.700 6.485 1.035 ;
        RECT  6.125 0.345 6.415 0.465 ;
        RECT  6.125 0.700 6.415 0.820 ;
        RECT  6.055 0.185 6.125 0.465 ;
        RECT  6.055 0.700 6.125 1.035 ;
        RECT  5.765 0.345 6.055 0.465 ;
        RECT  5.765 0.700 6.055 0.820 ;
        RECT  5.695 0.185 5.765 0.465 ;
        RECT  5.695 0.700 5.765 1.035 ;
        RECT  5.405 0.345 5.695 0.465 ;
        RECT  5.405 0.700 5.695 0.820 ;
        RECT  5.355 0.185 5.405 0.465 ;
        RECT  5.355 0.700 5.405 1.035 ;
        RECT  5.335 0.185 5.355 1.035 ;
        RECT  5.045 0.345 5.335 0.820 ;
        RECT  5.005 0.185 5.045 1.035 ;
        RECT  4.975 0.185 5.005 0.465 ;
        RECT  4.975 0.700 5.005 1.035 ;
        RECT  4.685 0.345 4.975 0.465 ;
        RECT  4.685 0.700 4.975 0.820 ;
        RECT  4.615 0.185 4.685 0.465 ;
        RECT  4.615 0.700 4.685 1.035 ;
        RECT  4.325 0.345 4.615 0.465 ;
        RECT  4.325 0.700 4.615 0.820 ;
        RECT  4.255 0.185 4.325 0.465 ;
        RECT  4.255 0.700 4.325 1.035 ;
        RECT  3.965 0.345 4.255 0.465 ;
        RECT  3.965 0.700 4.255 0.820 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.700 3.965 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.545 3.360 0.795 ;
        RECT  2.690 0.725 3.240 0.795 ;
        RECT  2.570 0.545 2.690 0.795 ;
        RECT  2.535 0.725 2.570 0.795 ;
        RECT  2.465 0.725 2.535 0.960 ;
        RECT  1.945 0.890 2.465 0.960 ;
        RECT  1.875 0.695 1.945 0.960 ;
        RECT  1.790 0.695 1.875 0.765 ;
        RECT  1.700 0.495 1.790 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 -0.115 6.720 0.115 ;
        RECT  6.595 -0.115 6.665 0.465 ;
        RECT  6.330 -0.115 6.595 0.115 ;
        RECT  6.210 -0.115 6.330 0.275 ;
        RECT  5.970 -0.115 6.210 0.115 ;
        RECT  5.850 -0.115 5.970 0.275 ;
        RECT  5.610 -0.115 5.850 0.115 ;
        RECT  5.490 -0.115 5.610 0.275 ;
        RECT  5.250 -0.115 5.490 0.115 ;
        RECT  5.130 -0.115 5.250 0.275 ;
        RECT  4.890 -0.115 5.130 0.115 ;
        RECT  4.770 -0.115 4.890 0.275 ;
        RECT  4.530 -0.115 4.770 0.115 ;
        RECT  4.410 -0.115 4.530 0.275 ;
        RECT  4.170 -0.115 4.410 0.115 ;
        RECT  4.050 -0.115 4.170 0.275 ;
        RECT  3.785 -0.115 4.050 0.115 ;
        RECT  3.715 -0.115 3.785 0.300 ;
        RECT  2.285 -0.115 3.715 0.115 ;
        RECT  2.215 -0.115 2.285 0.305 ;
        RECT  1.025 -0.115 2.215 0.115 ;
        RECT  0.955 -0.115 1.025 0.290 ;
        RECT  0.300 -0.115 0.955 0.115 ;
        RECT  0.230 -0.115 0.300 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.145 6.720 1.375 ;
        RECT  6.595 0.675 6.665 1.375 ;
        RECT  6.330 1.145 6.595 1.375 ;
        RECT  6.210 0.890 6.330 1.375 ;
        RECT  5.970 1.145 6.210 1.375 ;
        RECT  5.850 0.890 5.970 1.375 ;
        RECT  5.610 1.145 5.850 1.375 ;
        RECT  5.490 0.890 5.610 1.375 ;
        RECT  5.250 1.145 5.490 1.375 ;
        RECT  5.130 0.890 5.250 1.375 ;
        RECT  4.890 1.145 5.130 1.375 ;
        RECT  4.770 0.890 4.890 1.375 ;
        RECT  4.530 1.145 4.770 1.375 ;
        RECT  4.410 0.890 4.530 1.375 ;
        RECT  4.170 1.145 4.410 1.375 ;
        RECT  4.050 0.890 4.170 1.375 ;
        RECT  3.800 1.145 4.050 1.375 ;
        RECT  3.680 1.005 3.800 1.375 ;
        RECT  3.070 1.145 3.680 1.375 ;
        RECT  2.950 1.005 3.070 1.375 ;
        RECT  2.350 1.145 2.950 1.375 ;
        RECT  2.230 1.030 2.350 1.375 ;
        RECT  1.630 1.145 2.230 1.375 ;
        RECT  1.510 1.010 1.630 1.375 ;
        RECT  1.080 1.145 1.510 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.415 0.185 6.485 0.465 ;
        RECT  6.415 0.700 6.485 1.035 ;
        RECT  6.125 0.345 6.415 0.465 ;
        RECT  6.125 0.700 6.415 0.820 ;
        RECT  6.055 0.185 6.125 0.465 ;
        RECT  6.055 0.700 6.125 1.035 ;
        RECT  5.765 0.345 6.055 0.465 ;
        RECT  5.765 0.700 6.055 0.820 ;
        RECT  5.695 0.185 5.765 0.465 ;
        RECT  5.695 0.700 5.765 1.035 ;
        RECT  5.425 0.345 5.695 0.465 ;
        RECT  5.425 0.700 5.695 0.820 ;
        RECT  4.685 0.345 4.935 0.465 ;
        RECT  4.685 0.700 4.935 0.820 ;
        RECT  4.615 0.185 4.685 0.465 ;
        RECT  4.615 0.700 4.685 1.035 ;
        RECT  4.325 0.345 4.615 0.465 ;
        RECT  4.325 0.700 4.615 0.820 ;
        RECT  4.255 0.185 4.325 0.465 ;
        RECT  4.255 0.700 4.325 1.035 ;
        RECT  3.965 0.345 4.255 0.465 ;
        RECT  3.965 0.700 4.255 0.820 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.700 3.965 1.035 ;
        RECT  5.455 0.545 6.445 0.615 ;
        RECT  3.815 0.545 4.905 0.615 ;
        RECT  3.745 0.380 3.815 0.935 ;
        RECT  3.640 0.380 3.745 0.450 ;
        RECT  3.430 0.865 3.745 0.935 ;
        RECT  3.605 0.520 3.675 0.640 ;
        RECT  3.570 0.215 3.640 0.450 ;
        RECT  3.500 0.520 3.605 0.590 ;
        RECT  2.370 0.215 3.570 0.285 ;
        RECT  3.430 0.395 3.500 0.590 ;
        RECT  3.035 0.395 3.430 0.465 ;
        RECT  3.310 0.865 3.430 1.075 ;
        RECT  2.685 0.865 3.310 0.935 ;
        RECT  2.965 0.395 3.035 0.640 ;
        RECT  2.395 0.395 2.965 0.465 ;
        RECT  2.615 0.865 2.685 1.035 ;
        RECT  2.325 0.395 2.395 0.820 ;
        RECT  2.105 0.395 2.325 0.465 ;
        RECT  2.040 0.750 2.325 0.820 ;
        RECT  1.940 0.545 2.130 0.615 ;
        RECT  2.035 0.185 2.105 0.465 ;
        RECT  1.870 0.210 1.940 0.615 ;
        RECT  1.230 0.210 1.870 0.280 ;
        RECT  1.715 0.835 1.785 1.050 ;
        RECT  1.590 0.355 1.770 0.425 ;
        RECT  1.590 0.835 1.715 0.905 ;
        RECT  1.520 0.355 1.590 0.905 ;
        RECT  1.470 0.690 1.520 0.810 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.360 1.400 1.050 ;
        RECT  1.330 0.360 1.355 0.950 ;
        RECT  1.300 0.360 1.330 0.460 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.230 0.680 1.240 0.800 ;
        RECT  1.160 0.210 1.230 0.800 ;
        RECT  1.110 0.210 1.160 0.280 ;
        RECT  0.955 0.730 1.160 0.800 ;
        RECT  1.020 0.370 1.090 0.550 ;
        RECT  0.770 0.370 1.020 0.440 ;
        RECT  0.885 0.620 0.955 0.800 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.185 0.770 0.800 ;
        RECT  0.580 0.185 0.700 0.285 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.525 0.355 0.590 0.640 ;
        RECT  0.520 0.355 0.525 1.055 ;
        RECT  0.455 0.570 0.520 1.055 ;
        RECT  0.440 0.195 0.510 0.265 ;
        RECT  0.370 0.195 0.440 0.415 ;
        RECT  0.125 0.345 0.370 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD16BWP

MACRO CKLHQD1BWP
    CLASS CORE ;
    FOREIGN CKLHQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.185 2.905 1.045 ;
        RECT  2.815 0.185 2.835 0.465 ;
        RECT  2.815 0.745 2.835 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 1.795 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.940 0.115 ;
        RECT  2.640 -0.115 2.710 0.440 ;
        RECT  1.045 -0.115 2.640 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.145 2.940 1.375 ;
        RECT  2.610 1.005 2.730 1.375 ;
        RECT  1.650 1.145 2.610 1.375 ;
        RECT  1.530 1.000 1.650 1.375 ;
        RECT  1.100 1.145 1.530 1.375 ;
        RECT  0.980 1.020 1.100 1.375 ;
        RECT  0.130 1.145 0.980 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.745 0.520 2.765 0.640 ;
        RECT  2.675 0.520 2.745 0.920 ;
        RECT  1.985 0.850 2.675 0.920 ;
        RECT  2.500 0.330 2.570 0.780 ;
        RECT  2.455 0.330 2.500 0.450 ;
        RECT  2.235 0.710 2.500 0.780 ;
        RECT  2.385 0.530 2.430 0.630 ;
        RECT  2.315 0.195 2.385 0.630 ;
        RECT  1.270 0.195 2.315 0.265 ;
        RECT  2.165 0.520 2.235 0.780 ;
        RECT  1.985 0.355 2.170 0.425 ;
        RECT  1.915 0.355 1.985 1.035 ;
        RECT  1.585 0.355 1.810 0.425 ;
        RECT  1.735 0.860 1.805 1.035 ;
        RECT  1.585 0.860 1.735 0.930 ;
        RECT  1.515 0.355 1.585 0.930 ;
        RECT  1.480 0.665 1.515 0.785 ;
        RECT  1.410 0.885 1.445 1.025 ;
        RECT  1.340 0.345 1.410 1.025 ;
        RECT  0.835 0.880 1.340 0.950 ;
        RECT  1.200 0.195 1.270 0.810 ;
        RECT  1.130 0.195 1.200 0.265 ;
        RECT  0.935 0.740 1.200 0.810 ;
        RECT  1.060 0.370 1.130 0.640 ;
        RECT  0.770 0.370 1.060 0.440 ;
        RECT  0.865 0.520 0.935 0.810 ;
        RECT  0.765 0.880 0.835 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.525 0.985 0.765 1.055 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.345 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD1BWP

MACRO CKLHQD20BWP
    CLASS CORE ;
    FOREIGN CKLHQD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.0080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.255 0.185 7.325 0.465 ;
        RECT  7.255 0.700 7.325 1.035 ;
        RECT  6.965 0.345 7.255 0.465 ;
        RECT  6.965 0.700 7.255 0.820 ;
        RECT  6.895 0.185 6.965 0.465 ;
        RECT  6.895 0.700 6.965 1.035 ;
        RECT  6.605 0.345 6.895 0.465 ;
        RECT  6.605 0.700 6.895 0.820 ;
        RECT  6.535 0.185 6.605 0.465 ;
        RECT  6.535 0.700 6.605 1.035 ;
        RECT  6.245 0.345 6.535 0.465 ;
        RECT  6.245 0.700 6.535 0.820 ;
        RECT  6.175 0.185 6.245 0.465 ;
        RECT  6.175 0.700 6.245 1.035 ;
        RECT  5.885 0.345 6.175 0.465 ;
        RECT  5.885 0.700 6.175 0.820 ;
        RECT  5.815 0.185 5.885 0.465 ;
        RECT  5.815 0.700 5.885 1.035 ;
        RECT  5.775 0.345 5.815 0.465 ;
        RECT  5.775 0.700 5.815 0.820 ;
        RECT  5.525 0.345 5.775 0.820 ;
        RECT  5.455 0.185 5.525 1.035 ;
        RECT  5.425 0.345 5.455 0.820 ;
        RECT  5.165 0.345 5.425 0.465 ;
        RECT  5.165 0.700 5.425 0.820 ;
        RECT  5.095 0.185 5.165 0.465 ;
        RECT  5.095 0.700 5.165 1.035 ;
        RECT  4.805 0.345 5.095 0.465 ;
        RECT  4.805 0.700 5.095 0.820 ;
        RECT  4.735 0.185 4.805 0.465 ;
        RECT  4.735 0.700 4.805 1.035 ;
        RECT  4.445 0.345 4.735 0.465 ;
        RECT  4.445 0.700 4.735 0.820 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.700 4.445 1.035 ;
        RECT  4.065 0.345 4.375 0.465 ;
        RECT  4.085 0.700 4.375 0.820 ;
        RECT  4.015 0.700 4.085 1.035 ;
        RECT  3.995 0.185 4.065 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1048 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.545 3.490 0.795 ;
        RECT  2.790 0.725 3.370 0.795 ;
        RECT  2.670 0.545 2.790 0.795 ;
        RECT  2.605 0.725 2.670 0.795 ;
        RECT  2.535 0.725 2.605 0.960 ;
        RECT  2.020 0.890 2.535 0.960 ;
        RECT  1.950 0.835 2.020 0.960 ;
        RECT  1.795 0.835 1.950 0.905 ;
        RECT  1.695 0.495 1.795 0.905 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.505 -0.115 7.560 0.115 ;
        RECT  7.435 -0.115 7.505 0.465 ;
        RECT  7.170 -0.115 7.435 0.115 ;
        RECT  7.050 -0.115 7.170 0.275 ;
        RECT  6.810 -0.115 7.050 0.115 ;
        RECT  6.690 -0.115 6.810 0.275 ;
        RECT  6.450 -0.115 6.690 0.115 ;
        RECT  6.330 -0.115 6.450 0.275 ;
        RECT  6.090 -0.115 6.330 0.115 ;
        RECT  5.970 -0.115 6.090 0.275 ;
        RECT  5.730 -0.115 5.970 0.115 ;
        RECT  5.610 -0.115 5.730 0.275 ;
        RECT  5.370 -0.115 5.610 0.115 ;
        RECT  5.250 -0.115 5.370 0.275 ;
        RECT  5.010 -0.115 5.250 0.115 ;
        RECT  4.890 -0.115 5.010 0.275 ;
        RECT  4.650 -0.115 4.890 0.115 ;
        RECT  4.530 -0.115 4.650 0.275 ;
        RECT  4.280 -0.115 4.530 0.115 ;
        RECT  4.160 -0.115 4.280 0.275 ;
        RECT  2.365 -0.115 4.160 0.115 ;
        RECT  2.295 -0.115 2.365 0.305 ;
        RECT  1.045 -0.115 2.295 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.505 1.145 7.560 1.375 ;
        RECT  7.435 0.675 7.505 1.375 ;
        RECT  7.170 1.145 7.435 1.375 ;
        RECT  7.050 0.890 7.170 1.375 ;
        RECT  6.810 1.145 7.050 1.375 ;
        RECT  6.690 0.890 6.810 1.375 ;
        RECT  6.450 1.145 6.690 1.375 ;
        RECT  6.330 0.890 6.450 1.375 ;
        RECT  6.090 1.145 6.330 1.375 ;
        RECT  5.970 0.890 6.090 1.375 ;
        RECT  5.730 1.145 5.970 1.375 ;
        RECT  5.610 0.890 5.730 1.375 ;
        RECT  5.370 1.145 5.610 1.375 ;
        RECT  5.250 0.890 5.370 1.375 ;
        RECT  5.010 1.145 5.250 1.375 ;
        RECT  4.890 0.890 5.010 1.375 ;
        RECT  4.650 1.145 4.890 1.375 ;
        RECT  4.530 0.890 4.650 1.375 ;
        RECT  4.290 1.145 4.530 1.375 ;
        RECT  4.170 0.890 4.290 1.375 ;
        RECT  3.900 1.145 4.170 1.375 ;
        RECT  3.780 1.005 3.900 1.375 ;
        RECT  3.140 1.145 3.780 1.375 ;
        RECT  3.020 1.005 3.140 1.375 ;
        RECT  2.410 1.145 3.020 1.375 ;
        RECT  2.290 1.030 2.410 1.375 ;
        RECT  2.040 1.145 2.290 1.375 ;
        RECT  1.920 1.110 2.040 1.375 ;
        RECT  1.080 1.145 1.920 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.255 0.185 7.325 0.465 ;
        RECT  7.255 0.700 7.325 1.035 ;
        RECT  6.965 0.345 7.255 0.465 ;
        RECT  6.965 0.700 7.255 0.820 ;
        RECT  6.895 0.185 6.965 0.465 ;
        RECT  6.895 0.700 6.965 1.035 ;
        RECT  6.605 0.345 6.895 0.465 ;
        RECT  6.605 0.700 6.895 0.820 ;
        RECT  6.535 0.185 6.605 0.465 ;
        RECT  6.535 0.700 6.605 1.035 ;
        RECT  6.245 0.345 6.535 0.465 ;
        RECT  6.245 0.700 6.535 0.820 ;
        RECT  6.175 0.185 6.245 0.465 ;
        RECT  6.175 0.700 6.245 1.035 ;
        RECT  5.885 0.345 6.175 0.465 ;
        RECT  5.885 0.700 6.175 0.820 ;
        RECT  5.845 0.185 5.885 0.465 ;
        RECT  5.845 0.700 5.885 1.035 ;
        RECT  5.165 0.345 5.355 0.465 ;
        RECT  5.165 0.700 5.355 0.820 ;
        RECT  5.095 0.185 5.165 0.465 ;
        RECT  5.095 0.700 5.165 1.035 ;
        RECT  4.805 0.345 5.095 0.465 ;
        RECT  4.805 0.700 5.095 0.820 ;
        RECT  4.735 0.185 4.805 0.465 ;
        RECT  4.735 0.700 4.805 1.035 ;
        RECT  4.445 0.345 4.735 0.465 ;
        RECT  4.445 0.700 4.735 0.820 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.700 4.445 1.035 ;
        RECT  4.065 0.345 4.375 0.465 ;
        RECT  4.085 0.700 4.375 0.820 ;
        RECT  4.015 0.700 4.085 1.035 ;
        RECT  3.995 0.185 4.065 0.465 ;
        RECT  5.875 0.545 7.375 0.615 ;
        RECT  3.915 0.545 5.325 0.615 ;
        RECT  3.845 0.215 3.915 0.935 ;
        RECT  2.450 0.215 3.845 0.285 ;
        RECT  3.510 0.865 3.845 0.935 ;
        RECT  3.685 0.395 3.755 0.640 ;
        RECT  3.105 0.395 3.685 0.465 ;
        RECT  3.390 0.865 3.510 1.075 ;
        RECT  2.745 0.865 3.390 0.935 ;
        RECT  3.035 0.395 3.105 0.640 ;
        RECT  2.455 0.395 3.035 0.465 ;
        RECT  2.675 0.865 2.745 1.035 ;
        RECT  2.385 0.395 2.455 0.820 ;
        RECT  2.185 0.395 2.385 0.465 ;
        RECT  2.100 0.750 2.385 0.820 ;
        RECT  2.020 0.545 2.250 0.615 ;
        RECT  2.115 0.185 2.185 0.465 ;
        RECT  1.950 0.210 2.020 0.615 ;
        RECT  1.260 0.210 1.950 0.280 ;
        RECT  1.615 0.975 1.870 1.045 ;
        RECT  1.615 0.355 1.830 0.425 ;
        RECT  1.545 0.355 1.615 1.045 ;
        RECT  1.470 0.520 1.545 0.640 ;
        RECT  1.400 0.355 1.450 0.425 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.355 1.400 1.050 ;
        RECT  1.330 0.355 1.355 0.950 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.190 0.210 1.260 0.800 ;
        RECT  1.130 0.210 1.190 0.280 ;
        RECT  1.170 0.660 1.190 0.800 ;
        RECT  0.955 0.730 1.170 0.800 ;
        RECT  1.050 0.370 1.120 0.550 ;
        RECT  0.770 0.370 1.050 0.440 ;
        RECT  0.885 0.610 0.955 0.800 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.185 0.770 0.800 ;
        RECT  0.590 0.185 0.700 0.255 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.335 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.185 0.510 0.255 ;
        RECT  0.380 0.185 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD20BWP

MACRO CKLHQD24BWP
    CLASS CORE ;
    FOREIGN CKLHQD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.2096 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.375 0.185 8.445 0.465 ;
        RECT  8.375 0.700 8.445 1.045 ;
        RECT  8.085 0.345 8.375 0.465 ;
        RECT  8.085 0.700 8.375 0.820 ;
        RECT  8.015 0.185 8.085 0.465 ;
        RECT  8.015 0.700 8.085 1.045 ;
        RECT  7.725 0.345 8.015 0.465 ;
        RECT  7.725 0.700 8.015 0.820 ;
        RECT  7.655 0.185 7.725 0.465 ;
        RECT  7.655 0.700 7.725 1.045 ;
        RECT  7.365 0.345 7.655 0.465 ;
        RECT  7.365 0.700 7.655 0.820 ;
        RECT  7.295 0.185 7.365 0.465 ;
        RECT  7.295 0.700 7.365 1.045 ;
        RECT  7.005 0.345 7.295 0.465 ;
        RECT  7.005 0.700 7.295 0.820 ;
        RECT  6.935 0.185 7.005 0.465 ;
        RECT  6.935 0.700 7.005 1.045 ;
        RECT  6.645 0.345 6.935 0.465 ;
        RECT  6.645 0.700 6.935 0.820 ;
        RECT  6.575 0.185 6.645 0.465 ;
        RECT  6.575 0.700 6.645 1.045 ;
        RECT  6.475 0.345 6.575 0.465 ;
        RECT  6.475 0.700 6.575 0.820 ;
        RECT  6.285 0.345 6.475 0.820 ;
        RECT  6.215 0.185 6.285 1.045 ;
        RECT  6.125 0.345 6.215 0.820 ;
        RECT  5.925 0.345 6.125 0.465 ;
        RECT  5.925 0.700 6.125 0.820 ;
        RECT  5.855 0.185 5.925 0.465 ;
        RECT  5.855 0.700 5.925 1.045 ;
        RECT  5.545 0.345 5.855 0.465 ;
        RECT  5.565 0.700 5.855 0.820 ;
        RECT  5.495 0.700 5.565 1.045 ;
        RECT  5.475 0.185 5.545 0.465 ;
        RECT  5.205 0.700 5.495 0.820 ;
        RECT  5.165 0.345 5.475 0.465 ;
        RECT  5.135 0.700 5.205 1.045 ;
        RECT  5.095 0.185 5.165 0.465 ;
        RECT  4.845 0.700 5.135 0.820 ;
        RECT  4.785 0.345 5.095 0.465 ;
        RECT  4.775 0.700 4.845 1.045 ;
        RECT  4.715 0.185 4.785 0.465 ;
        RECT  4.485 0.700 4.775 0.820 ;
        RECT  4.405 0.345 4.715 0.465 ;
        RECT  4.415 0.700 4.485 1.045 ;
        RECT  4.335 0.185 4.405 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.1274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.495 4.055 0.795 ;
        RECT  3.360 0.725 3.955 0.795 ;
        RECT  3.240 0.545 3.360 0.795 ;
        RECT  2.690 0.725 3.240 0.795 ;
        RECT  2.570 0.545 2.690 0.795 ;
        RECT  2.535 0.725 2.570 0.795 ;
        RECT  2.465 0.725 2.535 0.960 ;
        RECT  1.960 0.890 2.465 0.960 ;
        RECT  1.890 0.695 1.960 0.960 ;
        RECT  1.790 0.695 1.890 0.765 ;
        RECT  1.700 0.495 1.790 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.625 -0.115 8.680 0.115 ;
        RECT  8.555 -0.115 8.625 0.475 ;
        RECT  8.290 -0.115 8.555 0.115 ;
        RECT  8.170 -0.115 8.290 0.275 ;
        RECT  7.930 -0.115 8.170 0.115 ;
        RECT  7.810 -0.115 7.930 0.275 ;
        RECT  7.570 -0.115 7.810 0.115 ;
        RECT  7.450 -0.115 7.570 0.275 ;
        RECT  7.210 -0.115 7.450 0.115 ;
        RECT  7.090 -0.115 7.210 0.275 ;
        RECT  6.850 -0.115 7.090 0.115 ;
        RECT  6.730 -0.115 6.850 0.275 ;
        RECT  6.490 -0.115 6.730 0.115 ;
        RECT  6.370 -0.115 6.490 0.275 ;
        RECT  6.130 -0.115 6.370 0.115 ;
        RECT  6.010 -0.115 6.130 0.275 ;
        RECT  5.760 -0.115 6.010 0.115 ;
        RECT  5.640 -0.115 5.760 0.275 ;
        RECT  5.380 -0.115 5.640 0.115 ;
        RECT  5.260 -0.115 5.380 0.275 ;
        RECT  5.000 -0.115 5.260 0.115 ;
        RECT  4.880 -0.115 5.000 0.275 ;
        RECT  4.620 -0.115 4.880 0.115 ;
        RECT  4.500 -0.115 4.620 0.275 ;
        RECT  2.285 -0.115 4.500 0.115 ;
        RECT  2.215 -0.115 2.285 0.305 ;
        RECT  1.025 -0.115 2.215 0.115 ;
        RECT  0.955 -0.115 1.025 0.290 ;
        RECT  0.300 -0.115 0.955 0.115 ;
        RECT  0.230 -0.115 0.300 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.625 1.145 8.680 1.375 ;
        RECT  8.555 0.675 8.625 1.375 ;
        RECT  8.290 1.145 8.555 1.375 ;
        RECT  8.170 0.890 8.290 1.375 ;
        RECT  7.930 1.145 8.170 1.375 ;
        RECT  7.810 0.890 7.930 1.375 ;
        RECT  7.570 1.145 7.810 1.375 ;
        RECT  7.450 0.890 7.570 1.375 ;
        RECT  7.210 1.145 7.450 1.375 ;
        RECT  7.090 0.890 7.210 1.375 ;
        RECT  6.850 1.145 7.090 1.375 ;
        RECT  6.730 0.890 6.850 1.375 ;
        RECT  6.490 1.145 6.730 1.375 ;
        RECT  6.370 0.890 6.490 1.375 ;
        RECT  6.130 1.145 6.370 1.375 ;
        RECT  6.010 0.890 6.130 1.375 ;
        RECT  5.770 1.145 6.010 1.375 ;
        RECT  5.650 0.890 5.770 1.375 ;
        RECT  5.410 1.145 5.650 1.375 ;
        RECT  5.290 0.890 5.410 1.375 ;
        RECT  5.050 1.145 5.290 1.375 ;
        RECT  4.930 0.890 5.050 1.375 ;
        RECT  4.690 1.145 4.930 1.375 ;
        RECT  4.570 0.890 4.690 1.375 ;
        RECT  4.330 1.145 4.570 1.375 ;
        RECT  4.210 1.020 4.330 1.375 ;
        RECT  3.790 1.145 4.210 1.375 ;
        RECT  3.670 1.005 3.790 1.375 ;
        RECT  3.070 1.145 3.670 1.375 ;
        RECT  2.950 1.005 3.070 1.375 ;
        RECT  2.350 1.145 2.950 1.375 ;
        RECT  2.230 1.030 2.350 1.375 ;
        RECT  1.630 1.145 2.230 1.375 ;
        RECT  1.510 1.010 1.630 1.375 ;
        RECT  1.080 1.145 1.510 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.375 0.185 8.445 0.465 ;
        RECT  8.375 0.700 8.445 1.045 ;
        RECT  8.085 0.345 8.375 0.465 ;
        RECT  8.085 0.700 8.375 0.820 ;
        RECT  8.015 0.185 8.085 0.465 ;
        RECT  8.015 0.700 8.085 1.045 ;
        RECT  7.725 0.345 8.015 0.465 ;
        RECT  7.725 0.700 8.015 0.820 ;
        RECT  7.655 0.185 7.725 0.465 ;
        RECT  7.655 0.700 7.725 1.045 ;
        RECT  7.365 0.345 7.655 0.465 ;
        RECT  7.365 0.700 7.655 0.820 ;
        RECT  7.295 0.185 7.365 0.465 ;
        RECT  7.295 0.700 7.365 1.045 ;
        RECT  7.005 0.345 7.295 0.465 ;
        RECT  7.005 0.700 7.295 0.820 ;
        RECT  6.935 0.185 7.005 0.465 ;
        RECT  6.935 0.700 7.005 1.045 ;
        RECT  6.645 0.345 6.935 0.465 ;
        RECT  6.645 0.700 6.935 0.820 ;
        RECT  6.575 0.185 6.645 0.465 ;
        RECT  6.575 0.700 6.645 1.045 ;
        RECT  6.545 0.345 6.575 0.465 ;
        RECT  6.545 0.700 6.575 0.820 ;
        RECT  5.925 0.345 6.055 0.465 ;
        RECT  5.925 0.700 6.055 0.820 ;
        RECT  5.855 0.185 5.925 0.465 ;
        RECT  5.855 0.700 5.925 1.045 ;
        RECT  5.545 0.345 5.855 0.465 ;
        RECT  5.565 0.700 5.855 0.820 ;
        RECT  5.495 0.700 5.565 1.045 ;
        RECT  5.475 0.185 5.545 0.465 ;
        RECT  5.205 0.700 5.495 0.820 ;
        RECT  5.165 0.345 5.475 0.465 ;
        RECT  5.135 0.700 5.205 1.045 ;
        RECT  5.095 0.185 5.165 0.465 ;
        RECT  4.845 0.700 5.135 0.820 ;
        RECT  4.785 0.345 5.095 0.465 ;
        RECT  4.775 0.700 4.845 1.045 ;
        RECT  4.715 0.185 4.785 0.465 ;
        RECT  4.485 0.700 4.775 0.820 ;
        RECT  4.405 0.345 4.715 0.465 ;
        RECT  4.415 0.700 4.485 1.045 ;
        RECT  4.335 0.185 4.405 0.465 ;
        RECT  6.575 0.545 8.415 0.615 ;
        RECT  4.205 0.545 6.025 0.615 ;
        RECT  4.135 0.215 4.205 0.935 ;
        RECT  2.370 0.215 4.135 0.285 ;
        RECT  3.430 0.865 4.135 0.935 ;
        RECT  3.670 0.395 3.750 0.640 ;
        RECT  3.035 0.395 3.670 0.465 ;
        RECT  3.310 0.865 3.430 1.075 ;
        RECT  2.685 0.865 3.310 0.935 ;
        RECT  2.965 0.395 3.035 0.640 ;
        RECT  2.395 0.395 2.965 0.465 ;
        RECT  2.615 0.865 2.685 1.035 ;
        RECT  2.325 0.395 2.395 0.820 ;
        RECT  2.105 0.395 2.325 0.465 ;
        RECT  2.050 0.750 2.325 0.820 ;
        RECT  1.940 0.545 2.140 0.615 ;
        RECT  2.035 0.185 2.105 0.465 ;
        RECT  1.870 0.210 1.940 0.615 ;
        RECT  1.230 0.210 1.870 0.280 ;
        RECT  1.715 0.835 1.785 1.050 ;
        RECT  1.590 0.355 1.770 0.425 ;
        RECT  1.590 0.835 1.715 0.905 ;
        RECT  1.520 0.355 1.590 0.905 ;
        RECT  1.470 0.690 1.520 0.810 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.360 1.400 1.050 ;
        RECT  1.330 0.360 1.355 0.950 ;
        RECT  1.300 0.360 1.330 0.460 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.230 0.680 1.240 0.800 ;
        RECT  1.160 0.210 1.230 0.800 ;
        RECT  1.110 0.210 1.160 0.280 ;
        RECT  0.955 0.730 1.160 0.800 ;
        RECT  1.020 0.370 1.090 0.550 ;
        RECT  0.770 0.370 1.020 0.440 ;
        RECT  0.885 0.620 0.955 0.800 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.185 0.770 0.800 ;
        RECT  0.580 0.185 0.700 0.285 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.525 0.355 0.590 0.640 ;
        RECT  0.520 0.355 0.525 1.055 ;
        RECT  0.455 0.570 0.520 1.055 ;
        RECT  0.440 0.195 0.510 0.265 ;
        RECT  0.370 0.195 0.440 0.415 ;
        RECT  0.125 0.345 0.370 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD24BWP

MACRO CKLHQD2BWP
    CLASS CORE ;
    FOREIGN CKLHQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.355 3.045 0.905 ;
        RECT  2.975 0.185 2.985 1.045 ;
        RECT  2.915 0.185 2.975 0.465 ;
        RECT  2.915 0.785 2.975 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 1.795 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.300 ;
        RECT  2.790 -0.115 3.095 0.115 ;
        RECT  2.710 -0.115 2.790 0.450 ;
        RECT  1.045 -0.115 2.710 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 1.145 3.220 1.375 ;
        RECT  3.095 0.960 3.165 1.375 ;
        RECT  2.810 1.145 3.095 1.375 ;
        RECT  2.690 1.005 2.810 1.375 ;
        RECT  2.410 1.145 2.690 1.375 ;
        RECT  2.290 1.000 2.410 1.375 ;
        RECT  1.650 1.145 2.290 1.375 ;
        RECT  1.530 1.000 1.650 1.375 ;
        RECT  1.100 1.145 1.530 1.375 ;
        RECT  0.980 1.020 1.100 1.375 ;
        RECT  0.130 1.145 0.980 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.775 0.520 2.845 0.920 ;
        RECT  2.025 0.850 2.775 0.920 ;
        RECT  2.540 0.330 2.610 0.780 ;
        RECT  2.515 0.330 2.540 0.450 ;
        RECT  2.275 0.710 2.540 0.780 ;
        RECT  2.425 0.520 2.470 0.640 ;
        RECT  2.355 0.195 2.425 0.640 ;
        RECT  1.270 0.195 2.355 0.265 ;
        RECT  2.205 0.520 2.275 0.780 ;
        RECT  2.025 0.355 2.230 0.425 ;
        RECT  1.955 0.355 2.025 1.035 ;
        RECT  1.585 0.355 1.850 0.425 ;
        RECT  1.755 0.860 1.825 1.035 ;
        RECT  1.585 0.860 1.755 0.930 ;
        RECT  1.515 0.355 1.585 0.930 ;
        RECT  1.500 0.665 1.515 0.785 ;
        RECT  1.410 0.885 1.445 1.025 ;
        RECT  1.340 0.345 1.410 1.025 ;
        RECT  0.835 0.880 1.340 0.950 ;
        RECT  1.200 0.195 1.270 0.810 ;
        RECT  1.130 0.195 1.200 0.265 ;
        RECT  0.935 0.740 1.200 0.810 ;
        RECT  1.060 0.370 1.130 0.640 ;
        RECT  0.770 0.370 1.060 0.440 ;
        RECT  0.865 0.520 0.935 0.810 ;
        RECT  0.765 0.880 0.835 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.525 0.985 0.765 1.055 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.345 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD2BWP

MACRO CKLHQD3BWP
    CLASS CORE ;
    FOREIGN CKLHQD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.185 3.305 0.485 ;
        RECT  3.235 0.700 3.305 1.035 ;
        RECT  3.115 0.355 3.235 0.485 ;
        RECT  3.115 0.700 3.235 0.820 ;
        RECT  2.945 0.355 3.115 0.820 ;
        RECT  2.905 0.185 2.945 1.035 ;
        RECT  2.875 0.185 2.905 0.485 ;
        RECT  2.875 0.700 2.905 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0370 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 1.795 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 -0.115 3.360 0.115 ;
        RECT  3.030 -0.115 3.150 0.280 ;
        RECT  2.770 -0.115 3.030 0.115 ;
        RECT  2.690 -0.115 2.770 0.440 ;
        RECT  1.045 -0.115 2.690 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.145 3.360 1.375 ;
        RECT  3.030 0.890 3.150 1.375 ;
        RECT  2.790 1.145 3.030 1.375 ;
        RECT  2.670 1.005 2.790 1.375 ;
        RECT  2.390 1.145 2.670 1.375 ;
        RECT  2.270 1.005 2.390 1.375 ;
        RECT  1.660 1.145 2.270 1.375 ;
        RECT  1.540 1.000 1.660 1.375 ;
        RECT  1.100 1.145 1.540 1.375 ;
        RECT  0.980 1.020 1.100 1.375 ;
        RECT  0.130 1.145 0.980 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.235 0.185 3.305 0.485 ;
        RECT  3.235 0.700 3.305 1.035 ;
        RECT  3.185 0.355 3.235 0.485 ;
        RECT  3.185 0.700 3.235 0.820 ;
        RECT  2.735 0.510 2.805 0.935 ;
        RECT  2.005 0.865 2.735 0.935 ;
        RECT  2.530 0.330 2.600 0.795 ;
        RECT  2.495 0.330 2.530 0.450 ;
        RECT  2.255 0.725 2.530 0.795 ;
        RECT  2.425 0.520 2.455 0.640 ;
        RECT  2.355 0.195 2.425 0.640 ;
        RECT  1.270 0.195 2.355 0.265 ;
        RECT  2.185 0.520 2.255 0.795 ;
        RECT  2.005 0.355 2.210 0.425 ;
        RECT  1.935 0.355 2.005 1.035 ;
        RECT  1.585 0.355 1.850 0.425 ;
        RECT  1.755 0.860 1.825 1.035 ;
        RECT  1.585 0.860 1.755 0.930 ;
        RECT  1.515 0.355 1.585 0.930 ;
        RECT  1.500 0.520 1.515 0.640 ;
        RECT  1.410 0.885 1.445 1.025 ;
        RECT  1.340 0.345 1.410 1.025 ;
        RECT  0.835 0.880 1.340 0.950 ;
        RECT  1.200 0.195 1.270 0.810 ;
        RECT  1.130 0.195 1.200 0.265 ;
        RECT  0.935 0.740 1.200 0.810 ;
        RECT  1.060 0.370 1.130 0.640 ;
        RECT  0.770 0.370 1.060 0.440 ;
        RECT  0.865 0.520 0.935 0.810 ;
        RECT  0.765 0.880 0.835 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.525 0.985 0.765 1.055 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.345 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD3BWP

MACRO CKLHQD4BWP
    CLASS CORE ;
    FOREIGN CKLHQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.455 0.185 3.530 0.465 ;
        RECT  3.455 0.700 3.525 1.035 ;
        RECT  3.395 0.355 3.455 0.465 ;
        RECT  3.395 0.700 3.455 0.820 ;
        RECT  3.185 0.355 3.395 0.820 ;
        RECT  3.145 0.355 3.185 0.465 ;
        RECT  3.145 0.700 3.185 0.820 ;
        RECT  3.075 0.185 3.145 0.465 ;
        RECT  3.075 0.700 3.145 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0596 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.545 2.605 0.615 ;
        RECT  2.365 0.545 2.435 0.920 ;
        RECT  1.790 0.850 2.365 0.920 ;
        RECT  1.700 0.495 1.790 0.920 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.705 -0.115 3.780 0.115 ;
        RECT  3.635 -0.115 3.705 0.465 ;
        RECT  3.360 -0.115 3.635 0.115 ;
        RECT  3.240 -0.115 3.360 0.280 ;
        RECT  1.045 -0.115 3.240 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.705 1.145 3.780 1.375 ;
        RECT  3.635 0.675 3.705 1.375 ;
        RECT  3.360 1.145 3.635 1.375 ;
        RECT  3.240 0.890 3.360 1.375 ;
        RECT  2.960 1.145 3.240 1.375 ;
        RECT  2.880 0.860 2.960 1.375 ;
        RECT  1.100 1.145 2.880 1.375 ;
        RECT  0.980 1.020 1.100 1.375 ;
        RECT  0.130 1.145 0.980 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.185 3.530 0.465 ;
        RECT  3.465 0.700 3.525 1.035 ;
        RECT  3.075 0.185 3.115 0.465 ;
        RECT  3.075 0.700 3.115 1.045 ;
        RECT  2.995 0.545 3.070 0.615 ;
        RECT  2.925 0.245 2.995 0.790 ;
        RECT  2.290 0.245 2.925 0.315 ;
        RECT  2.585 0.720 2.925 0.790 ;
        RECT  2.765 0.395 2.835 0.640 ;
        RECT  2.295 0.395 2.765 0.465 ;
        RECT  2.515 0.720 2.585 1.035 ;
        RECT  2.225 0.395 2.295 0.780 ;
        RECT  1.950 0.710 2.225 0.780 ;
        RECT  2.030 0.195 2.100 0.640 ;
        RECT  1.260 0.195 2.030 0.265 ;
        RECT  1.950 0.350 1.960 0.470 ;
        RECT  1.880 0.350 1.950 0.780 ;
        RECT  1.590 0.990 1.850 1.060 ;
        RECT  1.590 0.345 1.810 0.415 ;
        RECT  1.520 0.345 1.590 1.060 ;
        RECT  1.470 0.520 1.520 0.640 ;
        RECT  1.400 0.880 1.445 1.050 ;
        RECT  1.375 0.355 1.400 1.050 ;
        RECT  1.330 0.355 1.375 0.950 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.190 0.195 1.260 0.800 ;
        RECT  1.130 0.195 1.190 0.265 ;
        RECT  0.955 0.730 1.190 0.800 ;
        RECT  1.050 0.370 1.120 0.550 ;
        RECT  0.770 0.370 1.050 0.440 ;
        RECT  0.885 0.620 0.955 0.800 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.345 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD4BWP

MACRO CKLHQD6BWP
    CLASS CORE ;
    FOREIGN CKLHQD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.3024 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.755 0.700 3.825 1.035 ;
        RECT  3.535 0.335 3.755 0.465 ;
        RECT  3.535 0.700 3.755 0.820 ;
        RECT  3.465 0.335 3.535 0.820 ;
        RECT  3.395 0.185 3.465 1.035 ;
        RECT  3.325 0.335 3.395 0.820 ;
        RECT  3.105 0.335 3.325 0.465 ;
        RECT  3.105 0.700 3.325 0.820 ;
        RECT  3.035 0.185 3.105 0.465 ;
        RECT  3.035 0.700 3.105 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0596 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.545 2.565 0.615 ;
        RECT  2.345 0.545 2.415 0.920 ;
        RECT  1.790 0.850 2.345 0.920 ;
        RECT  1.700 0.550 1.790 0.920 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.465 ;
        RECT  3.670 -0.115 3.935 0.115 ;
        RECT  3.550 -0.115 3.670 0.255 ;
        RECT  3.310 -0.115 3.550 0.115 ;
        RECT  3.190 -0.115 3.310 0.255 ;
        RECT  1.045 -0.115 3.190 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.145 4.060 1.375 ;
        RECT  3.935 0.685 4.005 1.375 ;
        RECT  3.670 1.145 3.935 1.375 ;
        RECT  3.550 0.890 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 0.890 3.310 1.375 ;
        RECT  2.930 1.145 3.190 1.375 ;
        RECT  2.850 0.860 2.930 1.375 ;
        RECT  1.080 1.145 2.850 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.755 0.185 3.825 0.465 ;
        RECT  3.755 0.700 3.825 1.035 ;
        RECT  3.605 0.335 3.755 0.465 ;
        RECT  3.605 0.700 3.755 0.820 ;
        RECT  3.105 0.335 3.255 0.465 ;
        RECT  3.105 0.700 3.255 0.820 ;
        RECT  3.035 0.185 3.105 0.465 ;
        RECT  3.035 0.700 3.105 1.035 ;
        RECT  3.630 0.545 3.960 0.615 ;
        RECT  2.955 0.545 3.225 0.615 ;
        RECT  2.885 0.245 2.955 0.790 ;
        RECT  2.250 0.245 2.885 0.315 ;
        RECT  2.565 0.720 2.885 0.790 ;
        RECT  2.745 0.395 2.815 0.640 ;
        RECT  2.275 0.395 2.745 0.465 ;
        RECT  2.495 0.720 2.565 1.035 ;
        RECT  2.205 0.395 2.275 0.780 ;
        RECT  1.940 0.710 2.205 0.780 ;
        RECT  2.050 0.210 2.120 0.640 ;
        RECT  1.260 0.210 2.050 0.280 ;
        RECT  2.010 0.515 2.050 0.640 ;
        RECT  1.940 0.350 1.980 0.450 ;
        RECT  1.870 0.350 1.940 0.780 ;
        RECT  1.590 0.990 1.830 1.060 ;
        RECT  1.715 0.360 1.785 0.480 ;
        RECT  1.590 0.410 1.715 0.480 ;
        RECT  1.520 0.410 1.590 1.060 ;
        RECT  1.470 0.520 1.520 0.640 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.360 1.400 1.050 ;
        RECT  1.330 0.360 1.355 0.950 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.190 0.210 1.260 0.800 ;
        RECT  1.130 0.210 1.190 0.280 ;
        RECT  1.175 0.680 1.190 0.800 ;
        RECT  0.955 0.680 1.175 0.750 ;
        RECT  1.050 0.370 1.120 0.550 ;
        RECT  0.770 0.370 1.050 0.440 ;
        RECT  0.885 0.620 0.955 0.750 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.335 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD6BWP

MACRO CKLHQD8BWP
    CLASS CORE ;
    FOREIGN CKLHQD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.175 0.185 4.245 0.465 ;
        RECT  4.175 0.700 4.245 1.035 ;
        RECT  3.885 0.355 4.175 0.465 ;
        RECT  3.885 0.700 4.175 0.820 ;
        RECT  3.815 0.185 3.885 0.465 ;
        RECT  3.815 0.700 3.885 1.045 ;
        RECT  3.525 0.355 3.815 0.820 ;
        RECT  3.465 0.185 3.525 1.045 ;
        RECT  3.455 0.185 3.465 0.465 ;
        RECT  3.435 0.700 3.465 1.045 ;
        RECT  3.145 0.355 3.455 0.465 ;
        RECT  3.145 0.700 3.435 0.820 ;
        RECT  3.075 0.185 3.145 0.465 ;
        RECT  3.075 0.700 3.145 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.495 0.385 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.0596 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.545 2.605 0.615 ;
        RECT  2.365 0.545 2.435 0.925 ;
        RECT  1.790 0.855 2.365 0.925 ;
        RECT  1.700 0.550 1.790 0.925 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 -0.115 4.480 0.115 ;
        RECT  4.355 -0.115 4.425 0.465 ;
        RECT  4.090 -0.115 4.355 0.115 ;
        RECT  3.970 -0.115 4.090 0.275 ;
        RECT  3.730 -0.115 3.970 0.115 ;
        RECT  3.610 -0.115 3.730 0.275 ;
        RECT  3.360 -0.115 3.610 0.115 ;
        RECT  3.240 -0.115 3.360 0.275 ;
        RECT  1.045 -0.115 3.240 0.115 ;
        RECT  0.975 -0.115 1.045 0.290 ;
        RECT  0.310 -0.115 0.975 0.115 ;
        RECT  0.230 -0.115 0.310 0.265 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 1.145 4.480 1.375 ;
        RECT  4.355 0.675 4.425 1.375 ;
        RECT  4.090 1.145 4.355 1.375 ;
        RECT  3.970 0.890 4.090 1.375 ;
        RECT  3.730 1.145 3.970 1.375 ;
        RECT  3.610 0.890 3.730 1.375 ;
        RECT  3.360 1.145 3.610 1.375 ;
        RECT  3.240 0.890 3.360 1.375 ;
        RECT  2.955 1.145 3.240 1.375 ;
        RECT  2.885 0.860 2.955 1.375 ;
        RECT  1.080 1.145 2.885 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.130 1.145 0.960 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.175 0.185 4.245 0.465 ;
        RECT  4.175 0.700 4.245 1.035 ;
        RECT  3.885 0.355 4.175 0.465 ;
        RECT  3.885 0.700 4.175 0.820 ;
        RECT  3.145 0.355 3.395 0.465 ;
        RECT  3.145 0.700 3.395 0.820 ;
        RECT  3.075 0.185 3.145 0.465 ;
        RECT  3.075 0.700 3.145 1.035 ;
        RECT  3.915 0.545 4.255 0.615 ;
        RECT  2.975 0.545 3.365 0.615 ;
        RECT  2.905 0.245 2.975 0.790 ;
        RECT  2.290 0.245 2.905 0.315 ;
        RECT  2.585 0.720 2.905 0.790 ;
        RECT  2.765 0.395 2.835 0.640 ;
        RECT  2.295 0.395 2.765 0.465 ;
        RECT  2.515 0.720 2.585 1.035 ;
        RECT  2.225 0.395 2.295 0.785 ;
        RECT  1.965 0.715 2.225 0.785 ;
        RECT  2.075 0.210 2.145 0.640 ;
        RECT  1.260 0.210 2.075 0.280 ;
        RECT  2.040 0.520 2.075 0.640 ;
        RECT  1.895 0.350 1.965 0.785 ;
        RECT  1.590 0.995 1.870 1.065 ;
        RECT  1.715 0.360 1.785 0.480 ;
        RECT  1.590 0.410 1.715 0.480 ;
        RECT  1.520 0.410 1.590 1.065 ;
        RECT  1.470 0.520 1.520 0.640 ;
        RECT  1.400 0.880 1.425 1.050 ;
        RECT  1.355 0.360 1.400 1.050 ;
        RECT  1.330 0.360 1.355 0.950 ;
        RECT  0.855 0.880 1.330 0.950 ;
        RECT  1.190 0.210 1.260 0.800 ;
        RECT  1.130 0.210 1.190 0.280 ;
        RECT  1.175 0.680 1.190 0.800 ;
        RECT  0.955 0.680 1.175 0.750 ;
        RECT  1.050 0.370 1.120 0.550 ;
        RECT  0.770 0.370 1.050 0.440 ;
        RECT  0.885 0.610 0.955 0.750 ;
        RECT  0.785 0.880 0.855 1.055 ;
        RECT  0.525 0.985 0.785 1.055 ;
        RECT  0.700 0.195 0.770 0.800 ;
        RECT  0.590 0.195 0.700 0.265 ;
        RECT  0.685 0.730 0.700 0.800 ;
        RECT  0.615 0.730 0.685 0.905 ;
        RECT  0.530 0.335 0.600 0.640 ;
        RECT  0.525 0.570 0.530 0.640 ;
        RECT  0.455 0.570 0.525 1.055 ;
        RECT  0.450 0.195 0.510 0.265 ;
        RECT  0.380 0.195 0.450 0.415 ;
        RECT  0.125 0.345 0.380 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD8BWP

MACRO CKLNQD12BWP
    CLASS CORE ;
    FOREIGN CKLNQD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.5712 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.730 0.185 4.810 0.465 ;
        RECT  4.730 0.725 4.810 1.025 ;
        RECT  4.430 0.345 4.730 0.465 ;
        RECT  4.430 0.725 4.730 0.920 ;
        RECT  4.350 0.185 4.430 0.465 ;
        RECT  4.350 0.725 4.430 1.025 ;
        RECT  4.095 0.345 4.350 0.465 ;
        RECT  4.095 0.725 4.350 0.920 ;
        RECT  4.050 0.345 4.095 0.920 ;
        RECT  3.970 0.185 4.050 1.045 ;
        RECT  3.955 0.185 3.970 0.920 ;
        RECT  3.745 0.345 3.955 0.920 ;
        RECT  3.670 0.345 3.745 0.465 ;
        RECT  3.670 0.725 3.745 0.920 ;
        RECT  3.590 0.185 3.670 0.465 ;
        RECT  3.590 0.725 3.670 1.025 ;
        RECT  3.310 0.345 3.590 0.465 ;
        RECT  3.310 0.725 3.590 0.920 ;
        RECT  3.230 0.185 3.310 0.465 ;
        RECT  3.230 0.725 3.310 1.025 ;
        RECT  2.950 0.345 3.230 0.465 ;
        RECT  2.950 0.725 3.230 0.920 ;
        RECT  2.875 0.185 2.950 0.465 ;
        RECT  2.870 0.725 2.950 1.025 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0568 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.610 2.345 0.770 ;
        RECT  1.810 0.700 2.275 0.770 ;
        RECT  1.715 0.495 1.810 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.440 ;
        RECT  4.640 -0.115 4.910 0.115 ;
        RECT  4.520 -0.115 4.640 0.275 ;
        RECT  4.260 -0.115 4.520 0.115 ;
        RECT  4.140 -0.115 4.260 0.275 ;
        RECT  3.880 -0.115 4.140 0.115 ;
        RECT  3.760 -0.115 3.880 0.275 ;
        RECT  3.510 -0.115 3.760 0.115 ;
        RECT  3.390 -0.115 3.510 0.275 ;
        RECT  3.150 -0.115 3.390 0.115 ;
        RECT  3.030 -0.115 3.150 0.275 ;
        RECT  2.790 -0.115 3.030 0.115 ;
        RECT  2.670 -0.115 2.790 0.250 ;
        RECT  1.150 -0.115 2.670 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.675 4.990 1.375 ;
        RECT  4.640 1.145 4.910 1.375 ;
        RECT  4.520 1.000 4.640 1.375 ;
        RECT  4.260 1.145 4.520 1.375 ;
        RECT  4.140 1.000 4.260 1.375 ;
        RECT  3.880 1.145 4.140 1.375 ;
        RECT  3.760 1.000 3.880 1.375 ;
        RECT  3.510 1.145 3.760 1.375 ;
        RECT  3.390 1.000 3.510 1.375 ;
        RECT  3.150 1.145 3.390 1.375 ;
        RECT  3.030 1.000 3.150 1.375 ;
        RECT  2.770 1.145 3.030 1.375 ;
        RECT  2.690 0.980 2.770 1.375 ;
        RECT  2.410 1.145 2.690 1.375 ;
        RECT  2.330 0.980 2.410 1.375 ;
        RECT  2.050 1.145 2.330 1.375 ;
        RECT  1.970 0.840 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.185 4.810 0.465 ;
        RECT  4.730 0.725 4.810 1.025 ;
        RECT  4.430 0.345 4.730 0.465 ;
        RECT  4.430 0.725 4.730 0.920 ;
        RECT  4.350 0.185 4.430 0.465 ;
        RECT  4.350 0.725 4.430 1.025 ;
        RECT  4.165 0.345 4.350 0.465 ;
        RECT  4.165 0.725 4.350 0.920 ;
        RECT  3.670 0.345 3.675 0.465 ;
        RECT  3.670 0.725 3.675 0.920 ;
        RECT  3.590 0.185 3.670 0.465 ;
        RECT  3.590 0.725 3.670 1.025 ;
        RECT  3.310 0.345 3.590 0.465 ;
        RECT  3.310 0.725 3.590 0.920 ;
        RECT  3.230 0.185 3.310 0.465 ;
        RECT  3.230 0.725 3.310 1.025 ;
        RECT  2.950 0.345 3.230 0.465 ;
        RECT  2.950 0.725 3.230 0.920 ;
        RECT  2.875 0.185 2.950 0.465 ;
        RECT  2.870 0.725 2.950 1.025 ;
        RECT  4.230 0.545 4.780 0.615 ;
        RECT  2.790 0.545 3.590 0.615 ;
        RECT  2.720 0.320 2.790 0.910 ;
        RECT  2.405 0.320 2.720 0.390 ;
        RECT  2.585 0.840 2.720 0.910 ;
        RECT  2.580 0.460 2.650 0.640 ;
        RECT  2.515 0.840 2.585 1.075 ;
        RECT  2.155 0.460 2.580 0.530 ;
        RECT  2.250 0.840 2.515 0.910 ;
        RECT  2.335 0.215 2.405 0.390 ;
        RECT  2.130 0.840 2.250 1.050 ;
        RECT  2.085 0.205 2.155 0.630 ;
        RECT  1.330 0.205 2.085 0.275 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD12BWP

MACRO CKLNQD16BWP
    CLASS CORE ;
    FOREIGN CKLNQD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.7616 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.720 6.030 0.950 ;
        RECT  5.930 0.185 6.010 0.465 ;
        RECT  5.650 0.345 5.930 0.465 ;
        RECT  5.570 0.185 5.650 0.465 ;
        RECT  5.290 0.345 5.570 0.465 ;
        RECT  5.210 0.185 5.290 0.465 ;
        RECT  4.935 0.345 5.210 0.465 ;
        RECT  4.930 0.345 4.935 0.950 ;
        RECT  4.850 0.185 4.930 0.950 ;
        RECT  4.585 0.345 4.850 0.950 ;
        RECT  4.570 0.345 4.585 0.465 ;
        RECT  3.390 0.715 4.585 0.950 ;
        RECT  4.490 0.185 4.570 0.465 ;
        RECT  4.210 0.345 4.490 0.465 ;
        RECT  4.130 0.185 4.210 0.465 ;
        RECT  3.850 0.345 4.130 0.465 ;
        RECT  3.770 0.185 3.850 0.465 ;
        RECT  3.490 0.345 3.770 0.465 ;
        RECT  3.410 0.185 3.490 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0214 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0780 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.945 0.510 3.015 0.770 ;
        RECT  2.375 0.700 2.945 0.770 ;
        RECT  2.275 0.530 2.375 0.770 ;
        RECT  1.810 0.700 2.275 0.770 ;
        RECT  1.715 0.495 1.810 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.185 -0.115 6.300 0.115 ;
        RECT  6.115 -0.115 6.185 0.440 ;
        RECT  5.850 -0.115 6.115 0.115 ;
        RECT  5.730 -0.115 5.850 0.275 ;
        RECT  5.490 -0.115 5.730 0.115 ;
        RECT  5.370 -0.115 5.490 0.275 ;
        RECT  5.130 -0.115 5.370 0.115 ;
        RECT  5.010 -0.115 5.130 0.275 ;
        RECT  4.770 -0.115 5.010 0.115 ;
        RECT  4.650 -0.115 4.770 0.275 ;
        RECT  4.410 -0.115 4.650 0.115 ;
        RECT  4.290 -0.115 4.410 0.275 ;
        RECT  4.050 -0.115 4.290 0.115 ;
        RECT  3.930 -0.115 4.050 0.275 ;
        RECT  3.690 -0.115 3.930 0.115 ;
        RECT  3.570 -0.115 3.690 0.275 ;
        RECT  3.305 -0.115 3.570 0.115 ;
        RECT  3.235 -0.115 3.305 0.440 ;
        RECT  1.125 -0.115 3.235 0.115 ;
        RECT  1.055 -0.115 1.125 0.285 ;
        RECT  0.340 -0.115 1.055 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.185 1.145 6.300 1.375 ;
        RECT  6.115 0.680 6.185 1.375 ;
        RECT  5.850 1.145 6.115 1.375 ;
        RECT  5.730 1.020 5.850 1.375 ;
        RECT  5.490 1.145 5.730 1.375 ;
        RECT  5.370 1.020 5.490 1.375 ;
        RECT  5.130 1.145 5.370 1.375 ;
        RECT  5.010 1.020 5.130 1.375 ;
        RECT  4.770 1.145 5.010 1.375 ;
        RECT  4.650 1.020 4.770 1.375 ;
        RECT  4.410 1.145 4.650 1.375 ;
        RECT  4.290 1.020 4.410 1.375 ;
        RECT  4.050 1.145 4.290 1.375 ;
        RECT  3.930 1.020 4.050 1.375 ;
        RECT  3.690 1.145 3.930 1.375 ;
        RECT  3.570 1.020 3.690 1.375 ;
        RECT  3.305 1.145 3.570 1.375 ;
        RECT  3.235 0.700 3.305 1.375 ;
        RECT  3.130 1.145 3.235 1.375 ;
        RECT  3.050 0.980 3.130 1.375 ;
        RECT  2.790 1.145 3.050 1.375 ;
        RECT  2.670 1.000 2.790 1.375 ;
        RECT  2.410 1.145 2.670 1.375 ;
        RECT  2.330 0.980 2.410 1.375 ;
        RECT  2.050 1.145 2.330 1.375 ;
        RECT  1.970 0.860 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.050 1.010 1.120 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.005 0.720 6.030 0.950 ;
        RECT  5.930 0.185 6.010 0.465 ;
        RECT  5.650 0.345 5.930 0.465 ;
        RECT  5.570 0.185 5.650 0.465 ;
        RECT  5.290 0.345 5.570 0.465 ;
        RECT  5.210 0.185 5.290 0.465 ;
        RECT  5.005 0.345 5.210 0.465 ;
        RECT  4.490 0.185 4.515 0.465 ;
        RECT  3.390 0.715 4.515 0.950 ;
        RECT  4.210 0.345 4.490 0.465 ;
        RECT  4.130 0.185 4.210 0.465 ;
        RECT  3.850 0.345 4.130 0.465 ;
        RECT  3.770 0.185 3.850 0.465 ;
        RECT  3.490 0.345 3.770 0.465 ;
        RECT  3.410 0.185 3.490 0.465 ;
        RECT  5.090 0.545 6.040 0.615 ;
        RECT  3.160 0.545 4.430 0.615 ;
        RECT  3.090 0.240 3.160 0.910 ;
        RECT  2.290 0.240 3.090 0.310 ;
        RECT  2.945 0.840 3.090 0.910 ;
        RECT  2.875 0.840 2.945 1.075 ;
        RECT  2.585 0.840 2.875 0.910 ;
        RECT  2.680 0.380 2.780 0.630 ;
        RECT  2.115 0.380 2.680 0.450 ;
        RECT  2.515 0.840 2.585 1.075 ;
        RECT  2.250 0.840 2.515 0.910 ;
        RECT  2.130 0.840 2.250 1.050 ;
        RECT  2.045 0.205 2.115 0.630 ;
        RECT  1.310 0.205 2.045 0.275 ;
        RECT  1.640 0.355 1.870 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.685 1.570 0.805 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.970 0.870 1.410 0.940 ;
        RECT  1.240 0.205 1.310 0.800 ;
        RECT  1.020 0.730 1.240 0.800 ;
        RECT  1.100 0.495 1.170 0.630 ;
        RECT  0.980 0.495 1.100 0.565 ;
        RECT  0.900 0.635 1.020 0.800 ;
        RECT  0.910 0.195 0.980 0.565 ;
        RECT  0.900 0.870 0.970 1.065 ;
        RECT  0.620 0.195 0.910 0.265 ;
        RECT  0.830 0.495 0.910 0.565 ;
        RECT  0.530 0.995 0.900 1.065 ;
        RECT  0.665 0.355 0.830 0.425 ;
        RECT  0.760 0.495 0.830 0.925 ;
        RECT  0.600 0.825 0.760 0.925 ;
        RECT  0.595 0.355 0.665 0.750 ;
        RECT  0.530 0.680 0.595 0.750 ;
        RECT  0.460 0.680 0.530 1.065 ;
        RECT  0.445 0.185 0.515 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD16BWP

MACRO CKLNQD1BWP
    CLASS CORE ;
    FOREIGN CKLNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.0748 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.325 2.625 1.045 ;
        RECT  2.535 0.325 2.555 0.455 ;
        RECT  2.535 0.760 2.555 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0360 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.115 2.660 0.115 ;
        RECT  2.360 -0.115 2.430 0.440 ;
        RECT  1.150 -0.115 2.360 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.145 2.660 1.375 ;
        RECT  2.320 0.980 2.440 1.375 ;
        RECT  2.070 1.145 2.320 1.375 ;
        RECT  1.950 0.980 2.070 1.375 ;
        RECT  1.700 1.145 1.950 1.375 ;
        RECT  1.580 0.985 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.460 0.520 2.485 0.640 ;
        RECT  2.390 0.520 2.460 0.910 ;
        RECT  2.225 0.840 2.390 0.910 ;
        RECT  2.220 0.205 2.290 0.640 ;
        RECT  2.155 0.840 2.225 1.075 ;
        RECT  1.330 0.205 2.220 0.275 ;
        RECT  2.045 0.840 2.155 0.910 ;
        RECT  1.975 0.345 2.045 0.910 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.845 1.865 1.050 ;
        RECT  1.640 0.845 1.795 0.915 ;
        RECT  1.570 0.355 1.640 0.915 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD1BWP

MACRO CKLNQD20BWP
    CLASS CORE ;
    FOREIGN CKLNQD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.9520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.720 7.010 0.950 ;
        RECT  6.910 0.185 6.990 0.465 ;
        RECT  6.630 0.345 6.910 0.465 ;
        RECT  6.550 0.185 6.630 0.465 ;
        RECT  6.270 0.345 6.550 0.465 ;
        RECT  6.190 0.185 6.270 0.465 ;
        RECT  5.910 0.345 6.190 0.465 ;
        RECT  5.830 0.185 5.910 0.465 ;
        RECT  5.550 0.345 5.830 0.465 ;
        RECT  5.495 0.185 5.550 0.465 ;
        RECT  5.470 0.185 5.495 0.950 ;
        RECT  5.190 0.345 5.470 0.950 ;
        RECT  5.145 0.185 5.190 0.950 ;
        RECT  5.110 0.185 5.145 0.465 ;
        RECT  3.650 0.720 5.145 0.950 ;
        RECT  4.830 0.345 5.110 0.465 ;
        RECT  4.750 0.185 4.830 0.465 ;
        RECT  4.470 0.345 4.750 0.465 ;
        RECT  4.390 0.185 4.470 0.465 ;
        RECT  4.110 0.345 4.390 0.465 ;
        RECT  4.030 0.185 4.110 0.465 ;
        RECT  3.750 0.345 4.030 0.465 ;
        RECT  3.670 0.185 3.750 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0992 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.065 0.635 3.185 0.770 ;
        RECT  2.345 0.700 3.065 0.770 ;
        RECT  2.275 0.520 2.345 0.770 ;
        RECT  1.810 0.700 2.275 0.770 ;
        RECT  1.715 0.495 1.810 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.165 -0.115 7.280 0.115 ;
        RECT  7.095 -0.115 7.165 0.440 ;
        RECT  6.830 -0.115 7.095 0.115 ;
        RECT  6.710 -0.115 6.830 0.275 ;
        RECT  6.470 -0.115 6.710 0.115 ;
        RECT  6.350 -0.115 6.470 0.275 ;
        RECT  6.110 -0.115 6.350 0.115 ;
        RECT  5.990 -0.115 6.110 0.275 ;
        RECT  5.750 -0.115 5.990 0.115 ;
        RECT  5.630 -0.115 5.750 0.275 ;
        RECT  5.390 -0.115 5.630 0.115 ;
        RECT  5.270 -0.115 5.390 0.275 ;
        RECT  5.030 -0.115 5.270 0.115 ;
        RECT  4.910 -0.115 5.030 0.275 ;
        RECT  4.670 -0.115 4.910 0.115 ;
        RECT  4.550 -0.115 4.670 0.275 ;
        RECT  4.310 -0.115 4.550 0.115 ;
        RECT  4.190 -0.115 4.310 0.275 ;
        RECT  3.950 -0.115 4.190 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.560 -0.115 3.830 0.115 ;
        RECT  3.440 -0.115 3.560 0.260 ;
        RECT  1.150 -0.115 3.440 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.165 1.145 7.280 1.375 ;
        RECT  7.095 0.675 7.165 1.375 ;
        RECT  6.830 1.145 7.095 1.375 ;
        RECT  6.710 1.020 6.830 1.375 ;
        RECT  6.470 1.145 6.710 1.375 ;
        RECT  6.350 1.020 6.470 1.375 ;
        RECT  6.110 1.145 6.350 1.375 ;
        RECT  5.990 1.020 6.110 1.375 ;
        RECT  5.750 1.145 5.990 1.375 ;
        RECT  5.630 1.020 5.750 1.375 ;
        RECT  5.390 1.145 5.630 1.375 ;
        RECT  5.270 1.020 5.390 1.375 ;
        RECT  5.030 1.145 5.270 1.375 ;
        RECT  4.910 1.020 5.030 1.375 ;
        RECT  4.670 1.145 4.910 1.375 ;
        RECT  4.550 1.020 4.670 1.375 ;
        RECT  4.310 1.145 4.550 1.375 ;
        RECT  4.190 1.020 4.310 1.375 ;
        RECT  3.950 1.145 4.190 1.375 ;
        RECT  3.830 1.020 3.950 1.375 ;
        RECT  3.560 1.145 3.830 1.375 ;
        RECT  3.440 1.000 3.560 1.375 ;
        RECT  3.160 1.145 3.440 1.375 ;
        RECT  3.040 1.000 3.160 1.375 ;
        RECT  2.790 1.145 3.040 1.375 ;
        RECT  2.670 1.000 2.790 1.375 ;
        RECT  2.410 1.145 2.670 1.375 ;
        RECT  2.330 0.980 2.410 1.375 ;
        RECT  2.050 1.145 2.330 1.375 ;
        RECT  1.970 0.840 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.720 7.010 0.950 ;
        RECT  6.910 0.185 6.990 0.465 ;
        RECT  6.630 0.345 6.910 0.465 ;
        RECT  6.550 0.185 6.630 0.465 ;
        RECT  6.270 0.345 6.550 0.465 ;
        RECT  6.190 0.185 6.270 0.465 ;
        RECT  5.910 0.345 6.190 0.465 ;
        RECT  5.830 0.185 5.910 0.465 ;
        RECT  5.565 0.345 5.830 0.465 ;
        RECT  4.830 0.345 5.075 0.465 ;
        RECT  3.650 0.720 5.075 0.950 ;
        RECT  4.750 0.185 4.830 0.465 ;
        RECT  4.470 0.345 4.750 0.465 ;
        RECT  4.390 0.185 4.470 0.465 ;
        RECT  4.110 0.345 4.390 0.465 ;
        RECT  4.030 0.185 4.110 0.465 ;
        RECT  3.750 0.345 4.030 0.465 ;
        RECT  3.670 0.185 3.750 0.465 ;
        RECT  5.690 0.545 7.030 0.615 ;
        RECT  3.570 0.545 5.010 0.615 ;
        RECT  3.500 0.330 3.570 0.910 ;
        RECT  3.300 0.330 3.500 0.400 ;
        RECT  3.325 0.840 3.500 0.910 ;
        RECT  3.100 0.485 3.420 0.555 ;
        RECT  3.255 0.840 3.325 1.075 ;
        RECT  3.230 0.230 3.300 0.400 ;
        RECT  2.945 0.840 3.255 0.910 ;
        RECT  2.310 0.230 3.230 0.300 ;
        RECT  3.030 0.370 3.100 0.555 ;
        RECT  2.780 0.370 3.030 0.440 ;
        RECT  2.875 0.840 2.945 1.075 ;
        RECT  2.585 0.840 2.875 0.910 ;
        RECT  2.680 0.370 2.780 0.630 ;
        RECT  2.115 0.370 2.680 0.440 ;
        RECT  2.515 0.840 2.585 1.075 ;
        RECT  2.250 0.840 2.515 0.910 ;
        RECT  2.130 0.840 2.250 1.050 ;
        RECT  2.045 0.205 2.115 0.630 ;
        RECT  1.330 0.205 2.045 0.275 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD20BWP

MACRO CKLNQD24BWP
    CLASS CORE ;
    FOREIGN CKLNQD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.1424 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.720 7.750 0.950 ;
        RECT  7.650 0.185 7.730 0.465 ;
        RECT  7.350 0.345 7.650 0.465 ;
        RECT  7.270 0.185 7.350 0.465 ;
        RECT  6.990 0.345 7.270 0.465 ;
        RECT  6.910 0.185 6.990 0.465 ;
        RECT  6.630 0.345 6.910 0.465 ;
        RECT  6.550 0.185 6.630 0.465 ;
        RECT  6.270 0.345 6.550 0.465 ;
        RECT  6.190 0.185 6.270 0.465 ;
        RECT  5.910 0.345 6.190 0.465 ;
        RECT  5.830 0.185 5.910 0.465 ;
        RECT  5.550 0.345 5.830 0.465 ;
        RECT  5.495 0.185 5.550 0.465 ;
        RECT  5.470 0.185 5.495 0.950 ;
        RECT  5.190 0.345 5.470 0.950 ;
        RECT  5.145 0.185 5.190 0.950 ;
        RECT  5.110 0.185 5.145 0.465 ;
        RECT  3.630 0.720 5.145 0.950 ;
        RECT  4.830 0.345 5.110 0.465 ;
        RECT  4.750 0.185 4.830 0.465 ;
        RECT  4.470 0.345 4.750 0.465 ;
        RECT  4.390 0.185 4.470 0.465 ;
        RECT  4.110 0.345 4.390 0.465 ;
        RECT  4.030 0.185 4.110 0.465 ;
        RECT  3.730 0.345 4.030 0.465 ;
        RECT  3.650 0.185 3.730 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0992 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 0.635 3.200 0.770 ;
        RECT  2.485 0.700 3.080 0.770 ;
        RECT  2.415 0.520 2.485 0.770 ;
        RECT  1.810 0.700 2.415 0.770 ;
        RECT  1.715 0.495 1.810 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 -0.115 7.980 0.115 ;
        RECT  7.835 -0.115 7.905 0.440 ;
        RECT  7.560 -0.115 7.835 0.115 ;
        RECT  7.440 -0.115 7.560 0.275 ;
        RECT  7.190 -0.115 7.440 0.115 ;
        RECT  7.070 -0.115 7.190 0.275 ;
        RECT  6.830 -0.115 7.070 0.115 ;
        RECT  6.710 -0.115 6.830 0.275 ;
        RECT  6.470 -0.115 6.710 0.115 ;
        RECT  6.350 -0.115 6.470 0.275 ;
        RECT  6.110 -0.115 6.350 0.115 ;
        RECT  5.990 -0.115 6.110 0.275 ;
        RECT  5.750 -0.115 5.990 0.115 ;
        RECT  5.630 -0.115 5.750 0.275 ;
        RECT  5.390 -0.115 5.630 0.115 ;
        RECT  5.270 -0.115 5.390 0.275 ;
        RECT  5.030 -0.115 5.270 0.115 ;
        RECT  4.910 -0.115 5.030 0.275 ;
        RECT  4.670 -0.115 4.910 0.115 ;
        RECT  4.550 -0.115 4.670 0.275 ;
        RECT  4.310 -0.115 4.550 0.115 ;
        RECT  4.190 -0.115 4.310 0.275 ;
        RECT  3.940 -0.115 4.190 0.115 ;
        RECT  3.820 -0.115 3.940 0.275 ;
        RECT  3.560 -0.115 3.820 0.115 ;
        RECT  3.440 -0.115 3.560 0.240 ;
        RECT  1.150 -0.115 3.440 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 1.145 7.980 1.375 ;
        RECT  7.835 0.675 7.905 1.375 ;
        RECT  7.560 1.145 7.835 1.375 ;
        RECT  7.440 1.020 7.560 1.375 ;
        RECT  7.190 1.145 7.440 1.375 ;
        RECT  7.070 1.020 7.190 1.375 ;
        RECT  6.830 1.145 7.070 1.375 ;
        RECT  6.710 1.020 6.830 1.375 ;
        RECT  6.470 1.145 6.710 1.375 ;
        RECT  6.350 1.020 6.470 1.375 ;
        RECT  6.110 1.145 6.350 1.375 ;
        RECT  5.990 1.020 6.110 1.375 ;
        RECT  5.750 1.145 5.990 1.375 ;
        RECT  5.630 1.020 5.750 1.375 ;
        RECT  5.390 1.145 5.630 1.375 ;
        RECT  5.270 1.020 5.390 1.375 ;
        RECT  5.030 1.145 5.270 1.375 ;
        RECT  4.910 1.020 5.030 1.375 ;
        RECT  4.670 1.145 4.910 1.375 ;
        RECT  4.550 1.020 4.670 1.375 ;
        RECT  4.310 1.145 4.550 1.375 ;
        RECT  4.190 1.020 4.310 1.375 ;
        RECT  3.940 1.145 4.190 1.375 ;
        RECT  3.820 1.020 3.940 1.375 ;
        RECT  3.560 1.145 3.820 1.375 ;
        RECT  3.440 1.000 3.560 1.375 ;
        RECT  3.180 1.145 3.440 1.375 ;
        RECT  3.060 1.000 3.180 1.375 ;
        RECT  2.810 1.145 3.060 1.375 ;
        RECT  2.690 1.000 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.350 0.980 2.430 1.375 ;
        RECT  2.070 1.145 2.350 1.375 ;
        RECT  1.990 0.840 2.070 1.375 ;
        RECT  1.700 1.145 1.990 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.720 7.750 0.950 ;
        RECT  7.650 0.185 7.730 0.465 ;
        RECT  7.350 0.345 7.650 0.465 ;
        RECT  7.270 0.185 7.350 0.465 ;
        RECT  6.990 0.345 7.270 0.465 ;
        RECT  6.910 0.185 6.990 0.465 ;
        RECT  6.630 0.345 6.910 0.465 ;
        RECT  6.550 0.185 6.630 0.465 ;
        RECT  6.270 0.345 6.550 0.465 ;
        RECT  6.190 0.185 6.270 0.465 ;
        RECT  5.910 0.345 6.190 0.465 ;
        RECT  5.830 0.185 5.910 0.465 ;
        RECT  5.565 0.345 5.830 0.465 ;
        RECT  4.830 0.345 5.075 0.465 ;
        RECT  3.630 0.720 5.075 0.950 ;
        RECT  4.750 0.185 4.830 0.465 ;
        RECT  4.470 0.345 4.750 0.465 ;
        RECT  4.390 0.185 4.470 0.465 ;
        RECT  4.110 0.345 4.390 0.465 ;
        RECT  4.030 0.185 4.110 0.465 ;
        RECT  3.730 0.345 4.030 0.465 ;
        RECT  3.650 0.185 3.730 0.465 ;
        RECT  5.690 0.545 7.590 0.615 ;
        RECT  3.550 0.545 5.010 0.615 ;
        RECT  3.480 0.310 3.550 0.910 ;
        RECT  3.300 0.310 3.480 0.390 ;
        RECT  3.345 0.840 3.480 0.910 ;
        RECT  3.340 0.460 3.410 0.580 ;
        RECT  3.275 0.840 3.345 1.075 ;
        RECT  3.100 0.460 3.340 0.530 ;
        RECT  3.230 0.230 3.300 0.390 ;
        RECT  2.965 0.840 3.275 0.910 ;
        RECT  2.330 0.230 3.230 0.300 ;
        RECT  3.030 0.370 3.100 0.530 ;
        RECT  2.810 0.370 3.030 0.440 ;
        RECT  2.895 0.840 2.965 1.075 ;
        RECT  2.605 0.840 2.895 0.910 ;
        RECT  2.710 0.370 2.810 0.630 ;
        RECT  2.140 0.370 2.710 0.440 ;
        RECT  2.535 0.840 2.605 1.075 ;
        RECT  2.270 0.840 2.535 0.910 ;
        RECT  2.150 0.840 2.270 1.050 ;
        RECT  2.060 0.205 2.140 0.630 ;
        RECT  1.330 0.205 2.060 0.275 ;
        RECT  1.640 0.355 1.910 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD24BWP

MACRO CKLNQD2BWP
    CLASS CORE ;
    FOREIGN CKLNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.0952 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.565 0.355 2.625 0.905 ;
        RECT  2.555 0.200 2.565 1.045 ;
        RECT  2.495 0.200 2.555 0.430 ;
        RECT  2.495 0.785 2.555 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0214 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.300 ;
        RECT  2.390 -0.115 2.670 0.115 ;
        RECT  2.310 -0.115 2.390 0.380 ;
        RECT  1.125 -0.115 2.310 0.115 ;
        RECT  1.055 -0.115 1.125 0.285 ;
        RECT  0.340 -0.115 1.055 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.960 2.750 1.375 ;
        RECT  2.390 1.145 2.670 1.375 ;
        RECT  2.310 0.960 2.390 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.980 2.050 1.375 ;
        RECT  1.690 1.145 1.930 1.375 ;
        RECT  1.570 0.985 1.690 1.375 ;
        RECT  1.120 1.145 1.570 1.375 ;
        RECT  1.050 1.010 1.120 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.420 0.520 2.475 0.640 ;
        RECT  2.350 0.520 2.420 0.890 ;
        RECT  2.205 0.820 2.350 0.890 ;
        RECT  2.210 0.520 2.270 0.640 ;
        RECT  2.140 0.205 2.210 0.640 ;
        RECT  2.135 0.820 2.205 1.055 ;
        RECT  1.310 0.205 2.140 0.275 ;
        RECT  2.030 0.820 2.135 0.890 ;
        RECT  1.960 0.345 2.030 0.890 ;
        RECT  1.640 0.355 1.870 0.425 ;
        RECT  1.775 0.845 1.845 1.050 ;
        RECT  1.640 0.845 1.775 0.915 ;
        RECT  1.570 0.355 1.640 0.915 ;
        RECT  1.530 0.535 1.570 0.655 ;
        RECT  1.460 0.355 1.480 0.475 ;
        RECT  1.460 0.880 1.480 1.040 ;
        RECT  1.410 0.355 1.460 1.040 ;
        RECT  1.390 0.355 1.410 0.940 ;
        RECT  0.970 0.870 1.390 0.940 ;
        RECT  1.240 0.205 1.310 0.800 ;
        RECT  1.020 0.720 1.240 0.800 ;
        RECT  1.100 0.495 1.170 0.635 ;
        RECT  0.980 0.495 1.100 0.565 ;
        RECT  0.900 0.635 1.020 0.800 ;
        RECT  0.910 0.195 0.980 0.565 ;
        RECT  0.900 0.870 0.970 1.065 ;
        RECT  0.620 0.195 0.910 0.265 ;
        RECT  0.830 0.495 0.910 0.565 ;
        RECT  0.530 0.995 0.900 1.065 ;
        RECT  0.665 0.355 0.830 0.425 ;
        RECT  0.760 0.495 0.830 0.925 ;
        RECT  0.600 0.825 0.760 0.925 ;
        RECT  0.595 0.355 0.665 0.755 ;
        RECT  0.530 0.685 0.595 0.755 ;
        RECT  0.460 0.685 0.530 1.065 ;
        RECT  0.445 0.185 0.515 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD2BWP

MACRO CKLNQD3BWP
    CLASS CORE ;
    FOREIGN CKLNQD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.1836 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 0.290 3.030 0.465 ;
        RECT  2.950 0.700 3.030 1.050 ;
        RECT  2.845 0.375 2.950 0.465 ;
        RECT  2.845 0.700 2.950 0.820 ;
        RECT  2.635 0.375 2.845 0.820 ;
        RECT  2.600 0.375 2.635 0.465 ;
        RECT  2.600 0.700 2.635 0.820 ;
        RECT  2.520 0.290 2.600 0.465 ;
        RECT  2.520 0.700 2.600 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 3.080 0.115 ;
        RECT  2.720 -0.115 2.840 0.305 ;
        RECT  2.410 -0.115 2.720 0.115 ;
        RECT  2.330 -0.115 2.410 0.420 ;
        RECT  1.150 -0.115 2.330 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.145 3.080 1.375 ;
        RECT  2.720 0.890 2.840 1.375 ;
        RECT  2.430 1.145 2.720 1.375 ;
        RECT  2.310 0.980 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.970 0.960 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.985 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.290 3.030 0.465 ;
        RECT  2.950 0.700 3.030 1.050 ;
        RECT  2.905 0.375 2.950 0.465 ;
        RECT  2.905 0.700 2.950 0.820 ;
        RECT  2.520 0.290 2.575 0.465 ;
        RECT  2.520 0.700 2.575 1.050 ;
        RECT  2.440 0.540 2.555 0.620 ;
        RECT  2.370 0.540 2.440 0.890 ;
        RECT  2.225 0.820 2.370 0.890 ;
        RECT  2.230 0.520 2.290 0.640 ;
        RECT  2.160 0.205 2.230 0.640 ;
        RECT  2.155 0.820 2.225 1.055 ;
        RECT  1.330 0.205 2.160 0.275 ;
        RECT  2.050 0.820 2.155 0.890 ;
        RECT  1.970 0.345 2.050 0.890 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.845 1.865 1.050 ;
        RECT  1.640 0.845 1.795 0.915 ;
        RECT  1.570 0.355 1.640 0.915 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD3BWP

MACRO CKLNQD4BWP
    CLASS CORE ;
    FOREIGN CKLNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.2040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.915 0.280 2.990 0.465 ;
        RECT  2.915 0.700 2.990 1.045 ;
        RECT  2.835 0.365 2.915 0.465 ;
        RECT  2.835 0.700 2.915 0.820 ;
        RECT  2.625 0.365 2.835 0.820 ;
        RECT  2.595 0.365 2.625 0.465 ;
        RECT  2.595 0.700 2.625 0.820 ;
        RECT  2.525 0.280 2.595 0.465 ;
        RECT  2.525 0.700 2.595 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.490 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.295 ;
        RECT  2.410 -0.115 2.690 0.115 ;
        RECT  2.330 -0.115 2.410 0.410 ;
        RECT  1.160 -0.115 2.330 0.115 ;
        RECT  1.080 -0.115 1.160 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.675 3.170 1.375 ;
        RECT  2.820 1.145 3.090 1.375 ;
        RECT  2.700 0.890 2.820 1.375 ;
        RECT  2.430 1.145 2.700 1.375 ;
        RECT  2.310 0.980 2.430 1.375 ;
        RECT  2.070 1.145 2.310 1.375 ;
        RECT  1.950 0.980 2.070 1.375 ;
        RECT  1.700 1.145 1.950 1.375 ;
        RECT  1.580 0.985 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.915 0.280 2.990 0.465 ;
        RECT  2.915 0.700 2.990 1.045 ;
        RECT  2.905 0.365 2.915 0.465 ;
        RECT  2.905 0.700 2.915 0.820 ;
        RECT  2.525 0.280 2.555 0.465 ;
        RECT  2.525 0.700 2.555 1.045 ;
        RECT  2.440 0.540 2.535 0.620 ;
        RECT  2.370 0.540 2.440 0.890 ;
        RECT  2.225 0.820 2.370 0.890 ;
        RECT  2.230 0.520 2.290 0.640 ;
        RECT  2.160 0.205 2.230 0.640 ;
        RECT  2.155 0.820 2.225 1.055 ;
        RECT  1.330 0.205 2.160 0.275 ;
        RECT  2.050 0.820 2.155 0.890 ;
        RECT  1.970 0.345 2.050 0.890 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.845 1.865 1.050 ;
        RECT  1.640 0.845 1.795 0.915 ;
        RECT  1.570 0.355 1.640 0.915 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD4BWP

MACRO CKLNQD6BWP
    CLASS CORE ;
    FOREIGN CKLNQD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.2856 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.615 0.185 3.690 0.465 ;
        RECT  3.615 0.700 3.690 1.045 ;
        RECT  3.395 0.350 3.615 0.465 ;
        RECT  3.395 0.700 3.615 0.820 ;
        RECT  3.330 0.350 3.395 0.820 ;
        RECT  3.250 0.185 3.330 1.045 ;
        RECT  3.185 0.350 3.250 0.820 ;
        RECT  2.965 0.350 3.185 0.465 ;
        RECT  2.970 0.700 3.185 0.820 ;
        RECT  2.890 0.700 2.970 1.045 ;
        RECT  2.895 0.185 2.965 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0568 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.610 2.345 0.780 ;
        RECT  1.810 0.710 2.275 0.780 ;
        RECT  1.715 0.495 1.810 0.780 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.440 ;
        RECT  3.530 -0.115 3.790 0.115 ;
        RECT  3.410 -0.115 3.530 0.280 ;
        RECT  3.170 -0.115 3.410 0.115 ;
        RECT  3.050 -0.115 3.170 0.280 ;
        RECT  2.810 -0.115 3.050 0.115 ;
        RECT  2.690 -0.115 2.810 0.250 ;
        RECT  1.150 -0.115 2.690 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.760 3.870 1.375 ;
        RECT  3.530 1.145 3.790 1.375 ;
        RECT  3.410 0.890 3.530 1.375 ;
        RECT  3.170 1.145 3.410 1.375 ;
        RECT  3.050 0.890 3.170 1.375 ;
        RECT  2.780 1.145 3.050 1.375 ;
        RECT  2.700 0.990 2.780 1.375 ;
        RECT  2.410 1.145 2.700 1.375 ;
        RECT  2.330 0.990 2.410 1.375 ;
        RECT  2.050 1.145 2.330 1.375 ;
        RECT  1.970 0.920 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.615 0.185 3.690 0.465 ;
        RECT  3.615 0.700 3.690 1.045 ;
        RECT  3.465 0.350 3.615 0.465 ;
        RECT  3.465 0.700 3.615 0.820 ;
        RECT  2.965 0.350 3.115 0.465 ;
        RECT  2.970 0.700 3.115 0.820 ;
        RECT  2.890 0.700 2.970 1.045 ;
        RECT  2.895 0.185 2.965 0.465 ;
        RECT  3.475 0.545 3.815 0.615 ;
        RECT  2.820 0.545 3.100 0.615 ;
        RECT  2.750 0.320 2.820 0.920 ;
        RECT  2.425 0.320 2.750 0.390 ;
        RECT  2.610 0.850 2.750 0.920 ;
        RECT  2.600 0.460 2.670 0.640 ;
        RECT  2.490 0.850 2.610 1.060 ;
        RECT  2.140 0.460 2.600 0.530 ;
        RECT  2.250 0.850 2.490 0.920 ;
        RECT  2.355 0.215 2.425 0.390 ;
        RECT  2.130 0.850 2.250 1.060 ;
        RECT  2.060 0.205 2.140 0.640 ;
        RECT  1.330 0.205 2.060 0.275 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD6BWP

MACRO CKLNQD8BWP
    CLASS CORE ;
    FOREIGN CKLNQD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.3808 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.715 4.130 0.945 ;
        RECT  4.035 0.185 4.105 0.465 ;
        RECT  3.745 0.350 4.035 0.465 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.385 0.350 3.675 0.945 ;
        RECT  3.325 0.185 3.385 0.945 ;
        RECT  3.315 0.185 3.325 0.465 ;
        RECT  2.930 0.715 3.325 0.945 ;
        RECT  3.030 0.350 3.315 0.465 ;
        RECT  2.960 0.185 3.030 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0242 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.475 0.385 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.0568 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.610 2.485 0.770 ;
        RECT  1.810 0.700 2.415 0.770 ;
        RECT  1.715 0.495 1.810 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.440 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.280 ;
        RECT  3.590 -0.115 3.830 0.115 ;
        RECT  3.470 -0.115 3.590 0.280 ;
        RECT  3.230 -0.115 3.470 0.115 ;
        RECT  3.110 -0.115 3.230 0.280 ;
        RECT  2.860 -0.115 3.110 0.115 ;
        RECT  2.740 -0.115 2.860 0.250 ;
        RECT  1.150 -0.115 2.740 0.115 ;
        RECT  1.080 -0.115 1.150 0.295 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.675 4.290 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 1.015 3.950 1.375 ;
        RECT  3.590 1.145 3.830 1.375 ;
        RECT  3.470 1.015 3.590 1.375 ;
        RECT  3.230 1.145 3.470 1.375 ;
        RECT  3.110 1.015 3.230 1.375 ;
        RECT  2.860 1.145 3.110 1.375 ;
        RECT  2.740 1.000 2.860 1.375 ;
        RECT  2.480 1.145 2.740 1.375 ;
        RECT  2.360 1.000 2.480 1.375 ;
        RECT  2.070 1.145 2.360 1.375 ;
        RECT  1.990 0.910 2.070 1.375 ;
        RECT  1.700 1.145 1.990 1.375 ;
        RECT  1.580 0.990 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.020 1.120 1.375 ;
        RECT  0.130 1.145 1.000 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.715 4.130 0.945 ;
        RECT  4.035 0.185 4.105 0.465 ;
        RECT  3.745 0.350 4.035 0.465 ;
        RECT  3.030 0.350 3.255 0.465 ;
        RECT  2.930 0.715 3.255 0.945 ;
        RECT  2.960 0.185 3.030 0.465 ;
        RECT  3.775 0.545 4.140 0.615 ;
        RECT  2.860 0.545 3.225 0.615 ;
        RECT  2.790 0.320 2.860 0.910 ;
        RECT  2.445 0.320 2.790 0.390 ;
        RECT  2.645 0.840 2.790 0.910 ;
        RECT  2.640 0.460 2.710 0.640 ;
        RECT  2.575 0.840 2.645 1.075 ;
        RECT  2.155 0.460 2.640 0.530 ;
        RECT  2.290 0.840 2.575 0.910 ;
        RECT  2.375 0.215 2.445 0.390 ;
        RECT  2.170 0.840 2.290 1.050 ;
        RECT  2.085 0.205 2.155 0.630 ;
        RECT  1.330 0.205 2.085 0.275 ;
        RECT  1.640 0.355 1.890 0.425 ;
        RECT  1.795 0.850 1.865 1.050 ;
        RECT  1.640 0.850 1.795 0.920 ;
        RECT  1.570 0.355 1.640 0.920 ;
        RECT  1.550 0.535 1.570 0.655 ;
        RECT  1.480 0.355 1.500 0.475 ;
        RECT  1.410 0.355 1.480 1.040 ;
        RECT  0.855 0.880 1.410 0.950 ;
        RECT  1.260 0.205 1.330 0.810 ;
        RECT  1.005 0.740 1.260 0.810 ;
        RECT  1.120 0.395 1.190 0.640 ;
        RECT  1.010 0.395 1.120 0.465 ;
        RECT  0.940 0.245 1.010 0.465 ;
        RECT  0.935 0.595 1.005 0.810 ;
        RECT  0.690 0.245 0.940 0.315 ;
        RECT  0.855 0.395 0.870 0.515 ;
        RECT  0.785 0.395 0.855 1.055 ;
        RECT  0.550 0.985 0.785 1.055 ;
        RECT  0.620 0.245 0.690 0.905 ;
        RECT  0.480 0.590 0.550 1.055 ;
        RECT  0.445 0.220 0.525 0.375 ;
        RECT  0.130 0.305 0.445 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD8BWP

MACRO CKMUX2D0BWP
    CLASS CORE ;
    FOREIGN CKMUX2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.045 ;
        RECT  1.275 0.185 1.295 0.305 ;
        RECT  1.275 0.920 1.295 1.045 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.625 ;
        RECT  0.985 0.500 1.015 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 -0.115 1.400 0.115 ;
        RECT  1.080 -0.115 1.160 0.255 ;
        RECT  0.360 -0.115 1.080 0.115 ;
        RECT  0.240 -0.115 0.360 0.285 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.145 1.400 1.375 ;
        RECT  1.060 0.980 1.180 1.375 ;
        RECT  0.330 1.145 1.060 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.195 0.360 1.225 0.765 ;
        RECT  1.155 0.360 1.195 0.910 ;
        RECT  1.125 0.695 1.155 0.910 ;
        RECT  0.740 0.840 1.125 0.910 ;
        RECT  0.915 0.700 0.980 0.770 ;
        RECT  0.915 0.185 0.950 0.305 ;
        RECT  0.845 0.185 0.915 0.770 ;
        RECT  0.760 0.985 0.880 1.075 ;
        RECT  0.560 0.985 0.760 1.055 ;
        RECT  0.670 0.325 0.740 0.910 ;
        RECT  0.520 0.325 0.590 0.810 ;
        RECT  0.490 0.880 0.560 1.055 ;
        RECT  0.465 0.325 0.520 0.400 ;
        RECT  0.460 0.710 0.520 0.810 ;
        RECT  0.125 0.880 0.490 0.950 ;
        RECT  0.105 0.230 0.125 0.350 ;
        RECT  0.105 0.880 0.125 1.040 ;
        RECT  0.035 0.230 0.105 1.040 ;
    END
END CKMUX2D0BWP

MACRO CKMUX2D1BWP
    CLASS CORE ;
    FOREIGN CKMUX2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.045 ;
        RECT  1.275 0.185 1.295 0.465 ;
        RECT  1.275 0.920 1.295 1.045 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0170 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.625 ;
        RECT  0.970 0.500 1.015 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0162 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 -0.115 1.400 0.115 ;
        RECT  1.080 -0.115 1.160 0.255 ;
        RECT  0.360 -0.115 1.080 0.115 ;
        RECT  0.230 -0.115 0.360 0.280 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.145 1.400 1.375 ;
        RECT  1.060 0.980 1.180 1.375 ;
        RECT  0.330 1.145 1.060 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.195 0.520 1.225 0.765 ;
        RECT  1.155 0.520 1.195 0.910 ;
        RECT  1.125 0.695 1.155 0.910 ;
        RECT  0.740 0.840 1.125 0.910 ;
        RECT  0.900 0.700 0.980 0.770 ;
        RECT  0.900 0.185 0.950 0.305 ;
        RECT  0.830 0.185 0.900 0.770 ;
        RECT  0.760 0.985 0.880 1.075 ;
        RECT  0.560 0.985 0.760 1.055 ;
        RECT  0.670 0.325 0.740 0.910 ;
        RECT  0.520 0.325 0.590 0.810 ;
        RECT  0.490 0.880 0.560 1.055 ;
        RECT  0.465 0.325 0.520 0.400 ;
        RECT  0.460 0.710 0.520 0.810 ;
        RECT  0.125 0.880 0.490 0.950 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.880 0.125 1.040 ;
        RECT  0.035 0.210 0.105 1.040 ;
    END
END CKMUX2D1BWP

MACRO CKMUX2D2BWP
    CLASS CORE ;
    FOREIGN CKMUX2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.700 1.330 0.770 ;
        RECT  1.235 0.185 1.305 0.470 ;
        RECT  1.225 0.400 1.235 0.470 ;
        RECT  1.155 0.400 1.225 0.770 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0170 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.990 0.510 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0162 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.440 ;
        RECT  1.130 -0.115 1.410 0.115 ;
        RECT  1.050 -0.115 1.130 0.275 ;
        RECT  0.360 -0.115 1.050 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.980 1.490 1.375 ;
        RECT  0.330 1.145 1.410 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.410 0.540 1.480 0.910 ;
        RECT  1.310 0.540 1.410 0.620 ;
        RECT  0.740 0.840 1.410 0.910 ;
        RECT  0.900 0.700 0.970 0.770 ;
        RECT  0.900 0.185 0.940 0.305 ;
        RECT  0.830 0.185 0.900 0.770 ;
        RECT  0.760 0.985 0.880 1.075 ;
        RECT  0.560 0.985 0.760 1.055 ;
        RECT  0.670 0.325 0.740 0.910 ;
        RECT  0.520 0.325 0.590 0.810 ;
        RECT  0.490 0.880 0.560 1.055 ;
        RECT  0.460 0.325 0.520 0.400 ;
        RECT  0.460 0.710 0.520 0.810 ;
        RECT  0.125 0.880 0.490 0.950 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.880 0.125 1.040 ;
        RECT  0.035 0.210 0.105 1.040 ;
    END
END CKMUX2D2BWP

MACRO CKMUX2D4BWP
    CLASS CORE ;
    FOREIGN CKMUX2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.185 2.145 0.465 ;
        RECT  2.135 0.710 2.145 1.050 ;
        RECT  2.075 0.185 2.135 1.050 ;
        RECT  1.925 0.345 2.075 0.830 ;
        RECT  1.785 0.345 1.925 0.465 ;
        RECT  1.790 0.710 1.925 0.830 ;
        RECT  1.720 0.710 1.790 1.050 ;
        RECT  1.715 0.185 1.785 0.465 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.090 0.495 1.155 0.640 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.370 0.650 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.145 0.495 0.245 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.990 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.990 0.270 ;
        RECT  0.330 -0.115 1.870 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.145 2.380 1.375 ;
        RECT  2.250 0.675 2.330 1.375 ;
        RECT  1.990 1.145 2.250 1.375 ;
        RECT  1.870 0.900 1.990 1.375 ;
        RECT  1.630 1.145 1.870 1.375 ;
        RECT  1.510 1.020 1.630 1.375 ;
        RECT  1.270 1.145 1.510 1.375 ;
        RECT  1.150 1.020 1.270 1.375 ;
        RECT  0.310 1.145 1.150 1.375 ;
        RECT  0.230 0.985 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.345 1.855 0.465 ;
        RECT  1.790 0.710 1.855 0.830 ;
        RECT  1.720 0.710 1.790 1.050 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.650 0.545 1.760 0.615 ;
        RECT  1.580 0.545 1.650 0.950 ;
        RECT  0.665 0.880 1.580 0.950 ;
        RECT  1.440 0.205 1.510 0.800 ;
        RECT  0.820 0.205 1.440 0.275 ;
        RECT  1.330 0.730 1.440 0.800 ;
        RECT  1.010 0.730 1.070 0.800 ;
        RECT  1.010 0.345 1.050 0.415 ;
        RECT  0.940 0.345 1.010 0.800 ;
        RECT  0.930 0.345 0.940 0.620 ;
        RECT  0.890 0.500 0.930 0.620 ;
        RECT  0.820 0.690 0.860 0.810 ;
        RECT  0.750 0.205 0.820 0.810 ;
        RECT  0.595 0.200 0.665 0.995 ;
        RECT  0.415 0.200 0.485 0.990 ;
        RECT  0.125 0.350 0.415 0.420 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.240 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END CKMUX2D4BWP

MACRO CKND0BWP
    CLASS CORE ;
    FOREIGN CKND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0374 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.295 0.385 0.950 ;
        RECT  0.295 0.295 0.315 0.415 ;
        RECT  0.295 0.820 0.315 0.950 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0136 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 -0.115 0.420 0.115 ;
        RECT  0.100 -0.115 0.180 0.415 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.145 0.420 1.375 ;
        RECT  0.100 0.845 0.180 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
END CKND0BWP

MACRO CKND12BWP
    CLASS CORE ;
    FOREIGN CKND12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5829 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.715 2.170 0.945 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.325 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.325 1.715 0.465 ;
        RECT  1.355 0.185 1.425 0.465 ;
        RECT  1.295 0.325 1.355 0.465 ;
        RECT  1.065 0.325 1.295 0.945 ;
        RECT  0.995 0.185 1.065 0.945 ;
        RECT  0.945 0.325 0.995 0.945 ;
        RECT  0.705 0.325 0.945 0.465 ;
        RECT  0.210 0.715 0.945 0.945 ;
        RECT  0.635 0.185 0.705 0.465 ;
        RECT  0.345 0.325 0.635 0.465 ;
        RECT  0.275 0.185 0.345 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.845 0.625 ;
        RECT  0.035 0.200 0.125 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.990 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.990 0.255 ;
        RECT  1.630 -0.115 1.870 0.115 ;
        RECT  1.510 -0.115 1.630 0.255 ;
        RECT  1.270 -0.115 1.510 0.115 ;
        RECT  1.150 -0.115 1.270 0.255 ;
        RECT  0.910 -0.115 1.150 0.115 ;
        RECT  0.790 -0.115 0.910 0.255 ;
        RECT  0.550 -0.115 0.790 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.145 2.380 1.375 ;
        RECT  2.250 0.680 2.330 1.375 ;
        RECT  1.990 1.145 2.250 1.375 ;
        RECT  1.870 1.015 1.990 1.375 ;
        RECT  1.620 1.145 1.870 1.375 ;
        RECT  1.500 1.015 1.620 1.375 ;
        RECT  1.250 1.145 1.500 1.375 ;
        RECT  1.130 1.015 1.250 1.375 ;
        RECT  0.880 1.145 1.130 1.375 ;
        RECT  0.760 1.015 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.715 2.170 0.945 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.325 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.325 1.715 0.465 ;
        RECT  1.365 0.185 1.425 0.465 ;
        RECT  0.705 0.325 0.875 0.465 ;
        RECT  0.210 0.715 0.875 0.945 ;
        RECT  0.635 0.185 0.705 0.465 ;
        RECT  0.345 0.325 0.635 0.465 ;
        RECT  0.275 0.185 0.345 0.465 ;
        RECT  1.415 0.545 2.220 0.615 ;
    END
END CKND12BWP

MACRO CKND16BWP
    CLASS CORE ;
    FOREIGN CKND16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.715 2.870 0.945 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.125 0.305 2.415 0.465 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.765 0.305 2.055 0.465 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.695 0.185 1.715 0.945 ;
        RECT  1.405 0.305 1.695 0.945 ;
        RECT  1.365 0.185 1.405 0.945 ;
        RECT  1.335 0.185 1.365 0.465 ;
        RECT  0.210 0.715 1.365 0.945 ;
        RECT  1.045 0.305 1.335 0.465 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  0.625 0.305 0.975 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4352 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 1.265 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.115 3.080 0.115 ;
        RECT  2.955 -0.115 3.025 0.475 ;
        RECT  2.690 -0.115 2.955 0.115 ;
        RECT  2.570 -0.115 2.690 0.235 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.235 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.235 ;
        RECT  1.610 -0.115 1.850 0.115 ;
        RECT  1.490 -0.115 1.610 0.235 ;
        RECT  1.250 -0.115 1.490 0.115 ;
        RECT  1.130 -0.115 1.250 0.235 ;
        RECT  0.860 -0.115 1.130 0.115 ;
        RECT  0.740 -0.115 0.860 0.235 ;
        RECT  0.445 -0.115 0.740 0.115 ;
        RECT  0.375 -0.115 0.445 0.460 ;
        RECT  0.000 -0.115 0.375 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.675 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 1.015 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.015 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.015 1.970 1.375 ;
        RECT  1.610 1.145 1.850 1.375 ;
        RECT  1.490 1.015 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 1.015 1.250 1.375 ;
        RECT  0.880 1.145 1.130 1.375 ;
        RECT  0.760 1.015 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.715 2.870 0.945 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.125 0.305 2.415 0.465 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.785 0.305 2.055 0.465 ;
        RECT  1.045 0.305 1.295 0.465 ;
        RECT  0.210 0.715 1.295 0.945 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  0.625 0.305 0.975 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        RECT  1.815 0.545 2.805 0.615 ;
    END
END CKND16BWP

MACRO CKND1BWP
    CLASS CORE ;
    FOREIGN CKND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0748 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.215 0.385 1.075 ;
        RECT  0.295 0.215 0.315 0.355 ;
        RECT  0.295 0.815 0.315 1.075 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 -0.115 0.420 0.115 ;
        RECT  0.100 -0.115 0.180 0.355 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.145 0.420 1.375 ;
        RECT  0.100 0.850 0.180 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
END CKND1BWP

MACRO CKND20BWP
    CLASS CORE ;
    FOREIGN CKND20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.715 3.570 0.945 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.305 2.755 0.465 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.135 0.305 2.395 0.465 ;
        RECT  2.105 0.305 2.135 0.945 ;
        RECT  2.035 0.185 2.105 0.945 ;
        RECT  1.785 0.305 2.035 0.945 ;
        RECT  1.745 0.305 1.785 0.465 ;
        RECT  0.210 0.715 1.785 0.945 ;
        RECT  1.675 0.185 1.745 0.465 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.005 0.305 1.315 0.465 ;
        RECT  0.935 0.185 1.005 0.465 ;
        RECT  0.625 0.305 0.935 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.5440 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 1.685 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.115 3.780 0.115 ;
        RECT  3.655 -0.115 3.725 0.465 ;
        RECT  3.390 -0.115 3.655 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.235 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.235 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.235 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.235 ;
        RECT  1.220 -0.115 1.470 0.115 ;
        RECT  1.100 -0.115 1.220 0.235 ;
        RECT  0.840 -0.115 1.100 0.115 ;
        RECT  0.720 -0.115 0.840 0.235 ;
        RECT  0.450 -0.115 0.720 0.115 ;
        RECT  0.370 -0.115 0.450 0.460 ;
        RECT  0.000 -0.115 0.370 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.675 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.015 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.015 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.015 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 1.015 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 1.015 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.015 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.015 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.715 3.570 0.945 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.305 2.755 0.465 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.205 0.305 2.395 0.465 ;
        RECT  1.675 0.185 1.715 0.465 ;
        RECT  0.210 0.715 1.715 0.945 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.005 0.305 1.315 0.465 ;
        RECT  0.935 0.185 1.005 0.465 ;
        RECT  0.625 0.305 0.935 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        RECT  2.235 0.545 3.565 0.615 ;
    END
END CKND20BWP

MACRO CKND24BWP
    CLASS CORE ;
    FOREIGN CKND24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.1536 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.715 4.410 0.945 ;
        RECT  4.315 0.185 4.385 0.465 ;
        RECT  3.965 0.305 4.315 0.465 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.545 0.305 3.895 0.465 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.305 2.755 0.465 ;
        RECT  2.415 0.185 2.465 0.465 ;
        RECT  2.395 0.185 2.415 0.945 ;
        RECT  2.105 0.305 2.395 0.945 ;
        RECT  2.065 0.185 2.105 0.945 ;
        RECT  2.035 0.185 2.065 0.465 ;
        RECT  0.210 0.715 2.065 0.945 ;
        RECT  1.745 0.305 2.035 0.465 ;
        RECT  1.675 0.185 1.745 0.465 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.025 0.305 1.315 0.465 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.665 0.305 0.955 0.465 ;
        RECT  0.595 0.185 0.665 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6528 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 1.965 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.475 ;
        RECT  4.200 -0.115 4.490 0.115 ;
        RECT  4.080 -0.115 4.200 0.235 ;
        RECT  3.780 -0.115 4.080 0.115 ;
        RECT  3.660 -0.115 3.780 0.235 ;
        RECT  3.390 -0.115 3.660 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.235 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.235 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.235 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.235 ;
        RECT  1.230 -0.115 1.470 0.115 ;
        RECT  1.110 -0.115 1.230 0.235 ;
        RECT  0.870 -0.115 1.110 0.115 ;
        RECT  0.750 -0.115 0.870 0.235 ;
        RECT  0.000 -0.115 0.750 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.675 4.570 1.375 ;
        RECT  4.200 1.145 4.490 1.375 ;
        RECT  4.080 1.015 4.200 1.375 ;
        RECT  3.780 1.145 4.080 1.375 ;
        RECT  3.660 1.015 3.780 1.375 ;
        RECT  3.390 1.145 3.660 1.375 ;
        RECT  3.270 1.015 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.015 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.015 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 1.015 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 1.015 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.015 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.015 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.715 4.410 0.945 ;
        RECT  4.315 0.185 4.385 0.465 ;
        RECT  3.965 0.305 4.315 0.465 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.545 0.305 3.895 0.465 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.485 0.305 2.755 0.465 ;
        RECT  1.745 0.305 1.995 0.465 ;
        RECT  0.210 0.715 1.995 0.945 ;
        RECT  1.675 0.185 1.745 0.465 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.025 0.305 1.315 0.465 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.665 0.305 0.955 0.465 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  2.515 0.545 4.355 0.615 ;
    END
END CKND24BWP

MACRO CKND2BWP
    CLASS CORE ;
    FOREIGN CKND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.355 0.385 0.905 ;
        RECT  0.310 0.215 0.320 1.045 ;
        RECT  0.240 0.215 0.310 0.425 ;
        RECT  0.240 0.765 0.310 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.300 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 0.560 1.375 ;
        RECT  0.430 0.980 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END CKND2BWP

MACRO CKND2D0BWP
    CLASS CORE ;
    FOREIGN CKND2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0418 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 0.915 ;
        RECT  0.390 0.185 0.455 0.265 ;
        RECT  0.310 0.845 0.455 0.915 ;
        RECT  0.230 0.845 0.310 1.050 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0124 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.560 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.145 0.560 1.375 ;
        RECT  0.410 0.985 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.985 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END CKND2D0BWP

MACRO CKND2D1BWP
    CLASS CORE ;
    FOREIGN CKND2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0837 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.215 0.525 0.905 ;
        RECT  0.415 0.215 0.455 0.345 ;
        RECT  0.330 0.835 0.455 0.905 ;
        RECT  0.210 0.835 0.330 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.560 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.145 0.560 1.375 ;
        RECT  0.410 0.980 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END CKND2D1BWP

MACRO CKND2D2BWP
    CLASS CORE ;
    FOREIGN CKND2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1302 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.745 0.750 1.045 ;
        RECT  0.385 0.745 0.670 0.820 ;
        RECT  0.330 0.345 0.385 0.820 ;
        RECT  0.310 0.345 0.330 1.045 ;
        RECT  0.230 0.345 0.310 0.415 ;
        RECT  0.250 0.745 0.310 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0496 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.695 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0496 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.980 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.750 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.940 0.560 1.375 ;
        RECT  0.150 1.145 0.440 1.375 ;
        RECT  0.070 0.920 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.205 0.930 0.345 ;
        RECT  0.150 0.205 0.850 0.275 ;
        RECT  0.070 0.205 0.150 0.345 ;
    END
END CKND2D2BWP

MACRO CKND2D3BWP
    CLASS CORE ;
    FOREIGN CKND2D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2077 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.725 1.030 1.050 ;
        RECT  0.670 0.725 0.950 0.815 ;
        RECT  0.590 0.725 0.670 1.050 ;
        RECT  0.525 0.725 0.590 0.815 ;
        RECT  0.455 0.345 0.525 0.815 ;
        RECT  0.130 0.345 0.455 0.415 ;
        RECT  0.310 0.725 0.455 0.815 ;
        RECT  0.230 0.725 0.310 1.050 ;
        RECT  0.050 0.215 0.130 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0744 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.065 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0744 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.440 ;
        RECT  0.850 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.850 0.265 ;
        RECT  0.000 -0.115 0.770 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.735 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.940 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.940 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.930 0.205 1.050 0.415 ;
        RECT  0.665 0.345 0.930 0.415 ;
        RECT  0.595 0.205 0.665 0.415 ;
        RECT  0.210 0.205 0.595 0.275 ;
    END
END CKND2D3BWP

MACRO CKND2D4BWP
    CLASS CORE ;
    FOREIGN CKND2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2604 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.775 1.445 1.075 ;
        RECT  1.085 0.775 1.375 0.935 ;
        RECT  1.015 0.775 1.085 1.075 ;
        RECT  0.665 0.775 1.015 0.935 ;
        RECT  0.595 0.335 0.690 0.415 ;
        RECT  0.595 0.775 0.665 1.075 ;
        RECT  0.385 0.335 0.595 0.935 ;
        RECT  0.210 0.335 0.385 0.415 ;
        RECT  0.305 0.775 0.385 0.935 ;
        RECT  0.235 0.775 0.305 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0992 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.505 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0992 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.250 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 1.680 0.115 ;
        RECT  1.360 -0.115 1.460 0.270 ;
        RECT  1.100 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.100 0.270 ;
        RECT  0.000 -0.115 1.000 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.790 1.630 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 1.005 1.290 1.375 ;
        RECT  0.900 1.145 1.170 1.375 ;
        RECT  0.780 1.025 0.900 1.375 ;
        RECT  0.510 1.145 0.780 1.375 ;
        RECT  0.390 1.005 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.775 1.445 1.075 ;
        RECT  1.085 0.775 1.375 0.935 ;
        RECT  1.015 0.775 1.085 1.075 ;
        RECT  0.665 0.775 1.015 0.935 ;
        RECT  0.665 0.335 0.690 0.415 ;
        RECT  0.210 0.335 0.315 0.415 ;
        RECT  0.305 0.775 0.315 0.935 ;
        RECT  0.235 0.775 0.305 1.075 ;
        RECT  1.555 0.230 1.625 0.415 ;
        RECT  0.880 0.345 1.555 0.415 ;
        RECT  0.800 0.195 0.880 0.415 ;
        RECT  0.125 0.195 0.800 0.265 ;
        RECT  0.055 0.195 0.125 0.375 ;
    END
END CKND2D4BWP

MACRO CKND2D8BWP
    CLASS CORE ;
    FOREIGN CKND2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5208 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.780 2.845 1.075 ;
        RECT  2.485 0.780 2.775 0.935 ;
        RECT  2.415 0.780 2.485 1.075 ;
        RECT  2.125 0.780 2.415 0.935 ;
        RECT  2.055 0.780 2.125 1.075 ;
        RECT  1.765 0.780 2.055 0.935 ;
        RECT  1.695 0.780 1.765 1.075 ;
        RECT  1.385 0.780 1.695 0.935 ;
        RECT  1.295 0.335 1.410 0.425 ;
        RECT  1.315 0.780 1.385 1.075 ;
        RECT  1.295 0.780 1.315 0.935 ;
        RECT  1.085 0.335 1.295 0.935 ;
        RECT  0.210 0.335 1.085 0.425 ;
        RECT  1.025 0.780 1.085 0.935 ;
        RECT  0.955 0.780 1.025 1.075 ;
        RECT  0.665 0.780 0.955 0.935 ;
        RECT  0.595 0.780 0.665 1.075 ;
        RECT  0.305 0.780 0.595 0.935 ;
        RECT  0.235 0.780 0.305 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1984 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.635 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1984 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.955 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 -0.115 3.080 0.115 ;
        RECT  2.760 -0.115 2.860 0.270 ;
        RECT  2.500 -0.115 2.760 0.115 ;
        RECT  2.400 -0.115 2.500 0.270 ;
        RECT  2.140 -0.115 2.400 0.115 ;
        RECT  2.040 -0.115 2.140 0.270 ;
        RECT  1.780 -0.115 2.040 0.115 ;
        RECT  1.680 -0.115 1.780 0.270 ;
        RECT  0.000 -0.115 1.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.780 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.005 1.970 1.375 ;
        RECT  1.600 1.145 1.850 1.375 ;
        RECT  1.480 1.025 1.600 1.375 ;
        RECT  1.230 1.145 1.480 1.375 ;
        RECT  1.110 1.005 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.005 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 1.005 0.510 1.375 ;
        RECT  0.125 1.145 0.390 1.375 ;
        RECT  0.055 0.780 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.775 0.780 2.845 1.075 ;
        RECT  2.485 0.780 2.775 0.935 ;
        RECT  2.415 0.780 2.485 1.075 ;
        RECT  2.125 0.780 2.415 0.935 ;
        RECT  2.055 0.780 2.125 1.075 ;
        RECT  1.765 0.780 2.055 0.935 ;
        RECT  1.695 0.780 1.765 1.075 ;
        RECT  1.385 0.780 1.695 0.935 ;
        RECT  1.365 0.335 1.410 0.425 ;
        RECT  1.365 0.780 1.385 1.075 ;
        RECT  0.210 0.335 1.015 0.425 ;
        RECT  0.955 0.780 1.015 1.075 ;
        RECT  0.665 0.780 0.955 0.935 ;
        RECT  0.595 0.780 0.665 1.075 ;
        RECT  0.305 0.780 0.595 0.935 ;
        RECT  0.235 0.780 0.305 1.075 ;
        RECT  2.955 0.235 3.025 0.415 ;
        RECT  1.580 0.345 2.955 0.415 ;
        RECT  1.500 0.195 1.580 0.415 ;
        RECT  0.125 0.195 1.500 0.265 ;
        RECT  0.055 0.195 0.125 0.375 ;
    END
END CKND2D8BWP

MACRO CKND3BWP
    CLASS CORE ;
    FOREIGN CKND3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1972 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.215 0.765 0.415 ;
        RECT  0.695 0.700 0.765 1.050 ;
        RECT  0.595 0.295 0.695 0.415 ;
        RECT  0.595 0.700 0.695 0.820 ;
        RECT  0.385 0.295 0.595 0.820 ;
        RECT  0.325 0.295 0.385 0.415 ;
        RECT  0.325 0.700 0.385 0.820 ;
        RECT  0.255 0.215 0.325 0.415 ;
        RECT  0.255 0.700 0.325 1.050 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0816 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.580 0.225 ;
        RECT  0.150 -0.115 0.460 0.115 ;
        RECT  0.070 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.890 0.580 1.375 ;
        RECT  0.150 1.145 0.460 1.375 ;
        RECT  0.070 0.750 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.695 0.215 0.765 0.415 ;
        RECT  0.695 0.700 0.765 1.050 ;
        RECT  0.665 0.295 0.695 0.415 ;
        RECT  0.665 0.700 0.695 0.820 ;
        RECT  0.255 0.215 0.315 0.415 ;
        RECT  0.255 0.700 0.315 1.050 ;
    END
END CKND3BWP

MACRO CKND4BWP
    CLASS CORE ;
    FOREIGN CKND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1904 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.215 0.745 0.415 ;
        RECT  0.675 0.700 0.745 1.045 ;
        RECT  0.595 0.305 0.675 0.415 ;
        RECT  0.595 0.700 0.675 0.820 ;
        RECT  0.385 0.305 0.595 0.820 ;
        RECT  0.325 0.305 0.385 0.415 ;
        RECT  0.325 0.700 0.385 0.820 ;
        RECT  0.255 0.215 0.325 0.415 ;
        RECT  0.255 0.700 0.325 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1088 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.530 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.440 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.235 ;
        RECT  0.150 -0.115 0.440 0.115 ;
        RECT  0.070 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.675 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.150 1.145 0.440 1.375 ;
        RECT  0.070 0.750 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.675 0.215 0.745 0.415 ;
        RECT  0.675 0.700 0.745 1.045 ;
        RECT  0.665 0.305 0.675 0.415 ;
        RECT  0.665 0.700 0.675 0.820 ;
        RECT  0.255 0.215 0.315 0.415 ;
        RECT  0.255 0.700 0.315 1.045 ;
    END
END CKND4BWP

MACRO CKND6BWP
    CLASS CORE ;
    FOREIGN CKND6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2856 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.215 1.025 0.465 ;
        RECT  0.955 0.700 1.025 1.045 ;
        RECT  0.735 0.345 0.955 0.465 ;
        RECT  0.735 0.700 0.955 0.820 ;
        RECT  0.665 0.345 0.735 0.820 ;
        RECT  0.595 0.215 0.665 1.045 ;
        RECT  0.525 0.345 0.595 0.820 ;
        RECT  0.305 0.345 0.525 0.465 ;
        RECT  0.305 0.700 0.525 0.820 ;
        RECT  0.235 0.215 0.305 0.465 ;
        RECT  0.235 0.700 0.305 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1632 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.445 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.410 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.270 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.270 ;
        RECT  0.130 -0.115 0.390 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.750 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.890 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.890 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.760 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.215 1.025 0.465 ;
        RECT  0.955 0.700 1.025 1.045 ;
        RECT  0.805 0.345 0.955 0.465 ;
        RECT  0.805 0.700 0.955 0.820 ;
        RECT  0.305 0.345 0.455 0.465 ;
        RECT  0.305 0.700 0.455 0.820 ;
        RECT  0.235 0.215 0.305 0.465 ;
        RECT  0.235 0.700 0.305 1.045 ;
        RECT  0.815 0.545 1.155 0.615 ;
    END
END CKND6BWP

MACRO CKND8BWP
    CLASS CORE ;
    FOREIGN CKND8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3928 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.730 1.470 0.960 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.295 0.345 1.375 0.465 ;
        RECT  1.085 0.345 1.295 0.960 ;
        RECT  1.015 0.185 1.085 0.960 ;
        RECT  0.945 0.345 1.015 0.960 ;
        RECT  0.725 0.345 0.945 0.465 ;
        RECT  0.210 0.730 0.945 0.960 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.365 0.345 0.655 0.465 ;
        RECT  0.295 0.185 0.365 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2176 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 0.845 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.625 -0.115 1.680 0.115 ;
        RECT  1.555 -0.115 1.625 0.465 ;
        RECT  1.290 -0.115 1.555 0.115 ;
        RECT  1.170 -0.115 1.290 0.275 ;
        RECT  0.930 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.930 0.275 ;
        RECT  0.570 -0.115 0.810 0.115 ;
        RECT  0.450 -0.115 0.570 0.275 ;
        RECT  0.000 -0.115 0.450 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.675 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 1.030 1.280 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.780 1.030 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 1.030 0.520 1.375 ;
        RECT  0.130 1.145 0.400 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.730 1.470 0.960 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.365 0.345 1.375 0.465 ;
        RECT  0.725 0.345 0.875 0.465 ;
        RECT  0.210 0.730 0.875 0.960 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.365 0.345 0.655 0.465 ;
        RECT  0.295 0.185 0.365 0.465 ;
    END
END CKND8BWP

MACRO CKXOR2D0BWP
    CLASS CORE ;
    FOREIGN CKXOR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0437 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.215 1.365 1.070 ;
        RECT  1.275 0.215 1.295 0.360 ;
        RECT  1.230 0.990 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.085 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.165 -0.115 1.400 0.115 ;
        RECT  1.095 -0.115 1.165 0.360 ;
        RECT  0.260 -0.115 1.095 0.115 ;
        RECT  0.260 0.350 0.335 0.420 ;
        RECT  0.190 -0.115 0.260 0.420 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 1.400 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.640 1.225 0.905 ;
        RECT  1.145 0.835 1.155 0.905 ;
        RECT  1.075 0.835 1.145 1.050 ;
        RECT  0.775 0.980 1.075 1.050 ;
        RECT  0.915 0.265 1.010 0.335 ;
        RECT  0.915 0.840 0.970 0.910 ;
        RECT  0.845 0.205 0.915 0.910 ;
        RECT  0.470 0.205 0.845 0.275 ;
        RECT  0.705 0.355 0.775 1.050 ;
        RECT  0.630 0.710 0.705 0.790 ;
        RECT  0.550 0.870 0.620 1.070 ;
        RECT  0.125 0.870 0.550 0.940 ;
        RECT  0.475 0.350 0.545 0.800 ;
        RECT  0.340 0.195 0.470 0.275 ;
        RECT  0.105 0.870 0.125 1.020 ;
        RECT  0.105 0.295 0.120 0.415 ;
        RECT  0.035 0.295 0.105 1.020 ;
    END
END CKXOR2D0BWP

MACRO CKXOR2D1BWP
    CLASS CORE ;
    FOREIGN CKXOR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0874 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.070 ;
        RECT  1.275 0.185 1.295 0.445 ;
        RECT  1.230 0.990 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.970 0.495 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0310 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 -0.115 1.400 0.115 ;
        RECT  1.080 -0.115 1.160 0.410 ;
        RECT  0.260 -0.115 1.080 0.115 ;
        RECT  0.260 0.350 0.335 0.420 ;
        RECT  0.190 -0.115 0.260 0.420 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 1.400 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.520 1.225 0.915 ;
        RECT  1.145 0.845 1.155 0.915 ;
        RECT  1.075 0.845 1.145 1.050 ;
        RECT  0.760 0.980 1.075 1.050 ;
        RECT  0.900 0.330 0.980 0.410 ;
        RECT  0.900 0.840 0.970 0.910 ;
        RECT  0.830 0.205 0.900 0.910 ;
        RECT  0.460 0.205 0.830 0.275 ;
        RECT  0.690 0.355 0.760 1.050 ;
        RECT  0.630 0.715 0.690 0.795 ;
        RECT  0.550 0.870 0.620 1.060 ;
        RECT  0.125 0.870 0.550 0.940 ;
        RECT  0.475 0.350 0.545 0.800 ;
        RECT  0.435 0.350 0.475 0.470 ;
        RECT  0.340 0.195 0.460 0.275 ;
        RECT  0.105 0.870 0.125 1.020 ;
        RECT  0.105 0.295 0.120 0.415 ;
        RECT  0.035 0.295 0.105 1.020 ;
    END
END CKXOR2D1BWP

MACRO CKXOR2D2BWP
    CLASS CORE ;
    FOREIGN CKXOR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.920 ;
        RECT  1.330 0.355 1.435 0.425 ;
        RECT  1.210 0.850 1.435 0.920 ;
        RECT  1.210 0.215 1.330 0.425 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.990 0.520 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0462 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.285 ;
        RECT  1.130 -0.115 1.410 0.115 ;
        RECT  1.050 -0.115 1.130 0.275 ;
        RECT  0.260 -0.115 1.050 0.115 ;
        RECT  0.260 0.355 0.335 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.990 1.500 1.375 ;
        RECT  1.150 1.145 1.400 1.375 ;
        RECT  1.030 1.010 1.150 1.375 ;
        RECT  0.330 1.145 1.030 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.220 0.520 1.300 0.780 ;
        RECT  1.130 0.710 1.220 0.780 ;
        RECT  1.060 0.710 1.130 0.930 ;
        RECT  0.765 0.860 1.060 0.930 ;
        RECT  0.920 0.720 0.970 0.790 ;
        RECT  0.920 0.195 0.940 0.325 ;
        RECT  0.850 0.195 0.920 0.790 ;
        RECT  0.460 0.195 0.850 0.265 ;
        RECT  0.695 0.335 0.765 0.930 ;
        RECT  0.590 0.715 0.695 0.795 ;
        RECT  0.500 0.880 0.570 1.070 ;
        RECT  0.435 0.350 0.505 0.810 ;
        RECT  0.125 0.880 0.500 0.950 ;
        RECT  0.340 0.195 0.460 0.275 ;
        RECT  0.105 0.880 0.125 1.020 ;
        RECT  0.105 0.295 0.120 0.415 ;
        RECT  0.035 0.295 0.105 1.020 ;
    END
END CKXOR2D2BWP

MACRO CKXOR2D4BWP
    CLASS CORE ;
    FOREIGN CKXOR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.195 2.705 0.475 ;
        RECT  2.695 0.700 2.705 1.055 ;
        RECT  2.635 0.195 2.695 1.055 ;
        RECT  2.485 0.355 2.635 0.820 ;
        RECT  2.345 0.355 2.485 0.475 ;
        RECT  2.345 0.700 2.485 0.820 ;
        RECT  2.275 0.195 2.345 0.475 ;
        RECT  2.275 0.700 2.345 1.055 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.065 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.475 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.275 ;
        RECT  0.670 -0.115 2.430 0.115 ;
        RECT  0.590 -0.115 0.670 0.380 ;
        RECT  0.330 -0.115 0.590 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.675 2.890 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 0.890 2.550 1.375 ;
        RECT  0.310 1.145 2.430 1.375 ;
        RECT  0.230 0.985 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.475 ;
        RECT  2.345 0.700 2.415 0.820 ;
        RECT  2.275 0.195 2.345 0.475 ;
        RECT  2.275 0.700 2.345 1.055 ;
        RECT  2.205 0.545 2.385 0.615 ;
        RECT  2.135 0.210 2.205 1.050 ;
        RECT  1.960 0.210 2.135 0.280 ;
        RECT  1.690 0.980 2.135 1.050 ;
        RECT  1.855 0.350 1.990 0.420 ;
        RECT  1.855 0.840 1.990 0.910 ;
        RECT  1.890 0.195 1.960 0.280 ;
        RECT  1.430 0.195 1.890 0.265 ;
        RECT  1.785 0.350 1.855 0.910 ;
        RECT  1.640 0.335 1.710 0.860 ;
        RECT  1.510 0.335 1.640 0.405 ;
        RECT  1.605 0.790 1.640 0.860 ;
        RECT  1.535 0.790 1.605 1.060 ;
        RECT  1.400 0.500 1.570 0.570 ;
        RECT  0.490 0.990 1.535 1.060 ;
        RECT  1.350 0.195 1.430 0.405 ;
        RECT  1.350 0.710 1.430 0.910 ;
        RECT  1.330 0.500 1.400 0.630 ;
        RECT  1.010 0.335 1.350 0.405 ;
        RECT  1.010 0.710 1.350 0.780 ;
        RECT  1.080 0.560 1.330 0.630 ;
        RECT  0.870 0.850 1.270 0.920 ;
        RECT  0.870 0.195 1.250 0.265 ;
        RECT  0.940 0.335 1.010 0.780 ;
        RECT  0.800 0.195 0.870 0.920 ;
        RECT  0.780 0.195 0.800 0.340 ;
        RECT  0.490 0.520 0.730 0.640 ;
        RECT  0.410 0.185 0.490 1.060 ;
        RECT  0.130 0.330 0.410 0.405 ;
        RECT  0.130 0.845 0.410 0.915 ;
        RECT  0.050 0.240 0.130 0.405 ;
        RECT  0.050 0.845 0.130 0.985 ;
    END
END CKXOR2D4BWP

MACRO CMPE42D1BWP
    CLASS CORE ;
    FOREIGN CMPE42D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.860 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.755 0.185 6.825 1.045 ;
        RECT  6.735 0.185 6.755 0.465 ;
        RECT  6.740 0.735 6.755 1.045 ;
        END
    END S
    PIN D
        ANTENNAGATEAREA 0.0476 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.355 4.725 0.640 ;
        RECT  4.530 0.520 4.655 0.640 ;
        END
    END D
    PIN COX
        ANTENNADIFFAREA 0.0814 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.545 0.350 3.605 0.780 ;
        RECT  3.535 0.185 3.545 0.780 ;
        RECT  3.475 0.185 3.535 0.470 ;
        RECT  3.450 0.710 3.535 0.780 ;
        END
    END COX
    PIN CO
        ANTENNADIFFAREA 0.0814 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.405 0.680 6.450 0.780 ;
        RECT  6.405 0.185 6.425 0.465 ;
        RECT  6.355 0.185 6.405 0.780 ;
        RECT  6.335 0.395 6.355 0.780 ;
        END
    END CO
    PIN CIX
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.175 0.355 6.265 0.640 ;
        RECT  6.100 0.520 6.175 0.640 ;
        END
    END CIX
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.355 3.330 0.640 ;
        RECT  3.220 0.520 3.255 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.975 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.620 -0.115 6.860 0.115 ;
        RECT  6.540 -0.115 6.620 0.440 ;
        RECT  3.750 -0.115 6.540 0.115 ;
        RECT  3.630 -0.115 3.750 0.260 ;
        RECT  0.140 -0.115 3.630 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.640 1.145 6.860 1.375 ;
        RECT  6.520 1.005 6.640 1.375 ;
        RECT  4.690 1.145 6.520 1.375 ;
        RECT  4.570 1.030 4.690 1.375 ;
        RECT  0.890 1.145 4.570 1.375 ;
        RECT  0.770 1.000 0.890 1.375 ;
        RECT  0.500 1.145 0.770 1.375 ;
        RECT  0.420 0.860 0.500 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.660 0.520 6.685 0.640 ;
        RECT  6.590 0.520 6.660 0.920 ;
        RECT  5.630 0.850 6.590 0.920 ;
        RECT  5.250 0.990 6.340 1.060 ;
        RECT  6.030 0.200 6.270 0.270 ;
        RECT  6.030 0.710 6.230 0.780 ;
        RECT  5.960 0.200 6.030 0.780 ;
        RECT  5.490 0.200 5.960 0.280 ;
        RECT  5.890 0.520 5.960 0.640 ;
        RECT  5.820 0.370 5.890 0.440 ;
        RECT  5.750 0.370 5.820 0.765 ;
        RECT  5.700 0.695 5.750 0.765 ;
        RECT  5.630 0.350 5.670 0.470 ;
        RECT  5.560 0.350 5.630 0.920 ;
        RECT  5.490 0.850 5.560 0.920 ;
        RECT  5.420 0.200 5.490 0.630 ;
        RECT  5.390 0.560 5.420 0.630 ;
        RECT  5.320 0.560 5.390 0.890 ;
        RECT  5.250 0.210 5.295 0.470 ;
        RECT  5.225 0.210 5.250 1.060 ;
        RECT  5.180 0.395 5.225 1.060 ;
        RECT  5.140 0.930 5.180 1.060 ;
        RECT  5.040 0.360 5.110 0.850 ;
        RECT  5.025 0.780 5.040 0.850 ;
        RECT  4.955 0.780 5.025 1.035 ;
        RECT  4.900 0.185 5.020 0.275 ;
        RECT  4.885 0.520 4.970 0.640 ;
        RECT  4.490 0.890 4.955 0.960 ;
        RECT  4.090 0.205 4.900 0.275 ;
        RECT  4.880 0.345 4.885 0.640 ;
        RECT  4.810 0.345 4.880 0.810 ;
        RECT  4.750 0.740 4.810 0.810 ;
        RECT  4.460 0.370 4.520 0.440 ;
        RECT  4.460 0.745 4.490 1.035 ;
        RECT  4.410 0.370 4.460 1.035 ;
        RECT  4.390 0.370 4.410 0.815 ;
        RECT  4.320 0.540 4.390 0.610 ;
        RECT  4.250 0.345 4.320 0.460 ;
        RECT  4.260 0.690 4.300 0.960 ;
        RECT  4.250 0.690 4.260 1.050 ;
        RECT  4.190 0.345 4.250 1.050 ;
        RECT  4.180 0.345 4.190 0.770 ;
        RECT  3.745 0.980 4.190 1.050 ;
        RECT  4.090 0.810 4.120 0.910 ;
        RECT  4.020 0.205 4.090 0.910 ;
        RECT  3.905 0.365 3.950 0.905 ;
        RECT  3.880 0.185 3.905 0.905 ;
        RECT  3.835 0.185 3.880 0.445 ;
        RECT  3.830 0.835 3.880 0.905 ;
        RECT  3.745 0.520 3.810 0.640 ;
        RECT  3.675 0.520 3.745 1.050 ;
        RECT  2.755 0.850 3.675 0.920 ;
        RECT  2.330 0.990 3.460 1.060 ;
        RECT  3.150 0.210 3.390 0.280 ;
        RECT  3.150 0.710 3.350 0.780 ;
        RECT  3.080 0.210 3.150 0.780 ;
        RECT  2.605 0.210 3.080 0.280 ;
        RECT  3.000 0.520 3.080 0.640 ;
        RECT  2.930 0.360 3.010 0.430 ;
        RECT  2.860 0.360 2.930 0.780 ;
        RECT  2.755 0.350 2.780 0.470 ;
        RECT  2.685 0.350 2.755 0.920 ;
        RECT  2.590 0.850 2.685 0.920 ;
        RECT  2.535 0.210 2.605 0.630 ;
        RECT  2.505 0.560 2.535 0.630 ;
        RECT  2.435 0.560 2.505 0.890 ;
        RECT  2.330 0.195 2.395 0.495 ;
        RECT  2.325 0.195 2.330 1.060 ;
        RECT  2.260 0.425 2.325 1.060 ;
        RECT  2.120 0.210 2.190 1.000 ;
        RECT  1.600 0.210 2.120 0.280 ;
        RECT  2.050 0.930 2.120 1.000 ;
        RECT  2.010 0.520 2.050 0.640 ;
        RECT  2.000 0.355 2.010 0.640 ;
        RECT  1.965 0.355 2.000 0.805 ;
        RECT  1.930 0.355 1.965 1.035 ;
        RECT  1.880 0.355 1.930 0.425 ;
        RECT  1.895 0.735 1.930 1.035 ;
        RECT  1.775 0.520 1.860 0.640 ;
        RECT  1.705 0.520 1.775 1.050 ;
        RECT  1.230 0.980 1.705 1.050 ;
        RECT  1.525 0.210 1.600 0.910 ;
        RECT  1.515 0.520 1.525 0.910 ;
        RECT  1.450 0.520 1.515 0.640 ;
        RECT  1.380 0.210 1.420 0.330 ;
        RECT  1.380 0.740 1.405 0.860 ;
        RECT  1.310 0.210 1.380 0.860 ;
        RECT  0.480 0.210 1.310 0.280 ;
        RECT  1.150 0.350 1.230 1.050 ;
        RECT  0.790 0.350 1.070 0.420 ;
        RECT  0.975 0.845 1.045 1.035 ;
        RECT  0.790 0.845 0.975 0.920 ;
        RECT  0.720 0.350 0.790 0.920 ;
        RECT  0.590 0.350 0.720 0.420 ;
        RECT  0.685 0.765 0.720 0.920 ;
        RECT  0.615 0.765 0.685 1.035 ;
        RECT  0.480 0.520 0.635 0.640 ;
        RECT  0.410 0.210 0.480 0.790 ;
        RECT  0.305 0.395 0.410 0.465 ;
        RECT  0.305 0.720 0.410 0.790 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.720 0.305 1.035 ;
    END
END CMPE42D1BWP

MACRO CMPE42D2BWP
    CLASS CORE ;
    FOREIGN CMPE42D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.825 0.405 6.875 0.810 ;
        RECT  6.805 0.185 6.825 0.810 ;
        RECT  6.755 0.185 6.805 0.485 ;
        RECT  6.755 0.690 6.805 0.810 ;
        END
    END S
    PIN D
        ANTENNAGATEAREA 0.0476 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.355 4.865 0.640 ;
        RECT  4.750 0.520 4.795 0.640 ;
        END
    END D
    PIN COX
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.185 3.745 0.770 ;
        END
    END COX
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.185 0.355 7.245 0.905 ;
        RECT  7.175 0.185 7.185 1.045 ;
        RECT  7.115 0.185 7.175 0.465 ;
        RECT  7.115 0.785 7.175 1.045 ;
        END
    END CO
    PIN CIX
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.310 0.355 6.405 0.640 ;
        END
    END CIX
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.355 3.330 0.640 ;
        RECT  3.210 0.520 3.255 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.975 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.365 -0.115 7.420 0.115 ;
        RECT  7.295 -0.115 7.365 0.300 ;
        RECT  7.030 -0.115 7.295 0.115 ;
        RECT  6.910 -0.115 7.030 0.245 ;
        RECT  6.645 -0.115 6.910 0.115 ;
        RECT  6.575 -0.115 6.645 0.440 ;
        RECT  3.930 -0.115 6.575 0.115 ;
        RECT  3.850 -0.115 3.930 0.445 ;
        RECT  3.545 -0.115 3.850 0.115 ;
        RECT  3.475 -0.115 3.545 0.465 ;
        RECT  0.140 -0.115 3.475 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.365 1.145 7.420 1.375 ;
        RECT  7.295 0.960 7.365 1.375 ;
        RECT  7.030 1.145 7.295 1.375 ;
        RECT  6.910 1.020 7.030 1.375 ;
        RECT  4.900 1.145 6.910 1.375 ;
        RECT  4.780 1.025 4.900 1.375 ;
        RECT  0.890 1.145 4.780 1.375 ;
        RECT  0.770 0.990 0.890 1.375 ;
        RECT  0.500 1.145 0.770 1.375 ;
        RECT  0.420 0.860 0.500 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.025 0.545 7.100 0.615 ;
        RECT  6.955 0.545 7.025 0.950 ;
        RECT  6.840 0.880 6.955 0.950 ;
        RECT  6.770 0.880 6.840 1.060 ;
        RECT  5.470 0.990 6.770 1.060 ;
        RECT  6.605 0.520 6.675 0.920 ;
        RECT  5.865 0.850 6.605 0.920 ;
        RECT  6.240 0.210 6.490 0.280 ;
        RECT  6.240 0.710 6.490 0.780 ;
        RECT  6.170 0.210 6.240 0.780 ;
        RECT  5.725 0.210 6.170 0.280 ;
        RECT  6.125 0.520 6.170 0.640 ;
        RECT  6.055 0.350 6.100 0.450 ;
        RECT  5.985 0.350 6.055 0.765 ;
        RECT  5.935 0.695 5.985 0.765 ;
        RECT  5.865 0.350 5.900 0.470 ;
        RECT  5.795 0.350 5.865 0.920 ;
        RECT  5.710 0.845 5.795 0.920 ;
        RECT  5.655 0.210 5.725 0.630 ;
        RECT  5.610 0.560 5.655 0.630 ;
        RECT  5.540 0.560 5.610 0.910 ;
        RECT  5.470 0.200 5.495 0.460 ;
        RECT  5.400 0.200 5.470 1.060 ;
        RECT  5.330 0.990 5.400 1.060 ;
        RECT  5.260 0.385 5.330 0.850 ;
        RECT  5.190 0.385 5.260 0.455 ;
        RECT  5.245 0.780 5.260 0.850 ;
        RECT  5.175 0.780 5.245 1.035 ;
        RECT  5.120 0.185 5.240 0.275 ;
        RECT  5.110 0.530 5.190 0.650 ;
        RECT  4.680 0.885 5.175 0.955 ;
        RECT  4.300 0.205 5.120 0.275 ;
        RECT  5.100 0.345 5.110 0.650 ;
        RECT  5.030 0.345 5.100 0.790 ;
        RECT  4.970 0.720 5.030 0.790 ;
        RECT  4.680 0.355 4.710 0.425 ;
        RECT  4.610 0.355 4.680 1.035 ;
        RECT  4.590 0.355 4.610 0.640 ;
        RECT  4.550 0.520 4.590 0.640 ;
        RECT  4.470 0.345 4.505 0.465 ;
        RECT  4.470 0.700 4.500 0.960 ;
        RECT  4.400 0.345 4.470 1.050 ;
        RECT  3.945 0.980 4.400 1.050 ;
        RECT  4.300 0.810 4.330 0.910 ;
        RECT  4.230 0.205 4.300 0.910 ;
        RECT  4.105 0.365 4.160 0.905 ;
        RECT  4.090 0.185 4.105 0.905 ;
        RECT  4.035 0.185 4.090 0.445 ;
        RECT  4.030 0.835 4.090 0.905 ;
        RECT  3.945 0.520 4.010 0.640 ;
        RECT  3.875 0.520 3.945 1.050 ;
        RECT  2.755 0.850 3.875 0.920 ;
        RECT  3.340 0.990 3.460 1.075 ;
        RECT  3.140 0.210 3.400 0.280 ;
        RECT  3.140 0.710 3.350 0.780 ;
        RECT  2.330 0.990 3.340 1.060 ;
        RECT  3.070 0.210 3.140 0.780 ;
        RECT  2.605 0.210 3.070 0.280 ;
        RECT  2.990 0.520 3.070 0.640 ;
        RECT  2.920 0.350 3.000 0.450 ;
        RECT  2.850 0.350 2.920 0.780 ;
        RECT  2.755 0.350 2.780 0.470 ;
        RECT  2.685 0.350 2.755 0.920 ;
        RECT  2.590 0.850 2.685 0.920 ;
        RECT  2.535 0.210 2.605 0.630 ;
        RECT  2.505 0.560 2.535 0.630 ;
        RECT  2.435 0.560 2.505 0.890 ;
        RECT  2.330 0.195 2.395 0.495 ;
        RECT  2.325 0.195 2.330 1.060 ;
        RECT  2.260 0.425 2.325 1.060 ;
        RECT  2.120 0.210 2.190 1.000 ;
        RECT  1.600 0.210 2.120 0.280 ;
        RECT  2.050 0.930 2.120 1.000 ;
        RECT  2.010 0.520 2.050 0.640 ;
        RECT  2.000 0.355 2.010 0.640 ;
        RECT  1.965 0.355 2.000 0.805 ;
        RECT  1.930 0.355 1.965 1.035 ;
        RECT  1.880 0.355 1.930 0.425 ;
        RECT  1.895 0.735 1.930 1.035 ;
        RECT  1.775 0.520 1.860 0.640 ;
        RECT  1.705 0.520 1.775 1.050 ;
        RECT  1.230 0.980 1.705 1.050 ;
        RECT  1.525 0.210 1.600 0.910 ;
        RECT  1.515 0.520 1.525 0.910 ;
        RECT  1.450 0.520 1.515 0.640 ;
        RECT  1.380 0.210 1.420 0.330 ;
        RECT  1.380 0.740 1.405 0.860 ;
        RECT  1.310 0.210 1.380 0.860 ;
        RECT  0.480 0.210 1.310 0.280 ;
        RECT  1.150 0.350 1.230 1.050 ;
        RECT  0.790 0.350 1.070 0.420 ;
        RECT  0.975 0.845 1.045 1.025 ;
        RECT  0.790 0.845 0.975 0.920 ;
        RECT  0.720 0.350 0.790 0.920 ;
        RECT  0.590 0.350 0.720 0.420 ;
        RECT  0.685 0.765 0.720 0.920 ;
        RECT  0.615 0.765 0.685 1.025 ;
        RECT  0.480 0.520 0.635 0.640 ;
        RECT  0.410 0.210 0.480 0.790 ;
        RECT  0.305 0.395 0.410 0.465 ;
        RECT  0.305 0.720 0.410 0.790 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.720 0.305 1.035 ;
    END
END CMPE42D2BWP

MACRO DCAP16BWP
    CLASS CORE ;
    FOREIGN DCAP16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.375 -0.115 2.240 0.115 ;
        RECT  1.305 -0.115 1.375 0.360 ;
        RECT  0.760 -0.115 1.305 0.115 ;
        RECT  0.680 -0.115 0.760 0.360 ;
        RECT  0.145 -0.115 0.680 0.115 ;
        RECT  0.065 -0.115 0.145 0.360 ;
        RECT  0.000 -0.115 0.065 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.375 1.145 2.240 1.375 ;
        RECT  1.305 0.760 1.375 1.375 ;
        RECT  0.760 1.145 1.305 1.375 ;
        RECT  0.680 0.770 0.760 1.375 ;
        RECT  0.145 1.145 0.680 1.375 ;
        RECT  0.065 0.760 0.145 1.375 ;
        RECT  0.000 1.145 0.065 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.110 0.210 2.190 0.710 ;
        RECT  2.110 0.790 2.190 1.060 ;
        RECT  1.860 0.630 2.110 0.710 ;
        RECT  1.790 0.790 2.110 0.870 ;
        RECT  1.710 0.430 1.790 0.870 ;
        RECT  0.250 0.430 1.710 0.510 ;
    END
END DCAP16BWP

MACRO DCAP32BWP
    CLASS CORE ;
    FOREIGN DCAP32BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 -0.115 4.480 0.115 ;
        RECT  3.345 -0.115 3.415 0.360 ;
        RECT  2.595 -0.115 3.345 0.115 ;
        RECT  2.525 -0.115 2.595 0.360 ;
        RECT  1.775 -0.115 2.525 0.115 ;
        RECT  1.705 -0.115 1.775 0.360 ;
        RECT  0.955 -0.115 1.705 0.115 ;
        RECT  0.885 -0.115 0.955 0.360 ;
        RECT  0.135 -0.115 0.885 0.115 ;
        RECT  0.065 -0.115 0.135 0.360 ;
        RECT  0.000 -0.115 0.065 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.145 4.480 1.375 ;
        RECT  3.345 0.760 3.415 1.375 ;
        RECT  2.595 1.145 3.345 1.375 ;
        RECT  2.525 0.760 2.595 1.375 ;
        RECT  1.775 1.145 2.525 1.375 ;
        RECT  1.705 0.760 1.775 1.375 ;
        RECT  0.955 1.145 1.705 1.375 ;
        RECT  0.885 0.760 0.955 1.375 ;
        RECT  0.135 1.145 0.885 1.375 ;
        RECT  0.065 0.760 0.135 1.375 ;
        RECT  0.000 1.145 0.065 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.200 4.430 0.710 ;
        RECT  4.350 0.790 4.430 1.060 ;
        RECT  4.090 0.630 4.350 0.710 ;
        RECT  4.015 0.790 4.350 0.870 ;
        RECT  3.935 0.430 4.015 0.870 ;
        RECT  0.200 0.430 3.935 0.510 ;
    END
END DCAP32BWP

MACRO DCAP4BWP
    CLASS CORE ;
    FOREIGN DCAP4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 -0.115 0.560 0.115 ;
        RECT  0.250 -0.115 0.330 0.350 ;
        RECT  0.130 -0.115 0.250 0.115 ;
        RECT  0.050 -0.115 0.130 0.350 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 0.560 1.375 ;
        RECT  0.250 0.945 0.330 1.375 ;
        RECT  0.130 1.145 0.250 1.375 ;
        RECT  0.050 0.945 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.430 0.210 0.510 0.700 ;
        RECT  0.430 0.785 0.510 1.075 ;
        RECT  0.330 0.620 0.430 0.700 ;
        RECT  0.225 0.785 0.430 0.865 ;
        RECT  0.155 0.440 0.225 0.865 ;
    END
END DCAP4BWP

MACRO DCAP64BWP
    CLASS CORE ;
    FOREIGN DCAP64BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.885 -0.115 8.960 0.115 ;
        RECT  7.815 -0.115 7.885 0.360 ;
        RECT  7.115 -0.115 7.815 0.115 ;
        RECT  7.045 -0.115 7.115 0.360 ;
        RECT  6.345 -0.115 7.045 0.115 ;
        RECT  6.275 -0.115 6.345 0.360 ;
        RECT  5.575 -0.115 6.275 0.115 ;
        RECT  5.505 -0.115 5.575 0.360 ;
        RECT  4.805 -0.115 5.505 0.115 ;
        RECT  4.735 -0.115 4.805 0.360 ;
        RECT  4.035 -0.115 4.735 0.115 ;
        RECT  3.965 -0.115 4.035 0.360 ;
        RECT  3.265 -0.115 3.965 0.115 ;
        RECT  3.195 -0.115 3.265 0.360 ;
        RECT  2.495 -0.115 3.195 0.115 ;
        RECT  2.425 -0.115 2.495 0.360 ;
        RECT  1.725 -0.115 2.425 0.115 ;
        RECT  1.655 -0.115 1.725 0.360 ;
        RECT  0.955 -0.115 1.655 0.115 ;
        RECT  0.885 -0.115 0.955 0.360 ;
        RECT  0.185 -0.115 0.885 0.115 ;
        RECT  0.115 -0.115 0.185 0.360 ;
        RECT  0.000 -0.115 0.115 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.885 1.145 8.960 1.375 ;
        RECT  7.815 0.760 7.885 1.375 ;
        RECT  7.115 1.145 7.815 1.375 ;
        RECT  7.045 0.760 7.115 1.375 ;
        RECT  6.345 1.145 7.045 1.375 ;
        RECT  6.275 0.760 6.345 1.375 ;
        RECT  5.575 1.145 6.275 1.375 ;
        RECT  5.505 0.760 5.575 1.375 ;
        RECT  4.805 1.145 5.505 1.375 ;
        RECT  4.735 0.760 4.805 1.375 ;
        RECT  4.035 1.145 4.735 1.375 ;
        RECT  3.965 0.760 4.035 1.375 ;
        RECT  3.265 1.145 3.965 1.375 ;
        RECT  3.195 0.760 3.265 1.375 ;
        RECT  2.495 1.145 3.195 1.375 ;
        RECT  2.425 0.760 2.495 1.375 ;
        RECT  1.725 1.145 2.425 1.375 ;
        RECT  1.655 0.760 1.725 1.375 ;
        RECT  0.955 1.145 1.655 1.375 ;
        RECT  0.885 0.760 0.955 1.375 ;
        RECT  0.185 1.145 0.885 1.375 ;
        RECT  0.115 0.760 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.810 0.210 8.890 0.710 ;
        RECT  8.810 0.810 8.890 1.070 ;
        RECT  8.440 0.630 8.810 0.710 ;
        RECT  8.370 0.810 8.810 0.890 ;
        RECT  8.290 0.430 8.370 0.890 ;
        RECT  0.300 0.430 8.290 0.510 ;
    END
END DCAP64BWP

MACRO DCAP8BWP
    CLASS CORE ;
    FOREIGN DCAP8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.145 -0.115 1.120 0.115 ;
        RECT  0.065 -0.115 0.145 0.360 ;
        RECT  0.000 -0.115 0.065 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.145 1.145 1.120 1.375 ;
        RECT  0.065 0.770 0.145 1.375 ;
        RECT  0.000 1.145 0.065 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.210 1.070 0.710 ;
        RECT  0.990 0.790 1.070 1.050 ;
        RECT  0.740 0.630 0.990 0.710 ;
        RECT  0.670 0.790 0.990 0.870 ;
        RECT  0.590 0.430 0.670 0.870 ;
        RECT  0.250 0.430 0.590 0.510 ;
    END
END DCAP8BWP

MACRO DCAPBWP
    CLASS CORE ;
    FOREIGN DCAPBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.115 0.420 0.115 ;
        RECT  0.115 -0.115 0.185 0.345 ;
        RECT  0.000 -0.115 0.115 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.145 0.420 1.375 ;
        RECT  0.115 0.915 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.205 0.370 0.695 ;
        RECT  0.295 0.775 0.365 1.070 ;
        RECT  0.190 0.625 0.300 0.695 ;
        RECT  0.120 0.775 0.295 0.845 ;
        RECT  0.120 0.445 0.230 0.515 ;
        RECT  0.050 0.445 0.120 0.845 ;
    END
END DCAPBWP

MACRO DCAPX16BWP
    CLASS CORE ;
    FOREIGN DCAPX16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.165 -0.115 2.240 0.115 ;
        RECT  2.095 -0.115 2.165 0.370 ;
        RECT  1.565 -0.115 2.095 0.115 ;
        RECT  1.495 -0.115 1.565 0.370 ;
        RECT  0.955 -0.115 1.495 0.115 ;
        RECT  0.885 -0.115 0.955 0.370 ;
        RECT  0.355 -0.115 0.885 0.115 ;
        RECT  0.285 -0.115 0.355 0.370 ;
        RECT  0.215 -0.115 0.285 0.115 ;
        RECT  0.145 -0.115 0.215 0.190 ;
        RECT  0.000 -0.115 0.145 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.095 1.145 2.240 1.375 ;
        RECT  2.025 1.070 2.095 1.375 ;
        RECT  1.955 1.145 2.025 1.375 ;
        RECT  1.885 0.775 1.955 1.375 ;
        RECT  1.355 1.145 1.885 1.375 ;
        RECT  1.285 0.775 1.355 1.375 ;
        RECT  0.745 1.145 1.285 1.375 ;
        RECT  0.675 0.775 0.745 1.375 ;
        RECT  0.145 1.145 0.675 1.375 ;
        RECT  0.075 0.775 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
END DCAPX16BWP

MACRO DCAPX32BWP
    CLASS CORE ;
    FOREIGN DCAPX32BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.405 -0.115 4.480 0.115 ;
        RECT  4.335 -0.115 4.405 0.370 ;
        RECT  3.610 -0.115 4.335 0.115 ;
        RECT  3.530 -0.115 3.610 0.370 ;
        RECT  2.795 -0.115 3.530 0.115 ;
        RECT  2.725 -0.115 2.795 0.370 ;
        RECT  1.985 -0.115 2.725 0.115 ;
        RECT  1.915 -0.115 1.985 0.370 ;
        RECT  1.175 -0.115 1.915 0.115 ;
        RECT  1.105 -0.115 1.175 0.370 ;
        RECT  0.375 -0.115 1.105 0.115 ;
        RECT  0.305 -0.115 0.375 0.370 ;
        RECT  0.235 -0.115 0.305 0.115 ;
        RECT  0.165 -0.115 0.235 0.190 ;
        RECT  0.000 -0.115 0.165 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.315 1.145 4.480 1.375 ;
        RECT  4.245 1.070 4.315 1.375 ;
        RECT  4.175 1.145 4.245 1.375 ;
        RECT  4.105 0.785 4.175 1.375 ;
        RECT  3.375 1.145 4.105 1.375 ;
        RECT  3.305 0.785 3.375 1.375 ;
        RECT  2.565 1.145 3.305 1.375 ;
        RECT  2.495 0.785 2.565 1.375 ;
        RECT  1.755 1.145 2.495 1.375 ;
        RECT  1.685 0.785 1.755 1.375 ;
        RECT  0.950 1.145 1.685 1.375 ;
        RECT  0.870 0.785 0.950 1.375 ;
        RECT  0.145 1.145 0.870 1.375 ;
        RECT  0.075 0.785 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
END DCAPX32BWP

MACRO DCAPX4BWP
    CLASS CORE ;
    FOREIGN DCAPX4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.505 -0.115 0.560 0.115 ;
        RECT  0.435 -0.115 0.505 0.490 ;
        RECT  0.330 -0.115 0.435 0.115 ;
        RECT  0.260 -0.115 0.330 0.490 ;
        RECT  0.190 -0.115 0.260 0.115 ;
        RECT  0.120 -0.115 0.190 0.190 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.145 0.560 1.375 ;
        RECT  0.370 1.070 0.440 1.375 ;
        RECT  0.300 1.145 0.370 1.375 ;
        RECT  0.230 0.770 0.300 1.375 ;
        RECT  0.125 1.145 0.230 1.375 ;
        RECT  0.055 0.770 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
END DCAPX4BWP

MACRO DCAPX64BWP
    CLASS CORE ;
    FOREIGN DCAPX64BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.885 -0.115 8.960 0.115 ;
        RECT  8.815 -0.115 8.885 0.370 ;
        RECT  8.125 -0.115 8.815 0.115 ;
        RECT  8.055 -0.115 8.125 0.370 ;
        RECT  7.355 -0.115 8.055 0.115 ;
        RECT  7.285 -0.115 7.355 0.370 ;
        RECT  6.585 -0.115 7.285 0.115 ;
        RECT  6.515 -0.115 6.585 0.370 ;
        RECT  5.815 -0.115 6.515 0.115 ;
        RECT  5.745 -0.115 5.815 0.370 ;
        RECT  5.045 -0.115 5.745 0.115 ;
        RECT  4.975 -0.115 5.045 0.370 ;
        RECT  4.275 -0.115 4.975 0.115 ;
        RECT  4.205 -0.115 4.275 0.370 ;
        RECT  3.505 -0.115 4.205 0.115 ;
        RECT  3.435 -0.115 3.505 0.370 ;
        RECT  2.735 -0.115 3.435 0.115 ;
        RECT  2.665 -0.115 2.735 0.370 ;
        RECT  1.965 -0.115 2.665 0.115 ;
        RECT  1.895 -0.115 1.965 0.370 ;
        RECT  1.195 -0.115 1.895 0.115 ;
        RECT  1.125 -0.115 1.195 0.370 ;
        RECT  0.435 -0.115 1.125 0.115 ;
        RECT  0.365 -0.115 0.435 0.370 ;
        RECT  0.285 -0.115 0.365 0.115 ;
        RECT  0.205 -0.115 0.285 0.190 ;
        RECT  0.000 -0.115 0.205 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.755 1.145 8.960 1.375 ;
        RECT  8.675 1.080 8.755 1.375 ;
        RECT  8.605 1.145 8.675 1.375 ;
        RECT  8.535 0.775 8.605 1.375 ;
        RECT  7.835 1.145 8.535 1.375 ;
        RECT  7.765 0.775 7.835 1.375 ;
        RECT  7.065 1.145 7.765 1.375 ;
        RECT  6.995 0.775 7.065 1.375 ;
        RECT  6.295 1.145 6.995 1.375 ;
        RECT  6.225 0.775 6.295 1.375 ;
        RECT  5.525 1.145 6.225 1.375 ;
        RECT  5.455 0.775 5.525 1.375 ;
        RECT  4.755 1.145 5.455 1.375 ;
        RECT  4.685 0.775 4.755 1.375 ;
        RECT  3.985 1.145 4.685 1.375 ;
        RECT  3.915 0.775 3.985 1.375 ;
        RECT  3.215 1.145 3.915 1.375 ;
        RECT  3.145 0.775 3.215 1.375 ;
        RECT  2.445 1.145 3.145 1.375 ;
        RECT  2.375 0.775 2.445 1.375 ;
        RECT  1.675 1.145 2.375 1.375 ;
        RECT  1.605 0.775 1.675 1.375 ;
        RECT  0.905 1.145 1.605 1.375 ;
        RECT  0.835 0.775 0.905 1.375 ;
        RECT  0.145 1.145 0.835 1.375 ;
        RECT  0.075 0.775 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
END DCAPX64BWP

MACRO DCAPX8BWP
    CLASS CORE ;
    FOREIGN DCAPX8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.045 -0.115 1.120 0.115 ;
        RECT  0.975 -0.115 1.045 0.370 ;
        RECT  0.345 -0.115 0.975 0.115 ;
        RECT  0.275 -0.115 0.345 0.370 ;
        RECT  0.205 -0.115 0.275 0.115 ;
        RECT  0.135 -0.115 0.205 0.190 ;
        RECT  0.000 -0.115 0.135 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 1.145 1.120 1.375 ;
        RECT  0.915 1.070 0.985 1.375 ;
        RECT  0.845 1.145 0.915 1.375 ;
        RECT  0.775 0.770 0.845 1.375 ;
        RECT  0.145 1.145 0.775 1.375 ;
        RECT  0.075 0.770 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
END DCAPX8BWP

MACRO DCCKBD12BWP
    CLASS CORE ;
    FOREIGN DCCKBD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.5987 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 0.195 2.890 0.450 ;
        RECT  2.135 0.725 2.885 0.955 ;
        RECT  2.510 0.290 2.810 0.450 ;
        RECT  2.430 0.190 2.510 0.450 ;
        RECT  2.150 0.290 2.430 0.450 ;
        RECT  2.135 0.190 2.150 0.450 ;
        RECT  2.070 0.190 2.135 0.955 ;
        RECT  1.790 0.290 2.070 0.955 ;
        RECT  1.785 0.190 1.790 0.955 ;
        RECT  1.710 0.190 1.785 0.450 ;
        RECT  0.970 0.725 1.785 0.955 ;
        RECT  1.430 0.290 1.710 0.450 ;
        RECT  1.350 0.190 1.430 0.450 ;
        RECT  1.070 0.290 1.350 0.450 ;
        RECT  0.990 0.190 1.070 0.450 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1088 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.455 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.640 -0.115 5.880 0.115 ;
        RECT  5.560 -0.115 5.640 0.350 ;
        RECT  5.000 -0.115 5.560 0.115 ;
        RECT  4.920 -0.115 5.000 0.350 ;
        RECT  4.360 -0.115 4.920 0.115 ;
        RECT  4.280 -0.115 4.360 0.350 ;
        RECT  3.720 -0.115 4.280 0.115 ;
        RECT  3.640 -0.115 3.720 0.350 ;
        RECT  3.085 -0.115 3.640 0.115 ;
        RECT  3.005 -0.115 3.085 0.350 ;
        RECT  0.880 -0.115 3.005 0.115 ;
        RECT  0.800 -0.115 0.880 0.450 ;
        RECT  0.130 -0.115 0.800 0.115 ;
        RECT  0.050 -0.115 0.130 0.335 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.670 1.145 5.880 1.375 ;
        RECT  5.530 0.945 5.670 1.375 ;
        RECT  4.995 1.145 5.530 1.375 ;
        RECT  4.925 0.770 4.995 1.375 ;
        RECT  4.360 1.145 4.925 1.375 ;
        RECT  4.280 0.770 4.360 1.375 ;
        RECT  3.720 1.145 4.280 1.375 ;
        RECT  3.640 0.770 3.720 1.375 ;
        RECT  3.085 1.145 3.640 1.375 ;
        RECT  3.005 0.770 3.085 1.375 ;
        RECT  2.720 1.145 3.005 1.375 ;
        RECT  2.600 1.025 2.720 1.375 ;
        RECT  2.350 1.145 2.600 1.375 ;
        RECT  2.230 1.025 2.350 1.375 ;
        RECT  1.995 1.145 2.230 1.375 ;
        RECT  1.865 1.025 1.995 1.375 ;
        RECT  1.630 1.145 1.865 1.375 ;
        RECT  1.510 1.025 1.630 1.375 ;
        RECT  1.270 1.145 1.510 1.375 ;
        RECT  1.150 1.025 1.270 1.375 ;
        RECT  0.880 1.145 1.150 1.375 ;
        RECT  0.800 0.735 0.880 1.375 ;
        RECT  0.520 1.145 0.800 1.375 ;
        RECT  0.400 0.885 0.520 1.375 ;
        RECT  0.130 1.145 0.400 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.810 0.195 2.890 0.450 ;
        RECT  2.205 0.725 2.885 0.955 ;
        RECT  2.510 0.290 2.810 0.450 ;
        RECT  2.430 0.190 2.510 0.450 ;
        RECT  2.205 0.290 2.430 0.450 ;
        RECT  1.710 0.190 1.715 0.450 ;
        RECT  0.970 0.725 1.715 0.955 ;
        RECT  1.430 0.290 1.710 0.450 ;
        RECT  1.350 0.190 1.430 0.450 ;
        RECT  1.070 0.290 1.350 0.450 ;
        RECT  0.990 0.190 1.070 0.450 ;
        RECT  5.750 0.230 5.830 0.710 ;
        RECT  5.750 0.790 5.830 0.975 ;
        RECT  0.220 0.715 0.320 1.035 ;
        RECT  5.610 0.630 5.750 0.710 ;
        RECT  5.530 0.790 5.750 0.870 ;
        RECT  5.450 0.430 5.530 0.870 ;
        RECT  3.130 0.430 5.450 0.510 ;
        RECT  2.235 0.535 2.890 0.605 ;
        RECT  0.710 0.535 1.685 0.605 ;
        RECT  0.700 0.305 0.710 0.605 ;
        RECT  0.600 0.305 0.700 1.035 ;
        RECT  0.210 0.305 0.600 0.405 ;
        RECT  0.320 0.715 0.600 0.815 ;
    END
END DCCKBD12BWP

MACRO DCCKBD16BWP
    CLASS CORE ;
    FOREIGN DCCKBD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.7892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.195 3.730 0.455 ;
        RECT  2.695 0.725 3.725 0.955 ;
        RECT  3.370 0.295 3.650 0.455 ;
        RECT  3.290 0.195 3.370 0.455 ;
        RECT  3.010 0.295 3.290 0.455 ;
        RECT  2.930 0.195 3.010 0.455 ;
        RECT  2.695 0.295 2.930 0.455 ;
        RECT  2.650 0.295 2.695 0.955 ;
        RECT  2.555 0.195 2.650 0.955 ;
        RECT  2.345 0.295 2.555 0.955 ;
        RECT  2.290 0.295 2.345 0.455 ;
        RECT  1.110 0.725 2.345 0.955 ;
        RECT  2.210 0.195 2.290 0.455 ;
        RECT  1.930 0.295 2.210 0.455 ;
        RECT  1.850 0.195 1.930 0.455 ;
        RECT  1.570 0.295 1.850 0.455 ;
        RECT  1.490 0.195 1.570 0.455 ;
        RECT  1.210 0.295 1.490 0.455 ;
        RECT  1.130 0.195 1.210 0.455 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1360 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.625 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 -0.115 7.560 0.115 ;
        RECT  7.240 -0.115 7.320 0.350 ;
        RECT  6.640 -0.115 7.240 0.115 ;
        RECT  6.560 -0.115 6.640 0.350 ;
        RECT  5.960 -0.115 6.560 0.115 ;
        RECT  5.880 -0.115 5.960 0.350 ;
        RECT  5.280 -0.115 5.880 0.115 ;
        RECT  5.200 -0.115 5.280 0.350 ;
        RECT  4.600 -0.115 5.200 0.115 ;
        RECT  4.520 -0.115 4.600 0.350 ;
        RECT  3.925 -0.115 4.520 0.115 ;
        RECT  3.845 -0.115 3.925 0.350 ;
        RECT  1.030 -0.115 3.845 0.115 ;
        RECT  0.950 -0.115 1.030 0.455 ;
        RECT  0.000 -0.115 0.950 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.345 1.145 7.560 1.375 ;
        RECT  7.215 0.945 7.345 1.375 ;
        RECT  6.640 1.145 7.215 1.375 ;
        RECT  6.560 0.770 6.640 1.375 ;
        RECT  5.960 1.145 6.560 1.375 ;
        RECT  5.880 0.770 5.960 1.375 ;
        RECT  5.275 1.145 5.880 1.375 ;
        RECT  5.205 0.770 5.275 1.375 ;
        RECT  4.595 1.145 5.205 1.375 ;
        RECT  4.525 0.770 4.595 1.375 ;
        RECT  3.925 1.145 4.525 1.375 ;
        RECT  3.845 0.770 3.925 1.375 ;
        RECT  3.570 1.145 3.845 1.375 ;
        RECT  3.450 1.025 3.570 1.375 ;
        RECT  3.210 1.145 3.450 1.375 ;
        RECT  3.090 1.025 3.210 1.375 ;
        RECT  2.850 1.145 3.090 1.375 ;
        RECT  2.730 1.025 2.850 1.375 ;
        RECT  2.490 1.145 2.730 1.375 ;
        RECT  2.370 1.025 2.490 1.375 ;
        RECT  2.130 1.145 2.370 1.375 ;
        RECT  2.010 1.025 2.130 1.375 ;
        RECT  1.770 1.145 2.010 1.375 ;
        RECT  1.650 1.025 1.770 1.375 ;
        RECT  1.410 1.145 1.650 1.375 ;
        RECT  1.290 1.025 1.410 1.375 ;
        RECT  1.030 1.145 1.290 1.375 ;
        RECT  0.950 0.695 1.030 1.375 ;
        RECT  0.690 1.145 0.950 1.375 ;
        RECT  0.570 0.890 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.195 3.730 0.455 ;
        RECT  2.765 0.725 3.725 0.955 ;
        RECT  3.370 0.295 3.650 0.455 ;
        RECT  3.290 0.195 3.370 0.455 ;
        RECT  3.010 0.295 3.290 0.455 ;
        RECT  2.930 0.195 3.010 0.455 ;
        RECT  2.765 0.295 2.930 0.455 ;
        RECT  2.210 0.195 2.275 0.455 ;
        RECT  1.110 0.725 2.275 0.955 ;
        RECT  1.930 0.295 2.210 0.455 ;
        RECT  1.850 0.195 1.930 0.455 ;
        RECT  1.570 0.295 1.850 0.455 ;
        RECT  1.490 0.195 1.570 0.455 ;
        RECT  1.210 0.295 1.490 0.455 ;
        RECT  1.130 0.195 1.210 0.455 ;
        RECT  7.430 0.240 7.510 0.710 ;
        RECT  7.430 0.790 7.510 0.975 ;
        RECT  7.290 0.630 7.430 0.710 ;
        RECT  7.210 0.790 7.430 0.870 ;
        RECT  7.130 0.430 7.210 0.870 ;
        RECT  3.950 0.430 7.130 0.510 ;
        RECT  2.810 0.535 3.540 0.605 ;
        RECT  0.870 0.535 2.210 0.605 ;
        RECT  0.860 0.305 0.870 0.605 ;
        RECT  0.760 0.305 0.860 1.030 ;
        RECT  0.130 0.305 0.760 0.395 ;
        RECT  0.500 0.720 0.760 0.820 ;
        RECT  0.400 0.720 0.500 1.030 ;
        RECT  0.140 0.720 0.400 0.820 ;
        RECT  0.050 0.720 0.140 1.030 ;
        RECT  0.050 0.225 0.130 0.395 ;
    END
END DCCKBD16BWP

MACRO DCCKBD20BWP
    CLASS CORE ;
    FOREIGN DCCKBD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.710 4.330 0.940 ;
        RECT  4.220 0.190 4.300 0.450 ;
        RECT  3.910 0.310 4.220 0.450 ;
        RECT  3.830 0.190 3.910 0.450 ;
        RECT  3.550 0.310 3.830 0.450 ;
        RECT  3.470 0.190 3.550 0.450 ;
        RECT  3.190 0.310 3.470 0.450 ;
        RECT  3.115 0.190 3.190 0.450 ;
        RECT  3.110 0.190 3.115 0.940 ;
        RECT  2.830 0.310 3.110 0.940 ;
        RECT  2.765 0.190 2.830 0.940 ;
        RECT  2.750 0.190 2.765 0.450 ;
        RECT  1.290 0.710 2.765 0.940 ;
        RECT  2.470 0.310 2.750 0.450 ;
        RECT  2.390 0.190 2.470 0.450 ;
        RECT  2.110 0.310 2.390 0.450 ;
        RECT  2.030 0.190 2.110 0.450 ;
        RECT  1.750 0.310 2.030 0.450 ;
        RECT  1.670 0.190 1.750 0.450 ;
        RECT  1.390 0.310 1.670 0.450 ;
        RECT  1.310 0.190 1.390 0.450 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1632 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.785 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.980 -0.115 9.240 0.115 ;
        RECT  8.900 -0.115 8.980 0.350 ;
        RECT  8.260 -0.115 8.900 0.115 ;
        RECT  8.180 -0.115 8.260 0.350 ;
        RECT  7.560 -0.115 8.180 0.115 ;
        RECT  7.480 -0.115 7.560 0.350 ;
        RECT  6.860 -0.115 7.480 0.115 ;
        RECT  6.780 -0.115 6.860 0.350 ;
        RECT  6.160 -0.115 6.780 0.115 ;
        RECT  6.080 -0.115 6.160 0.350 ;
        RECT  5.460 -0.115 6.080 0.115 ;
        RECT  5.380 -0.115 5.460 0.350 ;
        RECT  4.765 -0.115 5.380 0.115 ;
        RECT  4.685 -0.115 4.765 0.350 ;
        RECT  4.490 -0.115 4.685 0.115 ;
        RECT  4.410 -0.115 4.490 0.450 ;
        RECT  4.120 -0.115 4.410 0.115 ;
        RECT  4.000 -0.115 4.120 0.240 ;
        RECT  3.750 -0.115 4.000 0.115 ;
        RECT  3.630 -0.115 3.750 0.240 ;
        RECT  3.390 -0.115 3.630 0.115 ;
        RECT  3.270 -0.115 3.390 0.240 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.240 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.240 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.240 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.240 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.240 ;
        RECT  1.210 -0.115 1.470 0.115 ;
        RECT  1.130 -0.115 1.210 0.450 ;
        RECT  0.130 -0.115 1.130 0.115 ;
        RECT  0.050 -0.115 0.130 0.350 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.015 1.145 9.240 1.375 ;
        RECT  8.865 0.945 9.015 1.375 ;
        RECT  8.265 1.145 8.865 1.375 ;
        RECT  8.185 0.770 8.265 1.375 ;
        RECT  7.560 1.145 8.185 1.375 ;
        RECT  7.480 0.770 7.560 1.375 ;
        RECT  6.860 1.145 7.480 1.375 ;
        RECT  6.780 0.770 6.860 1.375 ;
        RECT  6.165 1.145 6.780 1.375 ;
        RECT  6.075 0.770 6.165 1.375 ;
        RECT  5.465 1.145 6.075 1.375 ;
        RECT  5.375 0.770 5.465 1.375 ;
        RECT  4.765 1.145 5.375 1.375 ;
        RECT  4.685 0.770 4.765 1.375 ;
        RECT  4.485 1.145 4.685 1.375 ;
        RECT  4.415 0.750 4.485 1.375 ;
        RECT  4.120 1.145 4.415 1.375 ;
        RECT  4.000 1.010 4.120 1.375 ;
        RECT  3.750 1.145 4.000 1.375 ;
        RECT  3.630 1.010 3.750 1.375 ;
        RECT  3.390 1.145 3.630 1.375 ;
        RECT  3.270 1.010 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 1.010 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.010 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.010 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 1.010 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 1.010 1.590 1.375 ;
        RECT  1.210 1.145 1.470 1.375 ;
        RECT  1.130 0.695 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.910 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.910 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.705 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.710 4.330 0.940 ;
        RECT  4.220 0.190 4.300 0.450 ;
        RECT  3.910 0.310 4.220 0.450 ;
        RECT  3.830 0.190 3.910 0.450 ;
        RECT  3.550 0.310 3.830 0.450 ;
        RECT  3.470 0.190 3.550 0.450 ;
        RECT  3.190 0.310 3.470 0.450 ;
        RECT  3.185 0.190 3.190 0.450 ;
        RECT  2.470 0.310 2.695 0.450 ;
        RECT  1.290 0.710 2.695 0.940 ;
        RECT  2.390 0.190 2.470 0.450 ;
        RECT  2.110 0.310 2.390 0.450 ;
        RECT  2.030 0.190 2.110 0.450 ;
        RECT  1.750 0.310 2.030 0.450 ;
        RECT  1.670 0.190 1.750 0.450 ;
        RECT  1.390 0.310 1.670 0.450 ;
        RECT  1.310 0.190 1.390 0.450 ;
        RECT  9.110 0.240 9.190 0.710 ;
        RECT  9.110 0.790 9.190 0.975 ;
        RECT  8.970 0.630 9.110 0.710 ;
        RECT  8.860 0.790 9.110 0.870 ;
        RECT  8.780 0.430 8.860 0.870 ;
        RECT  4.805 0.430 8.780 0.510 ;
        RECT  3.245 0.525 4.295 0.595 ;
        RECT  1.050 0.525 2.635 0.595 ;
        RECT  0.940 0.290 1.050 1.035 ;
        RECT  0.210 0.290 0.940 0.390 ;
        RECT  0.680 0.740 0.940 0.840 ;
        RECT  0.580 0.740 0.680 1.035 ;
        RECT  0.320 0.740 0.580 0.840 ;
        RECT  0.220 0.740 0.320 1.035 ;
    END
END DCCKBD20BWP

MACRO DCCKBD4BWP
    CLASS CORE ;
    FOREIGN DCCKBD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1904 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.235 1.025 0.495 ;
        RECT  1.015 0.700 1.025 1.050 ;
        RECT  0.955 0.235 1.015 1.050 ;
        RECT  0.805 0.355 0.955 0.820 ;
        RECT  0.665 0.355 0.805 0.475 ;
        RECT  0.665 0.700 0.805 0.820 ;
        RECT  0.595 0.235 0.665 0.475 ;
        RECT  0.595 0.700 0.665 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 -0.115 2.520 0.115 ;
        RECT  2.210 -0.115 2.290 0.350 ;
        RECT  1.400 -0.115 2.210 0.115 ;
        RECT  1.320 -0.115 1.400 0.350 ;
        RECT  1.210 -0.115 1.320 0.115 ;
        RECT  1.130 -0.115 1.210 0.440 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.280 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.365 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.145 2.520 1.375 ;
        RECT  2.170 0.945 2.310 1.375 ;
        RECT  1.400 1.145 2.170 1.375 ;
        RECT  1.320 0.770 1.400 1.375 ;
        RECT  1.210 1.145 1.320 1.375 ;
        RECT  1.130 0.675 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.890 0.870 1.375 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.910 0.490 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.475 ;
        RECT  0.665 0.700 0.735 0.820 ;
        RECT  0.595 0.235 0.665 0.475 ;
        RECT  0.595 0.700 0.665 1.050 ;
        RECT  2.390 0.240 2.470 0.710 ;
        RECT  2.390 0.790 2.470 0.975 ;
        RECT  2.250 0.630 2.390 0.710 ;
        RECT  2.170 0.790 2.390 0.870 ;
        RECT  2.090 0.430 2.170 0.870 ;
        RECT  1.480 0.430 2.090 0.510 ;
        RECT  0.380 0.545 0.650 0.615 ;
        RECT  0.310 0.350 0.380 0.820 ;
        RECT  0.305 0.350 0.310 0.420 ;
        RECT  0.305 0.750 0.310 0.820 ;
        RECT  0.235 0.245 0.305 0.420 ;
        RECT  0.235 0.750 0.305 1.045 ;
    END
END DCCKBD4BWP

MACRO DCCKBD8BWP
    CLASS CORE ;
    FOREIGN DCCKBD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.3808 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.720 2.030 0.950 ;
        RECT  1.930 0.255 2.010 0.455 ;
        RECT  1.630 0.350 1.930 0.455 ;
        RECT  1.575 0.255 1.630 0.455 ;
        RECT  1.550 0.255 1.575 0.950 ;
        RECT  1.250 0.345 1.550 0.950 ;
        RECT  1.225 0.215 1.250 0.950 ;
        RECT  1.170 0.215 1.225 0.455 ;
        RECT  0.770 0.720 1.225 0.950 ;
        RECT  0.870 0.345 1.170 0.455 ;
        RECT  0.790 0.255 0.870 0.455 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0816 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.290 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 -0.115 4.480 0.115 ;
        RECT  4.160 -0.115 4.240 0.350 ;
        RECT  3.620 -0.115 4.160 0.115 ;
        RECT  3.540 -0.115 3.620 0.350 ;
        RECT  3.000 -0.115 3.540 0.115 ;
        RECT  2.920 -0.115 3.000 0.350 ;
        RECT  2.385 -0.115 2.920 0.115 ;
        RECT  2.305 -0.115 2.385 0.350 ;
        RECT  2.190 -0.115 2.305 0.115 ;
        RECT  2.110 -0.115 2.190 0.395 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.720 -0.115 1.840 0.275 ;
        RECT  1.460 -0.115 1.720 0.115 ;
        RECT  1.340 -0.115 1.460 0.275 ;
        RECT  1.080 -0.115 1.340 0.115 ;
        RECT  0.960 -0.115 1.080 0.275 ;
        RECT  0.690 -0.115 0.960 0.115 ;
        RECT  0.610 -0.115 0.690 0.460 ;
        RECT  0.340 -0.115 0.610 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 1.145 4.480 1.375 ;
        RECT  4.130 0.945 4.270 1.375 ;
        RECT  3.615 1.145 4.130 1.375 ;
        RECT  3.545 0.770 3.615 1.375 ;
        RECT  3.000 1.145 3.545 1.375 ;
        RECT  2.920 0.770 3.000 1.375 ;
        RECT  2.385 1.145 2.920 1.375 ;
        RECT  2.305 0.770 2.385 1.375 ;
        RECT  2.190 1.145 2.305 1.375 ;
        RECT  2.110 0.675 2.190 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.720 1.020 1.840 1.375 ;
        RECT  1.460 1.145 1.720 1.375 ;
        RECT  1.340 1.020 1.460 1.375 ;
        RECT  1.080 1.145 1.340 1.375 ;
        RECT  0.960 1.020 1.080 1.375 ;
        RECT  0.690 1.145 0.960 1.375 ;
        RECT  0.610 0.735 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.920 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.720 2.030 0.950 ;
        RECT  1.930 0.255 2.010 0.455 ;
        RECT  1.645 0.350 1.930 0.455 ;
        RECT  0.870 0.345 1.155 0.455 ;
        RECT  0.770 0.720 1.155 0.950 ;
        RECT  0.790 0.255 0.870 0.455 ;
        RECT  4.350 0.230 4.430 0.710 ;
        RECT  4.350 0.790 4.430 0.975 ;
        RECT  4.210 0.630 4.350 0.710 ;
        RECT  4.130 0.790 4.350 0.870 ;
        RECT  4.050 0.430 4.130 0.870 ;
        RECT  2.410 0.430 4.050 0.510 ;
        RECT  1.675 0.545 2.060 0.615 ;
        RECT  0.520 0.545 1.125 0.615 ;
        RECT  0.420 0.255 0.520 1.035 ;
        RECT  0.125 0.345 0.420 0.425 ;
        RECT  0.125 0.740 0.420 0.840 ;
        RECT  0.055 0.265 0.125 0.425 ;
        RECT  0.055 0.740 0.125 1.035 ;
    END
END DCCKBD8BWP

MACRO DCCKND12BWP
    CLASS CORE ;
    FOREIGN DCCKND12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5829 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.715 2.170 0.945 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.325 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.325 1.715 0.465 ;
        RECT  1.355 0.185 1.425 0.465 ;
        RECT  1.295 0.325 1.355 0.465 ;
        RECT  1.065 0.325 1.295 0.945 ;
        RECT  0.995 0.185 1.065 0.945 ;
        RECT  0.945 0.325 0.995 0.945 ;
        RECT  0.705 0.325 0.945 0.465 ;
        RECT  0.210 0.715 0.945 0.945 ;
        RECT  0.635 0.185 0.705 0.465 ;
        RECT  0.345 0.325 0.635 0.465 ;
        RECT  0.275 0.185 0.345 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.845 0.625 ;
        RECT  0.035 0.200 0.125 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.500 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.500 0.350 ;
        RECT  3.840 -0.115 4.420 0.115 ;
        RECT  3.760 -0.115 3.840 0.350 ;
        RECT  3.180 -0.115 3.760 0.115 ;
        RECT  3.100 -0.115 3.180 0.350 ;
        RECT  2.525 -0.115 3.100 0.115 ;
        RECT  2.445 -0.115 2.525 0.350 ;
        RECT  2.330 -0.115 2.445 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.990 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.990 0.255 ;
        RECT  1.630 -0.115 1.870 0.115 ;
        RECT  1.510 -0.115 1.630 0.255 ;
        RECT  1.270 -0.115 1.510 0.115 ;
        RECT  1.150 -0.115 1.270 0.255 ;
        RECT  0.910 -0.115 1.150 0.115 ;
        RECT  0.790 -0.115 0.910 0.255 ;
        RECT  0.550 -0.115 0.790 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.145 4.760 1.375 ;
        RECT  4.385 0.945 4.535 1.375 ;
        RECT  3.840 1.145 4.385 1.375 ;
        RECT  3.760 0.770 3.840 1.375 ;
        RECT  3.175 1.145 3.760 1.375 ;
        RECT  3.105 0.770 3.175 1.375 ;
        RECT  2.525 1.145 3.105 1.375 ;
        RECT  2.445 0.770 2.525 1.375 ;
        RECT  2.330 1.145 2.445 1.375 ;
        RECT  2.250 0.680 2.330 1.375 ;
        RECT  1.990 1.145 2.250 1.375 ;
        RECT  1.870 1.015 1.990 1.375 ;
        RECT  1.620 1.145 1.870 1.375 ;
        RECT  1.500 1.015 1.620 1.375 ;
        RECT  1.250 1.145 1.500 1.375 ;
        RECT  1.130 1.015 1.250 1.375 ;
        RECT  0.880 1.145 1.130 1.375 ;
        RECT  0.760 1.015 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.715 2.170 0.945 ;
        RECT  2.075 0.185 2.145 0.465 ;
        RECT  1.785 0.325 2.075 0.465 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.425 0.325 1.715 0.465 ;
        RECT  1.365 0.185 1.425 0.465 ;
        RECT  0.705 0.325 0.875 0.465 ;
        RECT  0.210 0.715 0.875 0.945 ;
        RECT  0.635 0.185 0.705 0.465 ;
        RECT  0.345 0.325 0.635 0.465 ;
        RECT  0.275 0.185 0.345 0.465 ;
        RECT  4.610 0.230 4.690 0.710 ;
        RECT  4.610 0.790 4.690 0.975 ;
        RECT  4.530 0.630 4.610 0.710 ;
        RECT  4.450 0.790 4.610 0.870 ;
        RECT  4.370 0.430 4.450 0.870 ;
        RECT  2.570 0.430 4.370 0.510 ;
        RECT  1.415 0.545 2.220 0.615 ;
    END
END DCCKND12BWP

MACRO DCCKND16BWP
    CLASS CORE ;
    FOREIGN DCCKND16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.7620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.715 2.870 0.945 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.125 0.305 2.415 0.465 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.765 0.305 2.055 0.465 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.695 0.185 1.715 0.945 ;
        RECT  1.405 0.305 1.695 0.945 ;
        RECT  1.365 0.185 1.405 0.945 ;
        RECT  1.335 0.185 1.365 0.465 ;
        RECT  0.210 0.715 1.365 0.945 ;
        RECT  1.045 0.305 1.335 0.465 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  0.625 0.305 0.975 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4352 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 1.265 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.920 -0.115 6.160 0.115 ;
        RECT  5.840 -0.115 5.920 0.350 ;
        RECT  5.245 -0.115 5.840 0.115 ;
        RECT  5.165 -0.115 5.245 0.350 ;
        RECT  4.570 -0.115 5.165 0.115 ;
        RECT  4.490 -0.115 4.570 0.350 ;
        RECT  3.895 -0.115 4.490 0.115 ;
        RECT  3.815 -0.115 3.895 0.350 ;
        RECT  3.225 -0.115 3.815 0.115 ;
        RECT  3.145 -0.115 3.225 0.350 ;
        RECT  3.025 -0.115 3.145 0.115 ;
        RECT  2.955 -0.115 3.025 0.475 ;
        RECT  2.690 -0.115 2.955 0.115 ;
        RECT  2.570 -0.115 2.690 0.235 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.235 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.235 ;
        RECT  1.610 -0.115 1.850 0.115 ;
        RECT  1.490 -0.115 1.610 0.235 ;
        RECT  1.250 -0.115 1.490 0.115 ;
        RECT  1.130 -0.115 1.250 0.235 ;
        RECT  0.860 -0.115 1.130 0.115 ;
        RECT  0.740 -0.115 0.860 0.235 ;
        RECT  0.445 -0.115 0.740 0.115 ;
        RECT  0.375 -0.115 0.445 0.460 ;
        RECT  0.000 -0.115 0.375 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.950 1.145 6.160 1.375 ;
        RECT  5.810 0.945 5.950 1.375 ;
        RECT  5.245 1.145 5.810 1.375 ;
        RECT  5.165 0.770 5.245 1.375 ;
        RECT  4.570 1.145 5.165 1.375 ;
        RECT  4.490 0.770 4.570 1.375 ;
        RECT  3.900 1.145 4.490 1.375 ;
        RECT  3.810 0.770 3.900 1.375 ;
        RECT  3.225 1.145 3.810 1.375 ;
        RECT  3.145 0.770 3.225 1.375 ;
        RECT  3.030 1.145 3.145 1.375 ;
        RECT  2.950 0.675 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 1.015 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.015 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.015 1.970 1.375 ;
        RECT  1.610 1.145 1.850 1.375 ;
        RECT  1.490 1.015 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 1.015 1.250 1.375 ;
        RECT  0.880 1.145 1.130 1.375 ;
        RECT  0.760 1.015 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.715 2.870 0.945 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.485 0.305 2.775 0.465 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.125 0.305 2.415 0.465 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.785 0.305 2.055 0.465 ;
        RECT  1.045 0.305 1.295 0.465 ;
        RECT  0.210 0.715 1.295 0.945 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  0.625 0.305 0.975 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        RECT  6.030 0.230 6.110 0.710 ;
        RECT  6.030 0.790 6.110 0.975 ;
        RECT  5.890 0.630 6.030 0.710 ;
        RECT  5.810 0.790 6.030 0.870 ;
        RECT  5.730 0.430 5.810 0.870 ;
        RECT  3.270 0.430 5.730 0.510 ;
        RECT  1.815 0.545 2.805 0.615 ;
    END
END DCCKND16BWP

MACRO DCCKND20BWP
    CLASS CORE ;
    FOREIGN DCCKND20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.9520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.715 3.570 0.945 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.305 2.755 0.465 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.135 0.305 2.395 0.465 ;
        RECT  2.105 0.305 2.135 0.945 ;
        RECT  2.035 0.185 2.105 0.945 ;
        RECT  1.785 0.305 2.035 0.945 ;
        RECT  1.745 0.305 1.785 0.465 ;
        RECT  0.210 0.715 1.785 0.945 ;
        RECT  1.675 0.185 1.745 0.465 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.005 0.305 1.315 0.465 ;
        RECT  0.935 0.185 1.005 0.465 ;
        RECT  0.625 0.305 0.935 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.5440 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 1.685 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.320 -0.115 7.560 0.115 ;
        RECT  7.240 -0.115 7.320 0.350 ;
        RECT  6.640 -0.115 7.240 0.115 ;
        RECT  6.560 -0.115 6.640 0.350 ;
        RECT  5.960 -0.115 6.560 0.115 ;
        RECT  5.880 -0.115 5.960 0.350 ;
        RECT  5.280 -0.115 5.880 0.115 ;
        RECT  5.200 -0.115 5.280 0.350 ;
        RECT  4.600 -0.115 5.200 0.115 ;
        RECT  4.520 -0.115 4.600 0.350 ;
        RECT  3.925 -0.115 4.520 0.115 ;
        RECT  3.845 -0.115 3.925 0.350 ;
        RECT  3.725 -0.115 3.845 0.115 ;
        RECT  3.655 -0.115 3.725 0.465 ;
        RECT  3.390 -0.115 3.655 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.235 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.235 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.235 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.235 ;
        RECT  1.220 -0.115 1.470 0.115 ;
        RECT  1.100 -0.115 1.220 0.235 ;
        RECT  0.840 -0.115 1.100 0.115 ;
        RECT  0.720 -0.115 0.840 0.235 ;
        RECT  0.450 -0.115 0.720 0.115 ;
        RECT  0.370 -0.115 0.450 0.460 ;
        RECT  0.000 -0.115 0.370 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.350 1.145 7.560 1.375 ;
        RECT  7.210 0.945 7.350 1.375 ;
        RECT  6.640 1.145 7.210 1.375 ;
        RECT  6.560 0.770 6.640 1.375 ;
        RECT  5.960 1.145 6.560 1.375 ;
        RECT  5.880 0.770 5.960 1.375 ;
        RECT  5.275 1.145 5.880 1.375 ;
        RECT  5.205 0.770 5.275 1.375 ;
        RECT  4.595 1.145 5.205 1.375 ;
        RECT  4.525 0.770 4.595 1.375 ;
        RECT  3.925 1.145 4.525 1.375 ;
        RECT  3.845 0.770 3.925 1.375 ;
        RECT  3.730 1.145 3.845 1.375 ;
        RECT  3.650 0.675 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.015 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.015 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.015 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 1.015 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 1.015 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.015 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.015 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 1.015 0.510 1.375 ;
        RECT  0.130 1.145 0.390 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.715 3.570 0.945 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.185 0.305 3.475 0.465 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  2.825 0.305 3.115 0.465 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.465 0.305 2.755 0.465 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.205 0.305 2.395 0.465 ;
        RECT  1.675 0.185 1.715 0.465 ;
        RECT  0.210 0.715 1.715 0.945 ;
        RECT  1.385 0.305 1.675 0.465 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.005 0.305 1.315 0.465 ;
        RECT  0.935 0.185 1.005 0.465 ;
        RECT  0.625 0.305 0.935 0.465 ;
        RECT  0.555 0.185 0.625 0.465 ;
        RECT  7.430 0.240 7.510 0.710 ;
        RECT  7.430 0.790 7.510 0.975 ;
        RECT  7.290 0.630 7.430 0.710 ;
        RECT  7.210 0.790 7.430 0.870 ;
        RECT  7.130 0.430 7.210 0.870 ;
        RECT  3.970 0.430 7.130 0.510 ;
        RECT  2.235 0.545 3.565 0.615 ;
    END
END DCCKND20BWP

MACRO DCCKND4BWP
    CLASS CORE ;
    FOREIGN DCCKND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1904 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.215 0.745 0.415 ;
        RECT  0.675 0.700 0.745 1.045 ;
        RECT  0.595 0.305 0.675 0.415 ;
        RECT  0.595 0.700 0.675 0.820 ;
        RECT  0.385 0.305 0.595 0.820 ;
        RECT  0.325 0.305 0.385 0.415 ;
        RECT  0.325 0.700 0.385 0.820 ;
        RECT  0.255 0.215 0.325 0.415 ;
        RECT  0.255 0.700 0.325 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1088 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.530 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.730 -0.115 1.960 0.115 ;
        RECT  1.650 -0.115 1.730 0.350 ;
        RECT  1.125 -0.115 1.650 0.115 ;
        RECT  1.045 -0.115 1.125 0.350 ;
        RECT  0.930 -0.115 1.045 0.115 ;
        RECT  0.850 -0.115 0.930 0.440 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.235 ;
        RECT  0.150 -0.115 0.440 0.115 ;
        RECT  0.070 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.145 1.960 1.375 ;
        RECT  1.610 0.945 1.750 1.375 ;
        RECT  1.125 1.145 1.610 1.375 ;
        RECT  1.045 0.770 1.125 1.375 ;
        RECT  0.930 1.145 1.045 1.375 ;
        RECT  0.850 0.675 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.150 1.145 0.440 1.375 ;
        RECT  0.070 0.750 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.675 0.215 0.745 0.415 ;
        RECT  0.675 0.700 0.745 1.045 ;
        RECT  0.665 0.305 0.675 0.415 ;
        RECT  0.665 0.700 0.675 0.820 ;
        RECT  0.255 0.215 0.315 0.415 ;
        RECT  0.255 0.700 0.315 1.045 ;
        RECT  1.830 0.240 1.910 0.710 ;
        RECT  1.830 0.790 1.910 0.970 ;
        RECT  1.690 0.630 1.830 0.710 ;
        RECT  1.610 0.790 1.830 0.870 ;
        RECT  1.530 0.430 1.610 0.870 ;
        RECT  1.150 0.430 1.530 0.510 ;
    END
END DCCKND4BWP

MACRO DCCKND8BWP
    CLASS CORE ;
    FOREIGN DCCKND8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3928 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.730 1.470 0.960 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.295 0.345 1.375 0.465 ;
        RECT  1.085 0.345 1.295 0.960 ;
        RECT  1.015 0.185 1.085 0.960 ;
        RECT  0.945 0.345 1.015 0.960 ;
        RECT  0.725 0.345 0.945 0.465 ;
        RECT  0.210 0.730 0.945 0.960 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.365 0.345 0.655 0.465 ;
        RECT  0.295 0.185 0.365 0.465 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2176 ;
        ANTENNADIFFAREA 0.0518 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.545 0.845 0.625 ;
        RECT  0.035 0.200 0.140 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 -0.115 3.360 0.115 ;
        RECT  3.040 -0.115 3.120 0.350 ;
        RECT  2.470 -0.115 3.040 0.115 ;
        RECT  2.390 -0.115 2.470 0.350 ;
        RECT  1.825 -0.115 2.390 0.115 ;
        RECT  1.745 -0.115 1.825 0.350 ;
        RECT  1.625 -0.115 1.745 0.115 ;
        RECT  1.555 -0.115 1.625 0.465 ;
        RECT  1.290 -0.115 1.555 0.115 ;
        RECT  1.170 -0.115 1.290 0.275 ;
        RECT  0.930 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.930 0.275 ;
        RECT  0.570 -0.115 0.810 0.115 ;
        RECT  0.450 -0.115 0.570 0.275 ;
        RECT  0.000 -0.115 0.450 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.145 3.360 1.375 ;
        RECT  3.010 0.945 3.150 1.375 ;
        RECT  2.470 1.145 3.010 1.375 ;
        RECT  2.390 0.770 2.470 1.375 ;
        RECT  1.825 1.145 2.390 1.375 ;
        RECT  1.745 0.770 1.825 1.375 ;
        RECT  1.630 1.145 1.745 1.375 ;
        RECT  1.550 0.675 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 1.030 1.280 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.780 1.030 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 1.030 0.520 1.375 ;
        RECT  0.130 1.145 0.400 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.730 1.470 0.960 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.365 0.345 1.375 0.465 ;
        RECT  0.725 0.345 0.875 0.465 ;
        RECT  0.210 0.730 0.875 0.960 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.365 0.345 0.655 0.465 ;
        RECT  0.295 0.185 0.365 0.465 ;
        RECT  3.230 0.230 3.310 0.710 ;
        RECT  3.230 0.790 3.310 0.975 ;
        RECT  3.090 0.630 3.230 0.710 ;
        RECT  3.010 0.790 3.230 0.870 ;
        RECT  2.930 0.430 3.010 0.870 ;
        RECT  1.860 0.430 2.930 0.510 ;
    END
END DCCKND8BWP

MACRO DEL025D1BWP
    CLASS CORE ;
    FOREIGN DEL025D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 0.215 0.665 0.905 ;
        RECT  0.595 0.215 0.615 1.035 ;
        RECT  0.520 0.215 0.595 0.285 ;
        RECT  0.545 0.735 0.595 1.035 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.765 ;
        RECT  0.260 0.495 0.315 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.430 -0.115 0.700 0.115 ;
        RECT  0.310 -0.115 0.430 0.270 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.405 1.145 0.700 1.375 ;
        RECT  0.335 0.845 0.405 1.375 ;
        RECT  0.000 1.145 0.335 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.455 0.355 0.525 0.650 ;
        RECT  0.190 0.355 0.455 0.425 ;
        RECT  0.120 0.185 0.190 1.035 ;
    END
END DEL025D1BWP

MACRO DEL050D1BWP
    CLASS CORE ;
    FOREIGN DEL050D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.195 0.805 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.725 0.525 1.045 ;
        RECT  0.405 0.725 0.455 0.795 ;
        RECT  0.335 0.520 0.405 0.795 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.575 0.210 0.645 0.640 ;
        RECT  0.125 0.210 0.575 0.280 ;
        RECT  0.265 0.365 0.370 0.435 ;
        RECT  0.265 0.875 0.370 0.945 ;
        RECT  0.195 0.365 0.265 0.945 ;
        RECT  0.055 0.210 0.125 0.980 ;
    END
END DEL050D1BWP

MACRO DEL075D1BWP
    CLASS CORE ;
    FOREIGN DEL075D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.085 1.045 ;
        RECT  0.995 0.185 1.015 0.465 ;
        RECT  0.995 0.725 1.015 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.320 ;
        RECT  0.340 -0.115 0.780 0.115 ;
        RECT  0.220 -0.115 0.340 0.285 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.800 0.900 0.880 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 0.945 0.640 ;
        RECT  0.850 0.395 0.920 0.805 ;
        RECT  0.685 0.395 0.850 0.465 ;
        RECT  0.685 0.735 0.850 0.805 ;
        RECT  0.530 0.545 0.780 0.615 ;
        RECT  0.615 0.225 0.685 0.465 ;
        RECT  0.615 0.735 0.685 1.020 ;
        RECT  0.460 0.225 0.530 1.020 ;
        RECT  0.435 0.225 0.460 0.345 ;
        RECT  0.435 0.900 0.460 1.020 ;
        RECT  0.335 0.520 0.390 0.640 ;
        RECT  0.265 0.355 0.335 0.920 ;
        RECT  0.125 0.355 0.265 0.425 ;
        RECT  0.125 0.850 0.265 0.920 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.060 ;
    END
END DEL075D1BWP

MACRO DEL100D1BWP
    CLASS CORE ;
    FOREIGN DEL100D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.045 ;
        RECT  1.275 0.185 1.295 0.465 ;
        RECT  1.275 0.735 1.295 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.130 -0.115 1.400 0.115 ;
        RECT  1.060 -0.115 1.130 0.325 ;
        RECT  0.375 -0.115 1.060 0.115 ;
        RECT  0.255 -0.115 0.375 0.285 ;
        RECT  0.000 -0.115 0.255 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.135 1.145 1.400 1.375 ;
        RECT  1.065 0.835 1.135 1.375 ;
        RECT  0.375 1.145 1.065 1.375 ;
        RECT  0.255 0.975 0.375 1.375 ;
        RECT  0.000 1.145 0.255 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.170 0.520 1.215 0.640 ;
        RECT  1.100 0.395 1.170 0.765 ;
        RECT  0.925 0.395 1.100 0.465 ;
        RECT  0.925 0.695 1.100 0.765 ;
        RECT  0.745 0.545 1.020 0.615 ;
        RECT  0.855 0.195 0.925 0.465 ;
        RECT  0.855 0.695 0.925 1.040 ;
        RECT  0.675 0.195 0.745 1.065 ;
        RECT  0.495 0.195 0.565 1.065 ;
        RECT  0.345 0.355 0.415 0.905 ;
        RECT  0.145 0.355 0.345 0.425 ;
        RECT  0.145 0.835 0.345 0.905 ;
        RECT  0.075 0.195 0.145 0.425 ;
        RECT  0.075 0.835 0.145 1.065 ;
    END
END DEL100D1BWP

MACRO DEL125D1BWP
    CLASS CORE ;
    FOREIGN DEL125D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.045 ;
        RECT  1.415 0.185 1.435 0.465 ;
        RECT  1.415 0.735 1.435 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.115 1.540 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 1.145 1.540 1.375 ;
        RECT  1.205 0.735 1.275 1.375 ;
        RECT  0.335 1.145 1.205 1.375 ;
        RECT  0.265 0.975 0.335 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.300 0.520 1.355 0.640 ;
        RECT  1.230 0.210 1.300 0.640 ;
        RECT  0.920 0.210 1.230 0.280 ;
        RECT  1.000 0.350 1.070 1.070 ;
        RECT  0.850 0.210 0.920 1.070 ;
        RECT  0.820 0.210 0.850 0.460 ;
        RECT  0.815 0.790 0.850 1.070 ;
        RECT  0.705 0.520 0.780 0.640 ;
        RECT  0.635 0.190 0.705 1.070 ;
        RECT  0.460 0.190 0.530 1.070 ;
        RECT  0.320 0.345 0.390 0.905 ;
        RECT  0.145 0.345 0.320 0.415 ;
        RECT  0.145 0.835 0.320 0.905 ;
        RECT  0.075 0.190 0.145 0.415 ;
        RECT  0.075 0.835 0.145 1.070 ;
    END
END DEL125D1BWP

MACRO DEL150D1BWP
    CLASS CORE ;
    FOREIGN DEL150D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.045 ;
        RECT  1.415 0.185 1.435 0.465 ;
        RECT  1.415 0.735 1.435 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0096 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.115 1.540 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 1.145 1.540 1.375 ;
        RECT  1.205 0.735 1.275 1.375 ;
        RECT  0.360 1.145 1.205 1.375 ;
        RECT  0.240 0.975 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.300 0.520 1.355 0.640 ;
        RECT  1.230 0.210 1.300 0.640 ;
        RECT  0.920 0.210 1.230 0.280 ;
        RECT  1.000 0.350 1.070 1.070 ;
        RECT  0.850 0.210 0.920 1.045 ;
        RECT  0.790 0.365 0.850 0.435 ;
        RECT  0.790 0.975 0.850 1.045 ;
        RECT  0.705 0.520 0.780 0.640 ;
        RECT  0.635 0.190 0.705 1.065 ;
        RECT  0.460 0.190 0.530 1.065 ;
        RECT  0.320 0.345 0.390 0.905 ;
        RECT  0.145 0.345 0.320 0.415 ;
        RECT  0.145 0.835 0.320 0.905 ;
        RECT  0.075 0.190 0.145 0.415 ;
        RECT  0.075 0.835 0.145 1.065 ;
    END
END DEL150D1BWP

MACRO DEL175D1BWP
    CLASS CORE ;
    FOREIGN DEL175D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.045 ;
        RECT  1.415 0.185 1.435 0.465 ;
        RECT  1.415 0.735 1.435 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.540 0.115 ;
        RECT  1.220 -0.115 1.300 0.310 ;
        RECT  0.340 -0.115 1.220 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.220 0.820 1.300 1.375 ;
        RECT  0.320 1.145 1.220 1.375 ;
        RECT  0.240 0.975 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.520 1.365 0.640 ;
        RECT  1.260 0.400 1.330 0.750 ;
        RECT  0.895 0.400 1.260 0.470 ;
        RECT  0.895 0.680 1.260 0.750 ;
        RECT  0.710 0.540 1.120 0.610 ;
        RECT  0.825 0.230 0.895 0.470 ;
        RECT  0.825 0.680 0.895 1.030 ;
        RECT  0.640 0.230 0.710 1.005 ;
        RECT  0.445 0.345 0.515 0.905 ;
        RECT  0.125 0.345 0.445 0.415 ;
        RECT  0.125 0.835 0.445 0.905 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.835 0.125 0.995 ;
    END
END DEL175D1BWP

MACRO DEL1D1BWP
    CLASS CORE ;
    FOREIGN DEL1D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.045 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.735 4.655 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 -0.115 4.760 0.115 ;
        RECT  4.450 -0.115 4.530 0.310 ;
        RECT  2.560 -0.115 4.450 0.115 ;
        RECT  2.430 -0.115 2.560 0.455 ;
        RECT  1.470 -0.115 2.430 0.115 ;
        RECT  1.350 -0.115 1.470 0.455 ;
        RECT  0.330 -0.115 1.350 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.145 4.760 1.375 ;
        RECT  4.450 0.820 4.530 1.375 ;
        RECT  2.530 1.145 4.450 1.375 ;
        RECT  2.450 0.830 2.530 1.375 ;
        RECT  1.450 1.145 2.450 1.375 ;
        RECT  1.370 0.805 1.450 1.375 ;
        RECT  0.310 1.145 1.370 1.375 ;
        RECT  0.230 0.835 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.520 4.585 0.640 ;
        RECT  4.235 0.195 4.305 1.065 ;
        RECT  3.820 0.195 4.235 0.265 ;
        RECT  3.605 0.995 4.235 1.065 ;
        RECT  3.985 0.390 4.055 0.920 ;
        RECT  3.425 0.545 3.910 0.615 ;
        RECT  3.740 0.195 3.820 0.455 ;
        RECT  3.510 0.385 3.740 0.455 ;
        RECT  3.535 0.805 3.605 1.065 ;
        RECT  3.355 0.360 3.425 0.990 ;
        RECT  2.900 0.360 2.980 0.990 ;
        RECT  2.350 0.545 2.830 0.615 ;
        RECT  2.270 0.360 2.350 0.965 ;
        RECT  1.825 0.360 1.895 0.965 ;
        RECT  1.265 0.545 1.750 0.615 ;
        RECT  1.195 0.360 1.265 0.990 ;
        RECT  0.400 0.545 0.670 0.615 ;
        RECT  0.330 0.345 0.400 0.765 ;
        RECT  0.125 0.345 0.330 0.415 ;
        RECT  0.125 0.695 0.330 0.765 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  0.055 0.695 0.125 1.035 ;
        RECT  0.745 0.360 0.815 0.990 ;
    END
END DEL1D1BWP

MACRO DEL1P5D1BWP
    CLASS CORE ;
    FOREIGN DEL1P5D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.185 5.145 1.045 ;
        RECT  5.055 0.185 5.075 0.465 ;
        RECT  5.055 0.735 5.075 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.950 -0.115 5.180 0.115 ;
        RECT  4.870 -0.115 4.950 0.310 ;
        RECT  2.770 -0.115 4.870 0.115 ;
        RECT  2.650 -0.115 2.770 0.465 ;
        RECT  1.580 -0.115 2.650 0.115 ;
        RECT  1.450 -0.115 1.580 0.465 ;
        RECT  0.330 -0.115 1.450 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.950 1.145 5.180 1.375 ;
        RECT  4.870 0.820 4.950 1.375 ;
        RECT  2.750 1.145 4.870 1.375 ;
        RECT  2.670 0.790 2.750 1.375 ;
        RECT  1.550 1.145 2.670 1.375 ;
        RECT  1.470 0.790 1.550 1.375 ;
        RECT  0.310 1.145 1.470 1.375 ;
        RECT  0.230 0.835 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.675 0.520 5.005 0.640 ;
        RECT  4.605 0.195 4.675 1.065 ;
        RECT  4.140 0.195 4.605 0.265 ;
        RECT  3.925 0.995 4.605 1.065 ;
        RECT  4.355 0.390 4.425 0.920 ;
        RECT  3.750 0.545 4.275 0.615 ;
        RECT  4.070 0.195 4.140 0.465 ;
        RECT  3.830 0.395 4.070 0.465 ;
        RECT  3.855 0.790 3.925 1.065 ;
        RECT  3.670 0.350 3.750 0.950 ;
        RECT  3.175 0.350 3.245 0.950 ;
        RECT  2.545 0.545 3.095 0.615 ;
        RECT  2.475 0.350 2.545 0.950 ;
        RECT  1.975 0.350 2.045 0.950 ;
        RECT  1.370 0.545 1.895 0.615 ;
        RECT  1.290 0.350 1.370 0.990 ;
        RECT  0.400 0.545 0.715 0.615 ;
        RECT  0.330 0.345 0.400 0.765 ;
        RECT  0.125 0.345 0.330 0.415 ;
        RECT  0.125 0.695 0.330 0.765 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  0.055 0.695 0.125 1.035 ;
        RECT  0.795 0.350 0.865 0.990 ;
    END
END DEL1P5D1BWP

MACRO DEL200D1BWP
    CLASS CORE ;
    FOREIGN DEL200D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.045 ;
        RECT  1.540 0.185 1.575 0.465 ;
        RECT  1.540 0.735 1.575 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.260 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 -0.115 1.680 0.115 ;
        RECT  1.320 -0.115 1.400 0.315 ;
        RECT  0.350 -0.115 1.320 0.115 ;
        RECT  0.230 -0.115 0.350 0.280 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.145 1.680 1.375 ;
        RECT  1.320 0.830 1.400 1.375 ;
        RECT  0.330 1.145 1.320 1.375 ;
        RECT  0.250 0.975 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.455 0.545 1.505 0.615 ;
        RECT  1.385 0.400 1.455 0.760 ;
        RECT  0.945 0.400 1.385 0.470 ;
        RECT  0.945 0.690 1.385 0.760 ;
        RECT  0.765 0.545 1.190 0.615 ;
        RECT  0.875 0.230 0.945 0.470 ;
        RECT  0.875 0.690 0.945 0.870 ;
        RECT  0.695 0.360 0.765 0.830 ;
        RECT  0.430 0.545 0.590 0.615 ;
        RECT  0.360 0.350 0.430 0.905 ;
        RECT  0.145 0.350 0.360 0.420 ;
        RECT  0.145 0.835 0.360 0.905 ;
        RECT  0.075 0.245 0.145 0.420 ;
        RECT  0.075 0.835 0.145 0.995 ;
    END
END DEL200D1BWP

MACRO DEL225D1BWP
    CLASS CORE ;
    FOREIGN DEL225D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.045 ;
        RECT  1.555 0.185 1.575 0.465 ;
        RECT  1.555 0.735 1.575 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 -0.115 1.680 0.115 ;
        RECT  1.360 -0.115 1.440 0.310 ;
        RECT  0.340 -0.115 1.360 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.145 1.680 1.375 ;
        RECT  1.360 0.830 1.440 1.375 ;
        RECT  0.320 1.145 1.360 1.375 ;
        RECT  0.240 0.975 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.470 0.520 1.505 0.640 ;
        RECT  1.400 0.400 1.470 0.760 ;
        RECT  0.965 0.400 1.400 0.470 ;
        RECT  0.965 0.690 1.400 0.760 ;
        RECT  0.790 0.545 1.290 0.615 ;
        RECT  0.895 0.230 0.965 0.470 ;
        RECT  0.895 0.690 0.965 1.030 ;
        RECT  0.720 0.265 0.790 1.005 ;
        RECT  0.410 0.545 0.650 0.615 ;
        RECT  0.340 0.345 0.410 0.905 ;
        RECT  0.125 0.345 0.340 0.415 ;
        RECT  0.125 0.835 0.340 0.905 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.835 0.125 0.995 ;
    END
END DEL225D1BWP

MACRO DEL250D1BWP
    CLASS CORE ;
    FOREIGN DEL250D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.185 1.785 1.045 ;
        RECT  1.695 0.185 1.715 0.465 ;
        RECT  1.695 0.735 1.715 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 -0.115 1.820 0.115 ;
        RECT  1.500 -0.115 1.580 0.310 ;
        RECT  0.340 -0.115 1.500 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 1.145 1.820 1.375 ;
        RECT  1.500 0.830 1.580 1.375 ;
        RECT  0.320 1.145 1.500 1.375 ;
        RECT  0.240 0.835 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.610 0.520 1.645 0.640 ;
        RECT  1.540 0.400 1.610 0.760 ;
        RECT  1.035 0.400 1.540 0.470 ;
        RECT  1.035 0.690 1.540 0.760 ;
        RECT  0.850 0.545 1.390 0.615 ;
        RECT  0.965 0.210 1.035 0.470 ;
        RECT  0.965 0.690 1.035 1.050 ;
        RECT  0.770 0.210 0.850 1.050 ;
        RECT  0.410 0.545 0.690 0.615 ;
        RECT  0.340 0.345 0.410 0.765 ;
        RECT  0.125 0.345 0.340 0.415 ;
        RECT  0.125 0.695 0.340 0.765 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.695 0.125 1.035 ;
    END
END DEL250D1BWP

MACRO DEL2D1BWP
    CLASS CORE ;
    FOREIGN DEL2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.455 0.185 7.525 1.045 ;
        RECT  7.435 0.185 7.455 0.465 ;
        RECT  7.435 0.735 7.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.330 -0.115 7.560 0.115 ;
        RECT  7.250 -0.115 7.330 0.310 ;
        RECT  5.150 -0.115 7.250 0.115 ;
        RECT  5.030 -0.115 5.150 0.465 ;
        RECT  3.960 -0.115 5.030 0.115 ;
        RECT  3.830 -0.115 3.960 0.465 ;
        RECT  2.770 -0.115 3.830 0.115 ;
        RECT  2.650 -0.115 2.770 0.465 ;
        RECT  1.580 -0.115 2.650 0.115 ;
        RECT  1.450 -0.115 1.580 0.465 ;
        RECT  0.330 -0.115 1.450 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.330 1.145 7.560 1.375 ;
        RECT  7.250 0.835 7.330 1.375 ;
        RECT  5.130 1.145 7.250 1.375 ;
        RECT  5.050 0.790 5.130 1.375 ;
        RECT  3.930 1.145 5.050 1.375 ;
        RECT  3.850 0.790 3.930 1.375 ;
        RECT  2.750 1.145 3.850 1.375 ;
        RECT  2.670 0.790 2.750 1.375 ;
        RECT  1.550 1.145 2.670 1.375 ;
        RECT  1.470 0.790 1.550 1.375 ;
        RECT  0.310 1.145 1.470 1.375 ;
        RECT  0.230 0.835 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.055 0.520 7.385 0.640 ;
        RECT  6.985 0.195 7.055 1.065 ;
        RECT  6.520 0.195 6.985 0.265 ;
        RECT  6.305 0.995 6.985 1.065 ;
        RECT  6.735 0.390 6.805 0.920 ;
        RECT  6.130 0.545 6.655 0.615 ;
        RECT  6.450 0.195 6.520 0.465 ;
        RECT  6.210 0.395 6.450 0.465 ;
        RECT  6.235 0.830 6.305 1.065 ;
        RECT  6.050 0.350 6.130 0.950 ;
        RECT  5.555 0.350 5.625 0.950 ;
        RECT  4.925 0.545 5.475 0.615 ;
        RECT  4.855 0.350 4.925 0.950 ;
        RECT  4.355 0.350 4.425 0.950 ;
        RECT  3.750 0.545 4.275 0.615 ;
        RECT  3.670 0.350 3.750 0.950 ;
        RECT  3.175 0.350 3.245 0.950 ;
        RECT  2.545 0.545 3.095 0.615 ;
        RECT  2.475 0.350 2.545 0.950 ;
        RECT  1.975 0.350 2.045 0.950 ;
        RECT  1.370 0.545 1.895 0.615 ;
        RECT  1.290 0.350 1.370 0.990 ;
        RECT  0.795 0.350 0.865 0.990 ;
        RECT  0.400 0.545 0.715 0.615 ;
        RECT  0.330 0.345 0.400 0.765 ;
        RECT  0.125 0.345 0.330 0.415 ;
        RECT  0.125 0.695 0.330 0.765 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  0.055 0.695 0.125 1.035 ;
    END
END DEL2D1BWP

MACRO DEL500D1BWP
    CLASS CORE ;
    FOREIGN DEL500D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.625 1.045 ;
        RECT  2.535 0.185 2.555 0.465 ;
        RECT  2.535 0.735 2.555 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.115 2.660 0.115 ;
        RECT  2.350 -0.115 2.430 0.310 ;
        RECT  0.330 -0.115 2.350 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.145 2.660 1.375 ;
        RECT  2.350 0.835 2.430 1.375 ;
        RECT  0.310 1.145 2.350 1.375 ;
        RECT  0.230 0.835 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.520 2.485 0.640 ;
        RECT  2.135 0.195 2.205 1.065 ;
        RECT  1.680 0.195 2.135 0.265 ;
        RECT  1.465 0.995 2.135 1.065 ;
        RECT  1.845 0.390 1.915 0.920 ;
        RECT  1.265 0.545 1.770 0.615 ;
        RECT  1.610 0.195 1.680 0.455 ;
        RECT  1.370 0.385 1.610 0.455 ;
        RECT  1.395 0.805 1.465 1.065 ;
        RECT  1.195 0.370 1.265 0.990 ;
        RECT  0.745 0.370 0.815 0.990 ;
        RECT  0.400 0.545 0.670 0.615 ;
        RECT  0.330 0.345 0.400 0.765 ;
        RECT  0.125 0.345 0.330 0.415 ;
        RECT  0.125 0.695 0.330 0.765 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  0.055 0.695 0.125 1.035 ;
    END
END DEL500D1BWP

MACRO DFCND1BWP
    CLASS CORE ;
    FOREIGN DFCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.045 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.520 0.730 3.535 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.415 3.310 0.785 ;
        RECT  3.205 0.415 3.240 0.485 ;
        RECT  3.110 0.715 3.240 0.785 ;
        RECT  3.115 0.205 3.205 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.630 ;
        RECT  2.645 0.510 2.695 0.630 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 -0.115 3.640 0.115 ;
        RECT  3.320 -0.115 3.400 0.335 ;
        RECT  2.615 -0.115 3.320 0.115 ;
        RECT  2.545 -0.115 2.615 0.360 ;
        RECT  1.570 -0.115 2.545 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.360 -0.115 0.595 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.145 3.640 1.375 ;
        RECT  3.300 1.010 3.420 1.375 ;
        RECT  0.000 1.145 3.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.450 0.520 3.460 0.640 ;
        RECT  3.380 0.520 3.450 0.935 ;
        RECT  2.910 0.865 3.380 0.935 ;
        RECT  3.005 0.555 3.150 0.625 ;
        RECT  2.935 0.230 3.005 0.775 ;
        RECT  2.510 0.705 2.935 0.775 ;
        RECT  2.840 0.845 2.910 0.935 ;
        RECT  2.770 1.005 2.880 1.075 ;
        RECT  2.370 0.845 2.840 0.915 ;
        RECT  2.700 0.985 2.770 1.075 ;
        RECT  2.230 0.985 2.700 1.055 ;
        RECT  2.440 0.520 2.510 0.775 ;
        RECT  2.410 0.520 2.440 0.640 ;
        RECT  2.340 0.380 2.430 0.450 ;
        RECT  2.340 0.700 2.370 0.915 ;
        RECT  2.300 0.380 2.340 0.915 ;
        RECT  1.710 0.200 2.330 0.270 ;
        RECT  2.270 0.380 2.300 0.770 ;
        RECT  2.130 0.380 2.270 0.450 ;
        RECT  2.175 0.830 2.230 1.055 ;
        RECT  2.160 0.660 2.175 1.055 ;
        RECT  2.105 0.660 2.160 0.900 ;
        RECT  2.045 0.660 2.105 0.730 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.350 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.535 1.700 0.605 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.845 1.590 0.915 ;
        RECT  1.390 0.500 1.460 0.605 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.330 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCND1BWP

MACRO DFCND2BWP
    CLASS CORE ;
    FOREIGN DFCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.355 4.025 0.800 ;
        RECT  3.955 0.185 3.965 1.035 ;
        RECT  3.895 0.185 3.955 0.465 ;
        RECT  3.895 0.730 3.955 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 0.785 ;
        RECT  3.475 0.185 3.535 0.465 ;
        RECT  3.440 0.715 3.535 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0524 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.640 ;
        RECT  2.595 0.510 2.695 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.300 ;
        RECT  3.755 -0.115 4.070 0.115 ;
        RECT  3.685 -0.115 3.755 0.465 ;
        RECT  3.365 -0.115 3.685 0.115 ;
        RECT  3.295 -0.115 3.365 0.420 ;
        RECT  2.605 -0.115 3.295 0.115 ;
        RECT  2.535 -0.115 2.605 0.430 ;
        RECT  1.570 -0.115 2.535 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.360 -0.115 0.595 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.145 4.200 1.375 ;
        RECT  4.060 0.870 4.160 1.375 ;
        RECT  3.780 1.145 4.060 1.375 ;
        RECT  3.660 1.030 3.780 1.375 ;
        RECT  3.380 1.145 3.660 1.375 ;
        RECT  3.260 1.030 3.380 1.375 ;
        RECT  0.000 1.145 3.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.780 0.545 3.880 0.615 ;
        RECT  3.710 0.545 3.780 0.925 ;
        RECT  2.370 0.855 3.710 0.925 ;
        RECT  3.200 0.545 3.460 0.615 ;
        RECT  3.130 0.325 3.200 0.785 ;
        RECT  2.890 0.325 3.130 0.395 ;
        RECT  2.510 0.715 3.130 0.785 ;
        RECT  2.720 0.995 2.840 1.075 ;
        RECT  2.230 0.995 2.720 1.065 ;
        RECT  2.440 0.520 2.510 0.785 ;
        RECT  2.340 0.375 2.450 0.445 ;
        RECT  2.410 0.520 2.440 0.640 ;
        RECT  2.340 0.700 2.370 0.925 ;
        RECT  1.710 0.200 2.350 0.270 ;
        RECT  2.300 0.375 2.340 0.925 ;
        RECT  2.270 0.375 2.300 0.770 ;
        RECT  2.130 0.375 2.270 0.445 ;
        RECT  2.175 0.830 2.230 1.065 ;
        RECT  2.160 0.660 2.175 1.065 ;
        RECT  2.105 0.660 2.160 0.900 ;
        RECT  2.045 0.660 2.105 0.730 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.350 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.330 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCND2BWP

MACRO DFCND4BWP
    CLASS CORE ;
    FOREIGN DFCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.665 0.485 ;
        RECT  4.655 0.765 4.665 1.065 ;
        RECT  4.595 0.185 4.655 1.065 ;
        RECT  4.445 0.355 4.595 0.905 ;
        RECT  4.310 0.355 4.445 0.485 ;
        RECT  4.305 0.765 4.445 0.905 ;
        RECT  4.240 0.185 4.310 0.485 ;
        RECT  4.235 0.765 4.305 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.705 3.960 0.785 ;
        RECT  3.855 0.185 3.925 0.475 ;
        RECT  3.815 0.355 3.855 0.475 ;
        RECT  3.605 0.355 3.815 0.785 ;
        RECT  3.545 0.355 3.605 0.475 ;
        RECT  3.440 0.705 3.605 0.785 ;
        RECT  3.475 0.185 3.545 0.475 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.640 ;
        RECT  2.595 0.510 2.695 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.115 4.900 0.115 ;
        RECT  4.770 -0.115 4.850 0.465 ;
        RECT  4.510 -0.115 4.770 0.115 ;
        RECT  4.390 -0.115 4.510 0.275 ;
        RECT  4.115 -0.115 4.390 0.115 ;
        RECT  4.045 -0.115 4.115 0.465 ;
        RECT  3.760 -0.115 4.045 0.115 ;
        RECT  3.640 -0.115 3.760 0.275 ;
        RECT  3.365 -0.115 3.640 0.115 ;
        RECT  3.295 -0.115 3.365 0.445 ;
        RECT  2.605 -0.115 3.295 0.115 ;
        RECT  2.535 -0.115 2.605 0.430 ;
        RECT  1.570 -0.115 2.535 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.145 4.900 1.375 ;
        RECT  4.770 0.680 4.850 1.375 ;
        RECT  4.485 1.145 4.770 1.375 ;
        RECT  4.415 0.975 4.485 1.375 ;
        RECT  4.140 1.145 4.415 1.375 ;
        RECT  4.020 1.010 4.140 1.375 ;
        RECT  3.760 1.145 4.020 1.375 ;
        RECT  3.640 1.010 3.760 1.375 ;
        RECT  3.380 1.145 3.640 1.375 ;
        RECT  3.260 1.010 3.380 1.375 ;
        RECT  0.690 1.145 3.260 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.310 0.355 4.375 0.485 ;
        RECT  4.305 0.765 4.375 0.905 ;
        RECT  4.240 0.185 4.310 0.485 ;
        RECT  4.235 0.765 4.305 1.065 ;
        RECT  3.885 0.705 3.960 0.785 ;
        RECT  3.885 0.185 3.925 0.475 ;
        RECT  3.475 0.185 3.535 0.475 ;
        RECT  3.440 0.705 3.535 0.785 ;
        RECT  4.130 0.545 4.200 0.615 ;
        RECT  4.060 0.545 4.130 0.925 ;
        RECT  2.370 0.855 4.060 0.925 ;
        RECT  3.200 0.545 3.470 0.615 ;
        RECT  3.130 0.325 3.200 0.785 ;
        RECT  2.890 0.325 3.130 0.395 ;
        RECT  2.510 0.715 3.130 0.785 ;
        RECT  2.720 0.995 2.840 1.075 ;
        RECT  2.230 0.995 2.720 1.065 ;
        RECT  2.440 0.520 2.510 0.785 ;
        RECT  2.340 0.375 2.450 0.445 ;
        RECT  2.410 0.520 2.440 0.640 ;
        RECT  2.340 0.700 2.370 0.925 ;
        RECT  1.710 0.200 2.350 0.270 ;
        RECT  2.300 0.375 2.340 0.925 ;
        RECT  2.270 0.375 2.300 0.770 ;
        RECT  2.130 0.375 2.270 0.445 ;
        RECT  2.175 0.830 2.230 1.065 ;
        RECT  2.160 0.660 2.175 1.065 ;
        RECT  2.105 0.660 2.160 0.900 ;
        RECT  2.045 0.660 2.105 0.730 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.350 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.860 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.790 0.870 0.860 1.055 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.330 0.870 0.790 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.465 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.465 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFCND4BWP

MACRO DFCNQD1BWP
    CLASS CORE ;
    FOREIGN DFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.185 1.045 ;
        RECT  3.095 0.185 3.115 0.465 ;
        RECT  3.095 0.735 3.115 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.545 2.700 0.625 ;
        RECT  2.555 0.355 2.625 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.980 0.290 ;
        RECT  2.405 -0.115 2.900 0.115 ;
        RECT  2.335 -0.115 2.405 0.450 ;
        RECT  1.570 -0.115 2.335 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 1.145 3.220 1.375 ;
        RECT  2.880 1.010 3.000 1.375 ;
        RECT  0.000 1.145 2.880 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.025 0.520 3.040 0.640 ;
        RECT  2.955 0.370 3.025 0.930 ;
        RECT  2.775 0.370 2.955 0.440 ;
        RECT  2.710 0.860 2.955 0.930 ;
        RECT  2.785 0.520 2.855 0.790 ;
        RECT  2.560 0.720 2.785 0.790 ;
        RECT  2.705 0.205 2.775 0.440 ;
        RECT  2.640 0.860 2.710 1.060 ;
        RECT  2.510 0.205 2.705 0.275 ;
        RECT  2.460 0.990 2.640 1.060 ;
        RECT  2.490 0.720 2.560 0.910 ;
        RECT  2.150 0.840 2.490 0.910 ;
        RECT  2.340 0.990 2.460 1.070 ;
        RECT  2.230 0.520 2.300 0.770 ;
        RECT  2.210 0.520 2.230 0.590 ;
        RECT  2.140 0.200 2.210 0.590 ;
        RECT  2.080 0.660 2.150 0.910 ;
        RECT  1.710 0.200 2.140 0.270 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  2.045 0.660 2.080 0.730 ;
        RECT  1.975 0.340 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.530 1.700 0.600 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.840 1.590 0.910 ;
        RECT  1.390 0.500 1.460 0.600 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.330 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCNQD1BWP

MACRO DFCNQD2BWP
    CLASS CORE ;
    FOREIGN DFCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.545 0.355 3.605 0.815 ;
        RECT  3.535 0.185 3.545 1.035 ;
        RECT  3.475 0.185 3.535 0.465 ;
        RECT  3.475 0.745 3.535 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.495 3.045 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.300 ;
        RECT  3.370 -0.115 3.650 0.115 ;
        RECT  3.300 -0.115 3.370 0.465 ;
        RECT  2.585 -0.115 3.300 0.115 ;
        RECT  2.515 -0.115 2.585 0.440 ;
        RECT  2.405 -0.115 2.515 0.115 ;
        RECT  2.335 -0.115 2.405 0.445 ;
        RECT  1.570 -0.115 2.335 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.895 3.730 1.375 ;
        RECT  3.380 1.145 3.650 1.375 ;
        RECT  3.260 1.010 3.380 1.375 ;
        RECT  3.000 1.145 3.260 1.375 ;
        RECT  2.880 1.010 3.000 1.375 ;
        RECT  0.000 1.145 2.880 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.405 0.545 3.460 0.615 ;
        RECT  3.335 0.545 3.405 0.940 ;
        RECT  2.870 0.870 3.335 0.940 ;
        RECT  3.160 0.205 3.230 0.660 ;
        RECT  2.730 0.205 3.160 0.275 ;
        RECT  2.870 0.345 2.995 0.415 ;
        RECT  2.800 0.345 2.870 0.940 ;
        RECT  2.640 0.870 2.800 0.940 ;
        RECT  2.675 0.205 2.730 0.640 ;
        RECT  2.660 0.205 2.675 0.800 ;
        RECT  2.605 0.520 2.660 0.800 ;
        RECT  2.570 0.870 2.640 1.050 ;
        RECT  2.470 0.730 2.605 0.800 ;
        RECT  2.460 0.980 2.570 1.050 ;
        RECT  2.400 0.730 2.470 0.910 ;
        RECT  2.340 0.980 2.460 1.060 ;
        RECT  2.160 0.840 2.400 0.910 ;
        RECT  2.230 0.530 2.320 0.760 ;
        RECT  2.220 0.530 2.230 0.600 ;
        RECT  2.150 0.200 2.220 0.600 ;
        RECT  2.090 0.695 2.160 0.910 ;
        RECT  1.710 0.200 2.150 0.270 ;
        RECT  2.045 0.695 2.090 0.765 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.340 2.045 0.765 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.330 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCNQD2BWP

MACRO DFCNQD4BWP
    CLASS CORE ;
    FOREIGN DFCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.465 ;
        RECT  3.955 0.765 3.965 1.065 ;
        RECT  3.895 0.185 3.955 1.065 ;
        RECT  3.745 0.355 3.895 0.905 ;
        RECT  3.585 0.355 3.745 0.465 ;
        RECT  3.585 0.765 3.745 0.905 ;
        RECT  3.515 0.185 3.585 0.465 ;
        RECT  3.515 0.765 3.585 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.495 3.045 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.475 ;
        RECT  3.800 -0.115 4.070 0.115 ;
        RECT  3.680 -0.115 3.800 0.275 ;
        RECT  3.410 -0.115 3.680 0.115 ;
        RECT  3.340 -0.115 3.410 0.465 ;
        RECT  2.585 -0.115 3.340 0.115 ;
        RECT  2.515 -0.115 2.585 0.440 ;
        RECT  2.405 -0.115 2.515 0.115 ;
        RECT  2.335 -0.115 2.405 0.445 ;
        RECT  1.570 -0.115 2.335 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.675 4.150 1.375 ;
        RECT  3.775 1.145 4.070 1.375 ;
        RECT  3.705 0.975 3.775 1.375 ;
        RECT  3.420 1.145 3.705 1.375 ;
        RECT  3.300 1.010 3.420 1.375 ;
        RECT  3.020 1.145 3.300 1.375 ;
        RECT  2.900 1.010 3.020 1.375 ;
        RECT  0.690 1.145 2.900 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.585 0.355 3.675 0.465 ;
        RECT  3.585 0.765 3.675 0.905 ;
        RECT  3.515 0.185 3.585 0.465 ;
        RECT  3.515 0.765 3.585 1.065 ;
        RECT  3.425 0.545 3.550 0.615 ;
        RECT  3.355 0.545 3.425 0.940 ;
        RECT  2.870 0.870 3.355 0.940 ;
        RECT  3.200 0.205 3.270 0.660 ;
        RECT  2.730 0.205 3.200 0.275 ;
        RECT  2.870 0.345 3.010 0.415 ;
        RECT  2.800 0.345 2.870 0.940 ;
        RECT  2.640 0.870 2.800 0.940 ;
        RECT  2.675 0.205 2.730 0.640 ;
        RECT  2.660 0.205 2.675 0.800 ;
        RECT  2.605 0.520 2.660 0.800 ;
        RECT  2.570 0.870 2.640 1.050 ;
        RECT  2.470 0.730 2.605 0.800 ;
        RECT  2.460 0.980 2.570 1.050 ;
        RECT  2.400 0.730 2.470 0.910 ;
        RECT  2.340 0.980 2.460 1.060 ;
        RECT  2.160 0.840 2.400 0.910 ;
        RECT  2.230 0.530 2.320 0.760 ;
        RECT  2.220 0.530 2.230 0.600 ;
        RECT  2.150 0.200 2.220 0.600 ;
        RECT  2.090 0.695 2.160 0.910 ;
        RECT  1.710 0.200 2.150 0.270 ;
        RECT  2.045 0.695 2.090 0.765 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.340 2.045 0.765 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.830 0.205 1.040 0.275 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.860 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.790 0.870 0.860 1.055 ;
        RECT  0.760 0.205 0.830 0.410 ;
        RECT  0.330 0.870 0.790 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.465 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.465 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFCNQD4BWP

MACRO DFCSND1BWP
    CLASS CORE ;
    FOREIGN DFCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.795 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.740 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0779 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.720 0.775 3.750 1.045 ;
        RECT  3.675 0.350 3.720 1.045 ;
        RECT  3.650 0.350 3.675 0.915 ;
        RECT  3.560 0.350 3.650 0.470 ;
        RECT  3.560 0.775 3.650 0.915 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.495 3.185 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.115 4.060 0.115 ;
        RECT  2.990 -0.115 3.110 0.275 ;
        RECT  1.620 -0.115 2.990 0.115 ;
        RECT  1.500 -0.115 1.620 0.210 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 4.060 1.375 ;
        RECT  2.600 1.030 2.720 1.375 ;
        RECT  2.010 1.145 2.600 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.010 1.650 1.375 ;
        RECT  0.000 1.145 1.530 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.880 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.260 0.210 3.790 0.280 ;
        RECT  3.480 0.545 3.570 0.615 ;
        RECT  3.410 0.355 3.480 1.045 ;
        RECT  3.340 0.355 3.410 0.425 ;
        RECT  2.860 0.975 3.410 1.045 ;
        RECT  3.270 0.520 3.340 0.905 ;
        RECT  2.345 0.835 3.270 0.905 ;
        RECT  3.190 0.210 3.260 0.425 ;
        RECT  2.485 0.355 3.190 0.425 ;
        RECT  2.485 0.695 2.910 0.765 ;
        RECT  1.790 0.200 2.490 0.270 ;
        RECT  2.415 0.355 2.485 0.765 ;
        RECT  2.250 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.905 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.850 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.580 0.850 2.120 0.920 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.200 1.790 0.350 ;
        RECT  1.670 0.420 1.760 0.640 ;
        RECT  1.380 0.280 1.720 0.350 ;
        RECT  1.080 0.420 1.670 0.490 ;
        RECT  1.530 0.560 1.600 0.780 ;
        RECT  1.530 0.850 1.580 0.940 ;
        RECT  1.220 0.560 1.530 0.630 ;
        RECT  1.360 0.870 1.530 0.940 ;
        RECT  1.360 0.700 1.460 0.800 ;
        RECT  1.310 0.195 1.380 0.350 ;
        RECT  1.220 0.730 1.360 0.800 ;
        RECT  1.290 0.870 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.330 0.980 1.290 1.050 ;
        RECT  1.150 0.730 1.220 0.900 ;
        RECT  1.010 0.340 1.080 0.885 ;
        RECT  0.930 0.340 1.010 0.420 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCSND1BWP

MACRO DFCSND2BWP
    CLASS CORE ;
    FOREIGN DFCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.790 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.385 0.355 4.445 0.810 ;
        RECT  4.375 0.185 4.385 1.040 ;
        RECT  4.315 0.185 4.375 0.465 ;
        RECT  4.315 0.740 4.375 1.040 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.355 4.025 1.045 ;
        RECT  3.920 0.355 3.955 0.455 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0584 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.690 0.640 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.300 ;
        RECT  3.040 -0.115 4.490 0.115 ;
        RECT  2.970 -0.115 3.040 0.270 ;
        RECT  1.620 -0.115 2.970 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.895 4.570 1.375 ;
        RECT  4.195 1.145 4.490 1.375 ;
        RECT  4.125 0.735 4.195 1.375 ;
        RECT  3.840 1.145 4.125 1.375 ;
        RECT  3.720 1.005 3.840 1.375 ;
        RECT  3.470 1.145 3.720 1.375 ;
        RECT  3.350 1.005 3.470 1.375 ;
        RECT  3.100 1.145 3.350 1.375 ;
        RECT  2.980 1.005 3.100 1.375 ;
        RECT  2.730 1.145 2.980 1.375 ;
        RECT  2.610 0.985 2.730 1.375 ;
        RECT  2.010 1.145 2.610 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.700 1.145 1.890 1.375 ;
        RECT  1.620 1.005 1.700 1.375 ;
        RECT  1.530 1.005 1.620 1.075 ;
        RECT  0.000 1.145 1.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.210 0.545 4.300 0.615 ;
        RECT  4.140 0.215 4.210 0.615 ;
        RECT  3.185 0.215 4.140 0.285 ;
        RECT  3.830 0.520 3.880 0.640 ;
        RECT  3.760 0.355 3.830 0.935 ;
        RECT  3.325 0.355 3.760 0.425 ;
        RECT  3.170 0.865 3.760 0.935 ;
        RECT  3.395 0.520 3.465 0.785 ;
        RECT  3.080 0.715 3.395 0.785 ;
        RECT  3.255 0.355 3.325 0.615 ;
        RECT  2.860 0.545 3.255 0.615 ;
        RECT  3.115 0.215 3.185 0.425 ;
        RECT  2.485 0.355 3.115 0.425 ;
        RECT  3.010 0.715 3.080 0.915 ;
        RECT  2.345 0.845 3.010 0.915 ;
        RECT  2.485 0.705 2.910 0.775 ;
        RECT  2.415 0.355 2.485 0.775 ;
        RECT  1.790 0.200 2.450 0.270 ;
        RECT  2.250 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.915 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.850 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.555 0.850 2.120 0.920 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.510 0.850 1.555 0.935 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.865 1.510 0.935 ;
        RECT  1.360 0.690 1.460 0.795 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.725 1.360 0.795 ;
        RECT  1.290 0.865 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.330 0.980 1.290 1.050 ;
        RECT  1.150 0.725 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCSND2BWP

MACRO DFCSND4BWP
    CLASS CORE ;
    FOREIGN DFCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.790 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.185 5.085 0.485 ;
        RECT  5.075 0.765 5.085 1.065 ;
        RECT  5.015 0.185 5.075 1.065 ;
        RECT  4.865 0.355 5.015 0.905 ;
        RECT  4.730 0.355 4.865 0.485 ;
        RECT  4.725 0.765 4.865 0.905 ;
        RECT  4.660 0.185 4.730 0.485 ;
        RECT  4.655 0.765 4.725 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.350 4.370 0.485 ;
        RECT  4.275 0.765 4.345 1.065 ;
        RECT  4.235 0.765 4.275 0.905 ;
        RECT  4.025 0.350 4.235 0.905 ;
        RECT  3.900 0.350 4.025 0.470 ;
        RECT  4.005 0.765 4.025 0.905 ;
        RECT  3.915 0.765 4.005 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0584 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.690 0.640 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.905 -0.115 5.190 0.115 ;
        RECT  4.835 -0.115 4.905 0.280 ;
        RECT  3.030 -0.115 4.835 0.115 ;
        RECT  2.960 -0.115 3.030 0.270 ;
        RECT  1.620 -0.115 2.960 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.675 5.270 1.375 ;
        RECT  4.905 1.145 5.190 1.375 ;
        RECT  4.835 0.975 4.905 1.375 ;
        RECT  4.535 1.145 4.835 1.375 ;
        RECT  4.465 0.745 4.535 1.375 ;
        RECT  4.170 1.145 4.465 1.375 ;
        RECT  4.090 0.975 4.170 1.375 ;
        RECT  3.830 1.145 4.090 1.375 ;
        RECT  3.710 1.005 3.830 1.375 ;
        RECT  3.470 1.145 3.710 1.375 ;
        RECT  3.350 1.005 3.470 1.375 ;
        RECT  3.100 1.145 3.350 1.375 ;
        RECT  2.980 1.005 3.100 1.375 ;
        RECT  2.730 1.145 2.980 1.375 ;
        RECT  2.610 0.985 2.730 1.375 ;
        RECT  2.010 1.145 2.610 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.000 1.650 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.355 4.795 0.485 ;
        RECT  4.725 0.765 4.795 0.905 ;
        RECT  4.660 0.185 4.730 0.485 ;
        RECT  4.655 0.765 4.725 1.065 ;
        RECT  4.305 0.350 4.370 0.485 ;
        RECT  4.305 0.765 4.345 1.065 ;
        RECT  3.900 0.350 3.955 0.470 ;
        RECT  3.915 0.765 3.955 1.065 ;
        RECT  4.550 0.545 4.620 0.615 ;
        RECT  4.480 0.210 4.550 0.615 ;
        RECT  3.185 0.210 4.480 0.280 ;
        RECT  3.830 0.545 3.930 0.615 ;
        RECT  3.760 0.355 3.830 0.935 ;
        RECT  3.325 0.355 3.760 0.425 ;
        RECT  3.170 0.865 3.760 0.935 ;
        RECT  3.395 0.520 3.465 0.785 ;
        RECT  3.080 0.715 3.395 0.785 ;
        RECT  3.255 0.355 3.325 0.615 ;
        RECT  2.860 0.545 3.255 0.615 ;
        RECT  3.115 0.210 3.185 0.425 ;
        RECT  2.485 0.355 3.115 0.425 ;
        RECT  3.010 0.715 3.080 0.915 ;
        RECT  2.345 0.845 3.010 0.915 ;
        RECT  2.485 0.705 2.910 0.775 ;
        RECT  1.790 0.205 2.500 0.275 ;
        RECT  2.415 0.355 2.485 0.775 ;
        RECT  2.250 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.915 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.850 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.565 0.850 2.120 0.920 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.205 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.510 0.850 1.565 0.930 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.860 1.510 0.930 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.860 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.790 0.870 0.860 1.050 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.330 0.870 0.790 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.475 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.475 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFCSND4BWP

MACRO DFCSNQD1BWP
    CLASS CORE ;
    FOREIGN DFCSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.625 ;
        RECT  2.690 0.545 2.835 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.195 3.885 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.495 3.185 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.685 -0.115 3.920 0.115 ;
        RECT  3.615 -0.115 3.685 0.465 ;
        RECT  3.120 -0.115 3.615 0.115 ;
        RECT  3.035 -0.115 3.120 0.315 ;
        RECT  1.620 -0.115 3.035 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.685 1.145 3.920 1.375 ;
        RECT  3.615 0.735 3.685 1.375 ;
        RECT  2.750 1.145 3.615 1.375 ;
        RECT  2.630 1.030 2.750 1.375 ;
        RECT  2.030 1.145 2.630 1.375 ;
        RECT  1.910 1.000 2.030 1.375 ;
        RECT  1.670 1.145 1.910 1.375 ;
        RECT  1.550 1.000 1.670 1.375 ;
        RECT  0.000 1.145 1.550 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.500 0.545 3.720 0.615 ;
        RECT  3.465 0.395 3.500 1.045 ;
        RECT  3.430 0.185 3.465 1.045 ;
        RECT  3.395 0.185 3.430 0.465 ;
        RECT  2.880 0.975 3.430 1.045 ;
        RECT  3.280 0.520 3.350 0.905 ;
        RECT  2.365 0.835 3.280 0.905 ;
        RECT  2.505 0.695 2.930 0.765 ;
        RECT  2.505 0.375 2.705 0.455 ;
        RECT  1.790 0.200 2.510 0.270 ;
        RECT  2.435 0.375 2.505 0.765 ;
        RECT  2.270 0.375 2.435 0.455 ;
        RECT  2.295 0.570 2.365 0.905 ;
        RECT  2.185 0.570 2.295 0.640 ;
        RECT  2.005 0.710 2.210 0.780 ;
        RECT  2.140 0.860 2.210 1.075 ;
        RECT  2.115 0.350 2.185 0.640 ;
        RECT  1.360 0.860 2.140 0.930 ;
        RECT  1.935 0.350 2.005 0.780 ;
        RECT  1.600 0.710 1.935 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.330 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCSNQD1BWP

MACRO DFCSNQD2BWP
    CLASS CORE ;
    FOREIGN DFCSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0396 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.215 2.905 0.620 ;
        RECT  2.590 0.550 2.835 0.620 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.355 4.025 0.805 ;
        RECT  3.955 0.185 3.965 1.035 ;
        RECT  3.895 0.185 3.955 0.465 ;
        RECT  3.895 0.735 3.955 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.520 3.675 0.640 ;
        RECT  3.535 0.355 3.605 0.640 ;
        RECT  3.185 0.355 3.535 0.425 ;
        RECT  3.115 0.355 3.185 0.640 ;
        RECT  3.075 0.495 3.115 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.300 ;
        RECT  3.045 -0.115 4.070 0.115 ;
        RECT  2.975 -0.115 3.045 0.410 ;
        RECT  1.620 -0.115 2.975 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.895 4.150 1.375 ;
        RECT  3.785 1.145 4.070 1.375 ;
        RECT  3.715 0.895 3.785 1.375 ;
        RECT  3.425 1.145 3.715 1.375 ;
        RECT  3.355 0.990 3.425 1.375 ;
        RECT  2.720 1.145 3.355 1.375 ;
        RECT  2.600 1.040 2.720 1.375 ;
        RECT  2.010 1.145 2.600 1.375 ;
        RECT  1.890 1.005 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.005 1.650 1.375 ;
        RECT  0.000 1.145 1.530 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.815 0.545 3.880 0.615 ;
        RECT  3.745 0.215 3.815 0.805 ;
        RECT  3.310 0.215 3.745 0.285 ;
        RECT  3.605 0.735 3.745 0.805 ;
        RECT  3.535 0.735 3.605 1.035 ;
        RECT  3.245 0.850 3.535 0.920 ;
        RECT  3.345 0.520 3.415 0.780 ;
        RECT  3.095 0.710 3.345 0.780 ;
        RECT  3.175 0.850 3.245 1.040 ;
        RECT  2.860 0.970 3.175 1.040 ;
        RECT  3.025 0.710 3.095 0.900 ;
        RECT  2.345 0.830 3.025 0.900 ;
        RECT  2.485 0.690 2.910 0.760 ;
        RECT  2.485 0.355 2.660 0.425 ;
        RECT  1.790 0.200 2.490 0.270 ;
        RECT  2.415 0.355 2.485 0.760 ;
        RECT  2.270 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.900 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.865 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.360 0.865 2.120 0.935 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.865 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.330 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFCSNQD2BWP

MACRO DFCSNQD4BWP
    CLASS CORE ;
    FOREIGN DFCSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.625 ;
        RECT  2.690 0.545 2.835 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.185 4.385 0.485 ;
        RECT  4.375 0.735 4.385 1.065 ;
        RECT  4.315 0.185 4.375 1.065 ;
        RECT  4.165 0.355 4.315 0.905 ;
        RECT  4.030 0.355 4.165 0.485 ;
        RECT  4.025 0.735 4.165 0.905 ;
        RECT  3.960 0.185 4.030 0.485 ;
        RECT  3.955 0.735 4.025 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.520 3.715 0.640 ;
        RECT  3.535 0.355 3.605 0.640 ;
        RECT  3.185 0.355 3.535 0.425 ;
        RECT  3.115 0.355 3.185 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.465 ;
        RECT  4.230 -0.115 4.490 0.115 ;
        RECT  4.110 -0.115 4.230 0.275 ;
        RECT  3.130 -0.115 4.110 0.115 ;
        RECT  3.010 -0.115 3.130 0.275 ;
        RECT  1.620 -0.115 3.010 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.665 -0.115 1.500 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.680 4.570 1.375 ;
        RECT  4.205 1.145 4.490 1.375 ;
        RECT  4.135 0.975 4.205 1.375 ;
        RECT  3.835 1.145 4.135 1.375 ;
        RECT  3.765 0.905 3.835 1.375 ;
        RECT  3.465 1.145 3.765 1.375 ;
        RECT  3.395 0.990 3.465 1.375 ;
        RECT  2.750 1.145 3.395 1.375 ;
        RECT  2.630 1.030 2.750 1.375 ;
        RECT  2.030 1.145 2.630 1.375 ;
        RECT  1.910 1.005 2.030 1.375 ;
        RECT  1.670 1.145 1.910 1.375 ;
        RECT  1.550 1.000 1.670 1.375 ;
        RECT  0.690 1.145 1.550 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.030 0.355 4.095 0.485 ;
        RECT  4.025 0.735 4.095 0.905 ;
        RECT  3.960 0.185 4.030 0.485 ;
        RECT  3.955 0.735 4.025 1.065 ;
        RECT  3.865 0.545 3.920 0.615 ;
        RECT  3.795 0.215 3.865 0.805 ;
        RECT  3.370 0.215 3.795 0.285 ;
        RECT  3.645 0.735 3.795 0.805 ;
        RECT  3.575 0.735 3.645 1.035 ;
        RECT  3.285 0.850 3.575 0.920 ;
        RECT  3.385 0.520 3.455 0.780 ;
        RECT  3.135 0.710 3.385 0.780 ;
        RECT  3.215 0.850 3.285 1.045 ;
        RECT  2.880 0.975 3.215 1.045 ;
        RECT  3.065 0.710 3.135 0.905 ;
        RECT  2.365 0.835 3.065 0.905 ;
        RECT  2.505 0.695 2.930 0.765 ;
        RECT  2.505 0.375 2.705 0.455 ;
        RECT  1.790 0.200 2.510 0.270 ;
        RECT  2.435 0.375 2.505 0.765 ;
        RECT  2.270 0.375 2.435 0.455 ;
        RECT  2.295 0.570 2.365 0.905 ;
        RECT  2.185 0.570 2.295 0.640 ;
        RECT  2.005 0.710 2.210 0.780 ;
        RECT  2.140 0.860 2.210 1.075 ;
        RECT  2.115 0.350 2.185 0.640 ;
        RECT  1.360 0.860 2.140 0.930 ;
        RECT  1.935 0.350 2.005 0.780 ;
        RECT  1.600 0.710 1.935 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  0.830 0.195 1.310 0.265 ;
        RECT  0.840 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.770 0.870 0.840 1.050 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.330 0.870 0.770 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.465 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.465 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFCSNQD4BWP

MACRO DFD1BWP
    CLASS CORE ;
    FOREIGN DFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.960 0.195 3.045 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.350 2.425 0.470 ;
        RECT  2.345 0.775 2.405 0.905 ;
        RECT  2.275 0.350 2.345 0.905 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.665 -0.115 3.080 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 3.080 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.820 0.210 2.890 0.640 ;
        RECT  2.140 0.210 2.820 0.280 ;
        RECT  2.680 0.520 2.750 1.050 ;
        RECT  2.650 0.520 2.680 0.640 ;
        RECT  1.860 0.980 2.680 1.050 ;
        RECT  2.580 0.375 2.640 0.445 ;
        RECT  2.580 0.775 2.605 0.905 ;
        RECT  2.510 0.375 2.580 0.905 ;
        RECT  2.430 0.545 2.510 0.615 ;
        RECT  2.070 0.210 2.140 0.910 ;
        RECT  1.950 0.295 2.070 0.415 ;
        RECT  1.930 0.820 2.070 0.910 ;
        RECT  1.880 0.675 1.980 0.745 ;
        RECT  1.810 0.195 1.880 0.745 ;
        RECT  1.790 0.840 1.860 1.050 ;
        RECT  1.710 0.195 1.810 0.265 ;
        RECT  1.740 0.840 1.790 0.910 ;
        RECT  1.670 0.345 1.740 0.910 ;
        RECT  1.600 0.985 1.720 1.075 ;
        RECT  1.570 0.185 1.710 0.265 ;
        RECT  1.530 0.345 1.600 0.905 ;
        RECT  0.330 0.985 1.600 1.055 ;
        RECT  1.160 0.195 1.570 0.265 ;
        RECT  1.280 0.345 1.530 0.415 ;
        RECT  1.520 0.785 1.530 0.905 ;
        RECT  1.430 0.520 1.460 0.640 ;
        RECT  1.360 0.520 1.430 0.905 ;
        RECT  1.130 0.835 1.360 0.905 ;
        RECT  1.210 0.345 1.280 0.640 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.910 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFD1BWP

MACRO DFD2BWP
    CLASS CORE ;
    FOREIGN DFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 0.355 3.325 0.805 ;
        RECT  3.265 0.185 3.270 0.805 ;
        RECT  3.255 0.185 3.265 1.035 ;
        RECT  3.200 0.185 3.255 0.465 ;
        RECT  3.195 0.735 3.255 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.910 0.785 ;
        RECT  2.790 0.355 2.835 0.425 ;
        RECT  2.790 0.715 2.835 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.300 ;
        RECT  0.665 -0.115 3.370 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.895 3.450 1.375 ;
        RECT  3.100 1.145 3.370 1.375 ;
        RECT  2.980 1.020 3.100 1.375 ;
        RECT  2.720 1.145 2.980 1.375 ;
        RECT  2.600 1.010 2.720 1.375 ;
        RECT  0.000 1.145 2.600 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.110 0.545 3.180 0.615 ;
        RECT  3.040 0.215 3.110 0.940 ;
        RECT  2.090 0.215 3.040 0.285 ;
        RECT  2.520 0.870 3.040 0.940 ;
        RECT  2.700 0.520 2.765 0.640 ;
        RECT  2.630 0.375 2.700 0.800 ;
        RECT  2.230 0.375 2.630 0.445 ;
        RECT  2.440 0.680 2.630 0.800 ;
        RECT  2.450 0.870 2.520 1.050 ;
        RECT  1.990 0.980 2.450 1.050 ;
        RECT  2.370 0.540 2.420 0.610 ;
        RECT  2.300 0.540 2.370 0.910 ;
        RECT  1.810 0.840 2.300 0.910 ;
        RECT  2.160 0.375 2.230 0.615 ;
        RECT  2.090 0.545 2.160 0.615 ;
        RECT  2.020 0.215 2.090 0.355 ;
        RECT  1.950 0.510 1.995 0.770 ;
        RECT  1.925 0.195 1.950 0.770 ;
        RECT  1.880 0.195 1.925 0.580 ;
        RECT  1.760 0.195 1.880 0.265 ;
        RECT  1.740 0.345 1.810 0.910 ;
        RECT  1.650 0.985 1.770 1.075 ;
        RECT  1.610 0.185 1.760 0.265 ;
        RECT  0.330 0.985 1.650 1.055 ;
        RECT  1.570 0.345 1.640 0.905 ;
        RECT  1.160 0.195 1.610 0.265 ;
        RECT  1.295 0.345 1.570 0.415 ;
        RECT  1.560 0.785 1.570 0.905 ;
        RECT  1.470 0.520 1.500 0.640 ;
        RECT  1.400 0.520 1.470 0.905 ;
        RECT  1.130 0.835 1.400 0.905 ;
        RECT  1.225 0.345 1.295 0.640 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.910 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFD2BWP

MACRO DFD4BWP
    CLASS CORE ;
    FOREIGN DFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.765 3.965 1.065 ;
        RECT  3.815 0.355 3.895 0.465 ;
        RECT  3.815 0.765 3.895 0.905 ;
        RECT  3.605 0.355 3.815 0.905 ;
        RECT  3.585 0.355 3.605 0.465 ;
        RECT  3.515 0.765 3.605 1.065 ;
        RECT  3.515 0.185 3.585 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.710 3.250 0.800 ;
        RECT  3.115 0.355 3.230 0.445 ;
        RECT  2.905 0.355 3.115 0.800 ;
        RECT  2.730 0.355 2.905 0.445 ;
        RECT  2.770 0.710 2.905 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.465 ;
        RECT  3.775 -0.115 4.070 0.115 ;
        RECT  3.705 -0.115 3.775 0.285 ;
        RECT  0.665 -0.115 3.705 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.680 4.150 1.375 ;
        RECT  3.775 1.145 4.070 1.375 ;
        RECT  3.705 0.975 3.775 1.375 ;
        RECT  3.430 1.145 3.705 1.375 ;
        RECT  3.310 1.010 3.430 1.375 ;
        RECT  3.070 1.145 3.310 1.375 ;
        RECT  2.950 1.010 3.070 1.375 ;
        RECT  2.700 1.145 2.950 1.375 ;
        RECT  2.580 1.010 2.700 1.375 ;
        RECT  0.690 1.145 2.580 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.765 3.965 1.065 ;
        RECT  3.885 0.355 3.895 0.465 ;
        RECT  3.885 0.765 3.895 0.905 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.515 0.765 3.535 1.065 ;
        RECT  3.185 0.710 3.250 0.800 ;
        RECT  3.185 0.355 3.230 0.445 ;
        RECT  2.730 0.355 2.835 0.445 ;
        RECT  2.770 0.710 2.835 0.800 ;
        RECT  3.390 0.545 3.510 0.615 ;
        RECT  3.320 0.215 3.390 0.940 ;
        RECT  2.050 0.215 3.320 0.285 ;
        RECT  2.495 0.870 3.320 0.940 ;
        RECT  2.620 0.545 2.800 0.615 ;
        RECT  2.550 0.365 2.620 0.800 ;
        RECT  2.190 0.365 2.550 0.435 ;
        RECT  2.400 0.700 2.550 0.800 ;
        RECT  2.425 0.870 2.495 1.030 ;
        RECT  2.330 0.545 2.470 0.615 ;
        RECT  1.950 0.960 2.425 1.030 ;
        RECT  2.260 0.545 2.330 0.890 ;
        RECT  1.770 0.820 2.260 0.890 ;
        RECT  2.120 0.365 2.190 0.630 ;
        RECT  2.090 0.530 2.120 0.630 ;
        RECT  1.980 0.215 2.050 0.385 ;
        RECT  1.910 0.675 2.010 0.745 ;
        RECT  1.840 0.195 1.910 0.745 ;
        RECT  1.740 0.195 1.840 0.265 ;
        RECT  1.700 0.345 1.770 0.890 ;
        RECT  1.630 0.985 1.750 1.075 ;
        RECT  1.590 0.185 1.740 0.265 ;
        RECT  0.830 0.985 1.630 1.055 ;
        RECT  1.550 0.345 1.620 0.905 ;
        RECT  1.160 0.195 1.590 0.265 ;
        RECT  1.295 0.345 1.550 0.415 ;
        RECT  1.540 0.785 1.550 0.905 ;
        RECT  1.450 0.520 1.480 0.640 ;
        RECT  1.380 0.520 1.450 0.905 ;
        RECT  1.130 0.835 1.380 0.905 ;
        RECT  1.225 0.345 1.295 0.640 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.910 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.760 0.870 0.830 1.055 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.330 0.870 0.760 0.940 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.465 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.465 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFD4BWP

MACRO DFKCND1BWP
    CLASS CORE ;
    FOREIGN DFKCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.185 3.325 1.045 ;
        RECT  3.235 0.185 3.255 0.465 ;
        RECT  3.235 0.745 3.255 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.025 0.765 3.050 1.045 ;
        RECT  2.955 0.350 3.025 1.045 ;
        RECT  2.860 0.350 2.955 0.470 ;
        RECT  2.860 0.765 2.955 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.355 0.950 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.690 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.360 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 1.145 3.360 1.375 ;
        RECT  3.020 1.120 3.140 1.375 ;
        RECT  1.635 1.145 3.020 1.375 ;
        RECT  1.565 0.830 1.635 1.375 ;
        RECT  0.000 1.145 1.565 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.165 0.520 3.180 0.640 ;
        RECT  3.095 0.210 3.165 0.640 ;
        RECT  2.340 0.210 3.095 0.280 ;
        RECT  2.790 0.550 2.880 0.620 ;
        RECT  2.720 0.355 2.790 0.975 ;
        RECT  2.480 0.355 2.720 0.425 ;
        RECT  2.640 0.905 2.720 0.975 ;
        RECT  2.580 0.520 2.650 0.800 ;
        RECT  2.550 0.730 2.580 0.800 ;
        RECT  2.480 0.730 2.550 1.060 ;
        RECT  2.410 0.355 2.480 0.640 ;
        RECT  2.050 0.990 2.480 1.060 ;
        RECT  2.340 0.780 2.390 0.910 ;
        RECT  2.270 0.210 2.340 0.910 ;
        RECT  2.130 0.200 2.200 0.910 ;
        RECT  2.020 0.200 2.130 0.270 ;
        RECT  2.050 0.350 2.060 0.470 ;
        RECT  1.980 0.350 2.050 1.060 ;
        RECT  1.900 0.185 2.020 0.270 ;
        RECT  1.875 0.340 1.910 0.870 ;
        RECT  1.480 0.200 1.900 0.270 ;
        RECT  1.840 0.340 1.875 1.060 ;
        RECT  1.595 0.340 1.840 0.410 ;
        RECT  1.805 0.800 1.840 1.060 ;
        RECT  1.745 0.510 1.770 0.640 ;
        RECT  1.675 0.510 1.745 0.760 ;
        RECT  1.345 0.690 1.675 0.760 ;
        RECT  1.525 0.340 1.595 0.620 ;
        RECT  1.360 0.185 1.480 0.270 ;
        RECT  1.240 0.980 1.360 1.075 ;
        RECT  1.275 0.340 1.345 0.910 ;
        RECT  1.150 0.840 1.275 0.910 ;
        RECT  0.330 0.980 1.240 1.050 ;
        RECT  1.095 0.195 1.165 0.500 ;
        RECT  1.080 0.570 1.160 0.770 ;
        RECT  0.330 0.195 1.095 0.265 ;
        RECT  0.520 0.700 1.080 0.770 ;
        RECT  0.570 0.840 1.070 0.910 ;
        RECT  0.485 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.485 0.910 ;
        RECT  0.435 0.345 0.450 0.465 ;
        RECT  0.415 0.695 0.450 0.910 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.195 0.330 1.050 ;
        RECT  0.055 0.295 0.260 0.415 ;
        RECT  0.050 0.850 0.260 0.970 ;
    END
END DFKCND1BWP

MACRO DFKCND2BWP
    CLASS CORE ;
    FOREIGN DFKCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.545 0.355 3.605 0.805 ;
        RECT  3.535 0.185 3.545 1.035 ;
        RECT  3.475 0.185 3.535 0.465 ;
        RECT  3.475 0.735 3.535 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.355 3.185 1.045 ;
        RECT  3.095 0.355 3.115 0.475 ;
        RECT  3.095 0.745 3.115 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.355 0.950 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.690 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.300 ;
        RECT  0.000 -0.115 3.650 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.895 3.730 1.375 ;
        RECT  3.355 1.145 3.650 1.375 ;
        RECT  3.285 0.745 3.355 1.375 ;
        RECT  3.000 1.145 3.285 1.375 ;
        RECT  2.880 1.010 3.000 1.375 ;
        RECT  2.620 1.145 2.880 1.375 ;
        RECT  2.500 1.010 2.620 1.375 ;
        RECT  1.655 1.145 2.500 1.375 ;
        RECT  1.585 0.850 1.655 1.375 ;
        RECT  0.000 1.145 1.585 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.370 0.545 3.460 0.615 ;
        RECT  3.300 0.215 3.370 0.615 ;
        RECT  2.400 0.215 3.300 0.285 ;
        RECT  2.980 0.520 3.040 0.640 ;
        RECT  2.910 0.365 2.980 0.940 ;
        RECT  2.540 0.365 2.910 0.435 ;
        RECT  2.680 0.870 2.910 0.940 ;
        RECT  2.645 0.520 2.715 0.800 ;
        RECT  2.590 0.730 2.645 0.800 ;
        RECT  2.520 0.730 2.590 0.940 ;
        RECT  2.470 0.365 2.540 0.640 ;
        RECT  2.430 0.870 2.520 0.940 ;
        RECT  2.360 0.870 2.430 1.060 ;
        RECT  2.330 0.195 2.400 0.790 ;
        RECT  2.080 0.990 2.360 1.060 ;
        RECT  2.170 0.200 2.240 0.910 ;
        RECT  2.060 0.200 2.170 0.270 ;
        RECT  2.150 0.790 2.170 0.910 ;
        RECT  2.080 0.350 2.100 0.470 ;
        RECT  2.010 0.350 2.080 1.060 ;
        RECT  1.940 0.185 2.060 0.270 ;
        RECT  1.480 0.200 1.940 0.270 ;
        RECT  1.905 0.340 1.930 0.890 ;
        RECT  1.860 0.340 1.905 1.060 ;
        RECT  1.610 0.340 1.860 0.410 ;
        RECT  1.835 0.800 1.860 1.060 ;
        RECT  1.760 0.510 1.790 0.640 ;
        RECT  1.690 0.510 1.760 0.780 ;
        RECT  1.345 0.710 1.690 0.780 ;
        RECT  1.540 0.340 1.610 0.640 ;
        RECT  1.360 0.185 1.480 0.270 ;
        RECT  1.240 0.980 1.360 1.075 ;
        RECT  1.275 0.340 1.345 0.910 ;
        RECT  1.150 0.840 1.275 0.910 ;
        RECT  0.330 0.980 1.240 1.050 ;
        RECT  1.095 0.195 1.165 0.500 ;
        RECT  1.080 0.570 1.160 0.770 ;
        RECT  0.330 0.195 1.095 0.265 ;
        RECT  0.520 0.700 1.080 0.770 ;
        RECT  0.570 0.840 1.070 0.910 ;
        RECT  0.485 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.485 0.910 ;
        RECT  0.435 0.345 0.450 0.465 ;
        RECT  0.415 0.695 0.450 0.910 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.195 0.330 1.050 ;
        RECT  0.055 0.295 0.260 0.415 ;
        RECT  0.050 0.850 0.260 0.970 ;
    END
END DFKCND2BWP

MACRO DFKCND4BWP
    CLASS CORE ;
    FOREIGN DFKCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.185 4.245 0.465 ;
        RECT  4.235 0.765 4.245 1.065 ;
        RECT  4.175 0.185 4.235 1.065 ;
        RECT  4.025 0.355 4.175 0.905 ;
        RECT  3.885 0.355 4.025 0.465 ;
        RECT  3.885 0.765 4.025 0.905 ;
        RECT  3.815 0.185 3.885 0.465 ;
        RECT  3.815 0.765 3.885 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.355 3.530 0.450 ;
        RECT  3.435 0.765 3.505 1.065 ;
        RECT  3.395 0.765 3.435 0.905 ;
        RECT  3.185 0.355 3.395 0.905 ;
        RECT  3.030 0.355 3.185 0.450 ;
        RECT  3.125 0.765 3.185 0.905 ;
        RECT  3.055 0.765 3.125 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.975 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.695 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.465 ;
        RECT  4.090 -0.115 4.350 0.115 ;
        RECT  3.970 -0.115 4.090 0.275 ;
        RECT  0.000 -0.115 3.970 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.680 4.430 1.375 ;
        RECT  4.065 1.145 4.350 1.375 ;
        RECT  3.995 0.975 4.065 1.375 ;
        RECT  3.695 1.145 3.995 1.375 ;
        RECT  3.625 0.745 3.695 1.375 ;
        RECT  3.325 1.145 3.625 1.375 ;
        RECT  3.235 0.975 3.325 1.375 ;
        RECT  1.655 1.145 3.235 1.375 ;
        RECT  1.585 0.850 1.655 1.375 ;
        RECT  0.000 1.145 1.585 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.355 3.955 0.465 ;
        RECT  3.885 0.765 3.955 0.905 ;
        RECT  3.815 0.185 3.885 0.465 ;
        RECT  3.815 0.765 3.885 1.065 ;
        RECT  3.465 0.355 3.530 0.450 ;
        RECT  3.465 0.765 3.505 1.065 ;
        RECT  3.030 0.355 3.115 0.450 ;
        RECT  3.055 0.765 3.115 1.065 ;
        RECT  3.700 0.545 3.850 0.615 ;
        RECT  3.630 0.215 3.700 0.615 ;
        RECT  2.360 0.215 3.630 0.285 ;
        RECT  2.910 0.545 3.060 0.615 ;
        RECT  2.840 0.355 2.910 1.000 ;
        RECT  2.500 0.355 2.840 0.425 ;
        RECT  2.650 0.930 2.840 1.000 ;
        RECT  2.675 0.510 2.745 0.850 ;
        RECT  2.540 0.780 2.675 0.850 ;
        RECT  2.470 0.780 2.540 1.060 ;
        RECT  2.430 0.355 2.500 0.640 ;
        RECT  2.070 0.990 2.470 1.060 ;
        RECT  2.290 0.195 2.360 0.800 ;
        RECT  2.150 0.200 2.220 0.920 ;
        RECT  2.020 0.200 2.150 0.270 ;
        RECT  2.070 0.350 2.080 0.470 ;
        RECT  2.000 0.350 2.070 1.060 ;
        RECT  1.900 0.185 2.020 0.270 ;
        RECT  1.895 0.350 1.930 0.840 ;
        RECT  1.480 0.200 1.900 0.270 ;
        RECT  1.860 0.350 1.895 1.060 ;
        RECT  1.595 0.350 1.860 0.420 ;
        RECT  1.825 0.770 1.860 1.060 ;
        RECT  1.755 0.510 1.790 0.640 ;
        RECT  1.685 0.510 1.755 0.780 ;
        RECT  1.345 0.710 1.685 0.780 ;
        RECT  1.525 0.350 1.595 0.640 ;
        RECT  1.360 0.185 1.480 0.270 ;
        RECT  1.260 0.980 1.380 1.075 ;
        RECT  1.275 0.340 1.345 0.910 ;
        RECT  1.170 0.840 1.275 0.910 ;
        RECT  0.350 0.980 1.260 1.050 ;
        RECT  1.105 0.570 1.175 0.770 ;
        RECT  1.095 0.215 1.165 0.500 ;
        RECT  0.515 0.700 1.105 0.770 ;
        RECT  0.350 0.215 1.095 0.285 ;
        RECT  0.590 0.840 1.090 0.910 ;
        RECT  0.505 0.355 0.515 0.770 ;
        RECT  0.445 0.355 0.505 0.910 ;
        RECT  0.435 0.355 0.445 0.475 ;
        RECT  0.435 0.695 0.445 0.910 ;
        RECT  0.350 0.520 0.375 0.640 ;
        RECT  0.280 0.215 0.350 1.050 ;
        RECT  0.055 0.215 0.280 0.335 ;
        RECT  0.050 0.930 0.280 1.050 ;
    END
END DFKCND4BWP

MACRO DFKCNQD1BWP
    CLASS CORE ;
    FOREIGN DFKCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.185 3.045 1.045 ;
        RECT  2.955 0.185 2.975 0.465 ;
        RECT  2.955 0.735 2.975 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.355 0.950 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.690 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 -0.115 3.080 0.115 ;
        RECT  2.740 -0.115 2.860 0.280 ;
        RECT  2.465 -0.115 2.740 0.115 ;
        RECT  2.395 -0.115 2.465 0.305 ;
        RECT  0.000 -0.115 2.395 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.835 1.145 3.080 1.375 ;
        RECT  2.765 0.905 2.835 1.375 ;
        RECT  1.635 1.145 2.765 1.375 ;
        RECT  1.565 0.850 1.635 1.375 ;
        RECT  0.000 1.145 1.565 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.885 0.520 2.905 0.640 ;
        RECT  2.815 0.375 2.885 0.805 ;
        RECT  2.645 0.375 2.815 0.445 ;
        RECT  2.650 0.735 2.815 0.805 ;
        RECT  2.510 0.545 2.740 0.615 ;
        RECT  2.580 0.735 2.650 1.035 ;
        RECT  2.575 0.185 2.645 0.445 ;
        RECT  2.370 0.375 2.575 0.445 ;
        RECT  2.440 0.545 2.510 1.060 ;
        RECT  2.050 0.990 2.440 1.060 ;
        RECT  2.300 0.375 2.370 0.640 ;
        RECT  2.140 0.200 2.210 0.910 ;
        RECT  2.020 0.200 2.140 0.270 ;
        RECT  2.050 0.350 2.065 0.470 ;
        RECT  1.980 0.350 2.050 1.060 ;
        RECT  1.900 0.185 2.020 0.270 ;
        RECT  1.885 0.360 1.910 0.840 ;
        RECT  1.480 0.200 1.900 0.270 ;
        RECT  1.840 0.360 1.885 1.060 ;
        RECT  1.595 0.360 1.840 0.430 ;
        RECT  1.815 0.770 1.840 1.060 ;
        RECT  1.745 0.510 1.770 0.640 ;
        RECT  1.675 0.510 1.745 0.780 ;
        RECT  1.345 0.710 1.675 0.780 ;
        RECT  1.525 0.360 1.595 0.640 ;
        RECT  1.360 0.185 1.480 0.270 ;
        RECT  1.240 0.980 1.360 1.075 ;
        RECT  1.275 0.340 1.345 0.910 ;
        RECT  1.150 0.840 1.275 0.910 ;
        RECT  0.330 0.980 1.240 1.050 ;
        RECT  1.095 0.195 1.165 0.500 ;
        RECT  1.080 0.570 1.160 0.770 ;
        RECT  0.330 0.195 1.095 0.265 ;
        RECT  0.520 0.700 1.080 0.770 ;
        RECT  0.570 0.840 1.070 0.910 ;
        RECT  0.485 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.485 0.910 ;
        RECT  0.435 0.345 0.450 0.465 ;
        RECT  0.415 0.695 0.450 0.910 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.195 0.330 1.050 ;
        RECT  0.055 0.295 0.260 0.415 ;
        RECT  0.050 0.850 0.260 0.970 ;
    END
END DFKCNQD1BWP

MACRO DFKCNQD2BWP
    CLASS CORE ;
    FOREIGN DFKCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.355 3.045 0.835 ;
        RECT  2.975 0.185 2.985 1.035 ;
        RECT  2.915 0.185 2.975 0.465 ;
        RECT  2.915 0.735 2.975 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.355 0.950 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.690 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.300 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.275 ;
        RECT  2.470 -0.115 2.710 0.115 ;
        RECT  2.350 -0.115 2.470 0.275 ;
        RECT  0.000 -0.115 2.350 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.905 3.170 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.010 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.380 0.950 2.450 1.375 ;
        RECT  1.645 1.145 2.380 1.375 ;
        RECT  1.575 0.835 1.645 1.375 ;
        RECT  0.000 1.145 1.575 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.545 2.900 0.615 ;
        RECT  2.680 0.370 2.750 0.940 ;
        RECT  2.625 0.370 2.680 0.440 ;
        RECT  2.530 0.870 2.680 0.940 ;
        RECT  2.555 0.185 2.625 0.440 ;
        RECT  2.355 0.370 2.555 0.440 ;
        RECT  2.485 0.510 2.555 0.790 ;
        RECT  2.310 0.720 2.485 0.790 ;
        RECT  2.285 0.370 2.355 0.640 ;
        RECT  2.240 0.720 2.310 1.060 ;
        RECT  2.030 0.990 2.240 1.060 ;
        RECT  2.170 0.200 2.185 0.620 ;
        RECT  2.115 0.200 2.170 0.910 ;
        RECT  2.000 0.200 2.115 0.270 ;
        RECT  2.100 0.550 2.115 0.910 ;
        RECT  2.030 0.350 2.045 0.470 ;
        RECT  1.960 0.350 2.030 1.060 ;
        RECT  1.870 0.185 2.000 0.270 ;
        RECT  1.820 0.345 1.890 0.930 ;
        RECT  1.430 0.200 1.870 0.270 ;
        RECT  1.575 0.345 1.820 0.415 ;
        RECT  1.730 0.860 1.820 0.930 ;
        RECT  1.680 0.500 1.750 0.765 ;
        RECT  1.290 0.695 1.680 0.765 ;
        RECT  1.505 0.345 1.575 0.625 ;
        RECT  1.360 0.200 1.430 0.320 ;
        RECT  1.240 0.980 1.360 1.075 ;
        RECT  1.220 0.185 1.290 0.910 ;
        RECT  0.330 0.980 1.240 1.050 ;
        RECT  1.180 0.185 1.220 0.305 ;
        RECT  1.150 0.840 1.220 0.910 ;
        RECT  1.090 0.370 1.150 0.500 ;
        RECT  1.070 0.570 1.140 0.770 ;
        RECT  1.020 0.195 1.090 0.500 ;
        RECT  0.520 0.700 1.070 0.770 ;
        RECT  0.570 0.840 1.070 0.910 ;
        RECT  0.330 0.195 1.020 0.265 ;
        RECT  0.485 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.485 0.910 ;
        RECT  0.435 0.345 0.450 0.465 ;
        RECT  0.415 0.695 0.450 0.910 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.195 0.330 1.050 ;
        RECT  0.055 0.295 0.260 0.415 ;
        RECT  0.050 0.850 0.260 0.970 ;
    END
END DFKCNQD2BWP

MACRO DFKCNQD4BWP
    CLASS CORE ;
    FOREIGN DFKCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.185 3.405 0.465 ;
        RECT  3.395 0.765 3.405 1.065 ;
        RECT  3.335 0.185 3.395 1.065 ;
        RECT  3.185 0.355 3.335 0.905 ;
        RECT  3.045 0.355 3.185 0.465 ;
        RECT  3.045 0.765 3.185 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.765 3.045 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.355 0.970 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.695 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.640 0.115 ;
        RECT  3.510 -0.115 3.590 0.465 ;
        RECT  3.250 -0.115 3.510 0.115 ;
        RECT  3.130 -0.115 3.250 0.275 ;
        RECT  2.890 -0.115 3.130 0.115 ;
        RECT  2.770 -0.115 2.890 0.275 ;
        RECT  2.530 -0.115 2.770 0.115 ;
        RECT  2.410 -0.115 2.530 0.275 ;
        RECT  0.000 -0.115 2.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.680 3.590 1.375 ;
        RECT  3.230 1.145 3.510 1.375 ;
        RECT  3.150 0.975 3.230 1.375 ;
        RECT  2.890 1.145 3.150 1.375 ;
        RECT  2.770 1.010 2.890 1.375 ;
        RECT  1.670 1.145 2.770 1.375 ;
        RECT  1.570 0.860 1.670 1.375 ;
        RECT  0.000 1.145 1.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.355 3.115 0.465 ;
        RECT  3.045 0.765 3.115 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.765 3.045 1.065 ;
        RECT  2.870 0.545 3.010 0.615 ;
        RECT  2.800 0.370 2.870 0.940 ;
        RECT  2.685 0.370 2.800 0.440 ;
        RECT  2.590 0.870 2.800 0.940 ;
        RECT  2.615 0.185 2.685 0.440 ;
        RECT  2.555 0.510 2.625 0.790 ;
        RECT  2.415 0.370 2.615 0.440 ;
        RECT  2.415 0.720 2.555 0.790 ;
        RECT  2.345 0.370 2.415 0.640 ;
        RECT  2.345 0.720 2.415 1.050 ;
        RECT  2.080 0.980 2.345 1.050 ;
        RECT  2.170 0.200 2.240 0.910 ;
        RECT  2.060 0.200 2.170 0.270 ;
        RECT  2.150 0.790 2.170 0.910 ;
        RECT  2.080 0.350 2.100 0.470 ;
        RECT  2.010 0.350 2.080 1.050 ;
        RECT  1.930 0.185 2.060 0.270 ;
        RECT  1.500 0.200 1.930 0.270 ;
        RECT  1.895 0.350 1.930 0.840 ;
        RECT  1.860 0.350 1.895 1.060 ;
        RECT  1.615 0.350 1.860 0.420 ;
        RECT  1.825 0.770 1.860 1.060 ;
        RECT  1.755 0.510 1.790 0.640 ;
        RECT  1.685 0.510 1.755 0.790 ;
        RECT  1.365 0.720 1.685 0.790 ;
        RECT  1.545 0.350 1.615 0.640 ;
        RECT  1.380 0.185 1.500 0.270 ;
        RECT  1.260 0.980 1.380 1.075 ;
        RECT  1.295 0.340 1.365 0.910 ;
        RECT  1.170 0.840 1.295 0.910 ;
        RECT  0.350 0.980 1.260 1.050 ;
        RECT  1.115 0.215 1.185 0.500 ;
        RECT  1.105 0.570 1.175 0.770 ;
        RECT  0.350 0.215 1.115 0.285 ;
        RECT  0.515 0.700 1.105 0.770 ;
        RECT  0.590 0.840 1.090 0.910 ;
        RECT  0.505 0.355 0.515 0.770 ;
        RECT  0.445 0.355 0.505 0.910 ;
        RECT  0.435 0.355 0.445 0.475 ;
        RECT  0.435 0.695 0.445 0.910 ;
        RECT  0.350 0.520 0.375 0.640 ;
        RECT  0.280 0.215 0.350 1.050 ;
        RECT  0.055 0.215 0.280 0.335 ;
        RECT  0.050 0.930 0.280 1.050 ;
    END
END DFKCNQD4BWP

MACRO DFKCSND1BWP
    CLASS CORE ;
    FOREIGN DFKCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.770 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.185 3.745 1.045 ;
        RECT  3.655 0.185 3.675 0.465 ;
        RECT  3.655 0.745 3.675 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.445 0.765 3.470 1.045 ;
        RECT  3.375 0.350 3.445 1.045 ;
        RECT  3.280 0.350 3.375 0.470 ;
        RECT  3.280 0.765 3.375 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.680 0.555 0.800 ;
        RECT  0.455 0.680 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.100 0.770 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.770 ;
        RECT  0.830 0.700 0.875 0.770 ;
        RECT  0.735 0.700 0.830 0.925 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.780 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.145 3.780 1.375 ;
        RECT  2.040 0.860 2.160 1.375 ;
        RECT  0.330 1.145 2.040 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.585 0.520 3.600 0.640 ;
        RECT  3.515 0.210 3.585 0.640 ;
        RECT  2.780 0.210 3.515 0.280 ;
        RECT  3.210 0.550 3.300 0.620 ;
        RECT  3.140 0.355 3.210 0.860 ;
        RECT  3.070 0.990 3.190 1.075 ;
        RECT  2.920 0.355 3.140 0.425 ;
        RECT  3.060 0.790 3.140 0.860 ;
        RECT  2.490 0.990 3.070 1.060 ;
        RECT  2.850 0.355 2.920 0.640 ;
        RECT  2.780 0.780 2.810 0.910 ;
        RECT  2.710 0.210 2.780 0.910 ;
        RECT  2.570 0.195 2.640 0.910 ;
        RECT  2.470 0.195 2.570 0.265 ;
        RECT  2.560 0.790 2.570 0.910 ;
        RECT  2.490 0.350 2.500 0.470 ;
        RECT  2.420 0.350 2.490 1.060 ;
        RECT  2.350 0.185 2.470 0.265 ;
        RECT  1.800 0.195 2.350 0.265 ;
        RECT  2.280 0.360 2.350 0.960 ;
        RECT  2.035 0.360 2.280 0.430 ;
        RECT  2.260 0.840 2.280 0.960 ;
        RECT  2.140 0.510 2.210 0.780 ;
        RECT  1.785 0.710 2.140 0.780 ;
        RECT  1.965 0.360 2.035 0.640 ;
        RECT  1.765 0.350 1.785 0.780 ;
        RECT  1.715 0.350 1.765 0.960 ;
        RECT  1.695 0.690 1.715 0.960 ;
        RECT  0.700 0.195 1.610 0.265 ;
        RECT  1.380 0.865 1.610 0.935 ;
        RECT  1.505 0.345 1.575 0.785 ;
        RECT  1.310 0.345 1.505 0.415 ;
        RECT  1.310 0.715 1.505 0.785 ;
        RECT  1.310 0.865 1.380 1.065 ;
        RECT  1.240 0.545 1.340 0.615 ;
        RECT  0.665 0.995 1.310 1.065 ;
        RECT  1.170 0.345 1.240 0.925 ;
        RECT  0.950 0.345 1.170 0.415 ;
        RECT  0.930 0.855 1.170 0.925 ;
        RECT  0.780 0.360 0.880 0.460 ;
        RECT  0.500 0.390 0.780 0.460 ;
        RECT  0.375 0.540 0.780 0.610 ;
        RECT  0.580 0.195 0.700 0.310 ;
        RECT  0.595 0.925 0.665 1.065 ;
        RECT  0.400 0.360 0.500 0.460 ;
        RECT  0.330 0.540 0.375 0.940 ;
        RECT  0.305 0.310 0.330 0.940 ;
        RECT  0.260 0.310 0.305 0.610 ;
        RECT  0.125 0.870 0.305 0.940 ;
        RECT  0.125 0.310 0.260 0.380 ;
        RECT  0.055 0.230 0.125 0.380 ;
        RECT  0.055 0.870 0.125 1.030 ;
    END
END DFKCSND1BWP

MACRO DFKCSND2BWP
    CLASS CORE ;
    FOREIGN DFKCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.770 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.355 4.025 0.805 ;
        RECT  3.955 0.185 3.965 1.035 ;
        RECT  3.895 0.185 3.955 0.465 ;
        RECT  3.895 0.735 3.955 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.350 3.605 1.045 ;
        RECT  3.515 0.350 3.535 0.470 ;
        RECT  3.515 0.735 3.535 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.680 0.555 0.800 ;
        RECT  0.455 0.680 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.100 0.770 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0156 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.770 ;
        RECT  0.830 0.700 0.875 0.770 ;
        RECT  0.735 0.700 0.830 0.925 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.300 ;
        RECT  0.000 -0.115 4.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.895 4.150 1.375 ;
        RECT  3.775 1.145 4.070 1.375 ;
        RECT  3.705 0.735 3.775 1.375 ;
        RECT  2.180 1.145 3.705 1.375 ;
        RECT  2.060 0.860 2.180 1.375 ;
        RECT  0.330 1.145 2.060 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.800 0.545 3.880 0.615 ;
        RECT  3.730 0.210 3.800 0.615 ;
        RECT  2.800 0.210 3.730 0.280 ;
        RECT  3.380 0.520 3.465 0.640 ;
        RECT  3.310 0.365 3.380 1.000 ;
        RECT  2.940 0.365 3.310 0.435 ;
        RECT  3.110 0.930 3.310 1.000 ;
        RECT  3.065 0.520 3.135 0.860 ;
        RECT  3.020 0.790 3.065 0.860 ;
        RECT  2.950 0.790 3.020 1.010 ;
        RECT  2.810 0.940 2.950 1.010 ;
        RECT  2.870 0.365 2.940 0.640 ;
        RECT  2.800 0.730 2.830 0.860 ;
        RECT  2.740 0.940 2.810 1.060 ;
        RECT  2.730 0.210 2.800 0.860 ;
        RECT  2.510 0.990 2.740 1.060 ;
        RECT  2.590 0.195 2.660 0.910 ;
        RECT  2.490 0.195 2.590 0.265 ;
        RECT  2.580 0.790 2.590 0.910 ;
        RECT  2.510 0.350 2.520 0.470 ;
        RECT  2.440 0.350 2.510 1.060 ;
        RECT  2.360 0.185 2.490 0.265 ;
        RECT  2.300 0.360 2.370 0.960 ;
        RECT  1.800 0.195 2.360 0.265 ;
        RECT  2.055 0.360 2.300 0.430 ;
        RECT  2.280 0.840 2.300 0.960 ;
        RECT  2.160 0.510 2.230 0.780 ;
        RECT  1.785 0.710 2.160 0.780 ;
        RECT  1.985 0.360 2.055 0.640 ;
        RECT  1.765 0.350 1.785 0.780 ;
        RECT  1.715 0.350 1.765 0.960 ;
        RECT  1.695 0.690 1.715 0.960 ;
        RECT  0.700 0.195 1.610 0.265 ;
        RECT  1.380 0.865 1.610 0.935 ;
        RECT  1.505 0.345 1.575 0.785 ;
        RECT  1.310 0.345 1.505 0.415 ;
        RECT  1.310 0.715 1.505 0.785 ;
        RECT  1.310 0.865 1.380 1.065 ;
        RECT  1.240 0.545 1.340 0.615 ;
        RECT  0.665 0.995 1.310 1.065 ;
        RECT  1.170 0.345 1.240 0.925 ;
        RECT  0.950 0.345 1.170 0.415 ;
        RECT  0.930 0.855 1.170 0.925 ;
        RECT  0.780 0.360 0.880 0.460 ;
        RECT  0.500 0.390 0.780 0.460 ;
        RECT  0.375 0.540 0.780 0.610 ;
        RECT  0.580 0.195 0.700 0.310 ;
        RECT  0.595 0.925 0.665 1.065 ;
        RECT  0.400 0.360 0.500 0.460 ;
        RECT  0.330 0.540 0.375 0.940 ;
        RECT  0.305 0.310 0.330 0.940 ;
        RECT  0.260 0.310 0.305 0.610 ;
        RECT  0.125 0.870 0.305 0.940 ;
        RECT  0.125 0.310 0.260 0.380 ;
        RECT  0.055 0.230 0.125 0.380 ;
        RECT  0.055 0.870 0.125 1.030 ;
    END
END DFKCSND2BWP

MACRO DFKCSND4BWP
    CLASS CORE ;
    FOREIGN DFKCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.770 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.805 0.465 ;
        RECT  4.795 0.765 4.805 1.065 ;
        RECT  4.735 0.185 4.795 1.065 ;
        RECT  4.585 0.355 4.735 0.905 ;
        RECT  4.445 0.355 4.585 0.465 ;
        RECT  4.445 0.765 4.585 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.765 4.445 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.355 4.050 0.455 ;
        RECT  3.955 0.765 4.025 1.065 ;
        RECT  3.745 0.355 3.955 0.905 ;
        RECT  3.550 0.355 3.745 0.455 ;
        RECT  3.645 0.765 3.745 0.905 ;
        RECT  3.575 0.765 3.645 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.680 0.555 0.800 ;
        RECT  0.455 0.680 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.110 0.770 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0156 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.770 ;
        RECT  0.830 0.700 0.875 0.770 ;
        RECT  0.735 0.700 0.830 0.920 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.465 ;
        RECT  4.650 -0.115 4.910 0.115 ;
        RECT  4.530 -0.115 4.650 0.275 ;
        RECT  0.000 -0.115 4.530 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.675 4.990 1.375 ;
        RECT  4.625 1.145 4.910 1.375 ;
        RECT  4.555 0.975 4.625 1.375 ;
        RECT  4.240 1.145 4.555 1.375 ;
        RECT  4.160 0.735 4.240 1.375 ;
        RECT  3.835 1.145 4.160 1.375 ;
        RECT  3.765 0.975 3.835 1.375 ;
        RECT  3.480 1.145 3.765 1.375 ;
        RECT  3.360 1.010 3.480 1.375 ;
        RECT  3.080 1.145 3.360 1.375 ;
        RECT  2.960 1.010 3.080 1.375 ;
        RECT  2.200 1.145 2.960 1.375 ;
        RECT  2.080 0.860 2.200 1.375 ;
        RECT  0.330 1.145 2.080 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.355 4.515 0.465 ;
        RECT  4.445 0.765 4.515 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.765 4.445 1.065 ;
        RECT  4.025 0.355 4.050 0.455 ;
        RECT  3.550 0.355 3.675 0.455 ;
        RECT  3.645 0.765 3.675 0.905 ;
        RECT  3.575 0.765 3.645 1.065 ;
        RECT  4.250 0.545 4.410 0.615 ;
        RECT  4.180 0.215 4.250 0.615 ;
        RECT  2.845 0.215 4.180 0.285 ;
        RECT  3.430 0.545 3.580 0.615 ;
        RECT  3.360 0.365 3.430 0.940 ;
        RECT  2.985 0.365 3.360 0.435 ;
        RECT  3.160 0.870 3.360 0.940 ;
        RECT  3.195 0.520 3.265 0.790 ;
        RECT  3.090 0.720 3.195 0.790 ;
        RECT  3.020 0.720 3.090 0.940 ;
        RECT  2.820 0.870 3.020 0.940 ;
        RECT  2.915 0.365 2.985 0.640 ;
        RECT  2.775 0.185 2.845 0.800 ;
        RECT  2.750 0.870 2.820 1.060 ;
        RECT  2.530 0.990 2.750 1.060 ;
        RECT  2.610 0.195 2.680 0.910 ;
        RECT  2.510 0.195 2.610 0.265 ;
        RECT  2.600 0.790 2.610 0.910 ;
        RECT  2.530 0.350 2.540 0.470 ;
        RECT  2.460 0.350 2.530 1.060 ;
        RECT  2.380 0.185 2.510 0.265 ;
        RECT  2.320 0.360 2.390 0.950 ;
        RECT  1.820 0.195 2.380 0.265 ;
        RECT  2.075 0.360 2.320 0.430 ;
        RECT  2.300 0.830 2.320 0.950 ;
        RECT  2.180 0.510 2.250 0.780 ;
        RECT  1.805 0.710 2.180 0.780 ;
        RECT  2.005 0.360 2.075 0.640 ;
        RECT  1.785 0.350 1.805 0.780 ;
        RECT  1.735 0.350 1.785 0.960 ;
        RECT  1.715 0.690 1.735 0.960 ;
        RECT  0.580 0.200 1.640 0.270 ;
        RECT  1.400 0.865 1.630 0.935 ;
        RECT  1.525 0.350 1.595 0.785 ;
        RECT  1.330 0.350 1.525 0.420 ;
        RECT  1.330 0.715 1.525 0.785 ;
        RECT  1.330 0.865 1.400 1.060 ;
        RECT  1.260 0.545 1.340 0.615 ;
        RECT  0.665 0.990 1.330 1.060 ;
        RECT  1.190 0.350 1.260 0.920 ;
        RECT  0.950 0.350 1.190 0.420 ;
        RECT  0.950 0.850 1.190 0.920 ;
        RECT  0.795 0.350 0.865 0.470 ;
        RECT  0.485 0.350 0.795 0.420 ;
        RECT  0.375 0.540 0.780 0.610 ;
        RECT  0.595 0.920 0.665 1.060 ;
        RECT  0.415 0.350 0.485 0.470 ;
        RECT  0.330 0.540 0.375 0.940 ;
        RECT  0.305 0.310 0.330 0.940 ;
        RECT  0.260 0.310 0.305 0.610 ;
        RECT  0.125 0.870 0.305 0.940 ;
        RECT  0.125 0.310 0.260 0.380 ;
        RECT  0.055 0.230 0.125 0.380 ;
        RECT  0.055 0.870 0.125 1.030 ;
    END
END DFKCSND4BWP

MACRO DFKSND1BWP
    CLASS CORE ;
    FOREIGN DFKSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.720 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.045 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.515 0.745 3.535 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.305 0.765 3.330 1.045 ;
        RECT  3.235 0.350 3.305 1.045 ;
        RECT  3.140 0.350 3.235 0.470 ;
        RECT  3.140 0.765 3.235 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.640 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.145 3.640 1.375 ;
        RECT  3.300 1.120 3.420 1.375 ;
        RECT  2.050 1.145 3.300 1.375 ;
        RECT  1.930 0.845 2.050 1.375 ;
        RECT  0.000 1.145 1.930 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.445 0.520 3.460 0.640 ;
        RECT  3.375 0.210 3.445 0.640 ;
        RECT  2.640 0.210 3.375 0.280 ;
        RECT  3.070 0.550 3.160 0.620 ;
        RECT  3.000 0.355 3.070 0.860 ;
        RECT  2.930 0.990 3.050 1.075 ;
        RECT  2.780 0.355 3.000 0.425 ;
        RECT  2.920 0.790 3.000 0.860 ;
        RECT  2.350 0.990 2.930 1.060 ;
        RECT  2.710 0.355 2.780 0.620 ;
        RECT  2.570 0.210 2.640 0.780 ;
        RECT  2.430 0.195 2.500 0.920 ;
        RECT  2.320 0.195 2.430 0.265 ;
        RECT  2.350 0.350 2.360 0.470 ;
        RECT  2.280 0.350 2.350 1.060 ;
        RECT  2.200 0.185 2.320 0.265 ;
        RECT  2.140 0.360 2.210 1.020 ;
        RECT  1.700 0.195 2.200 0.265 ;
        RECT  1.855 0.360 2.140 0.430 ;
        RECT  2.000 0.510 2.070 0.770 ;
        RECT  1.635 0.700 2.000 0.770 ;
        RECT  1.785 0.360 1.855 0.600 ;
        RECT  1.340 0.995 1.760 1.065 ;
        RECT  1.580 0.185 1.700 0.265 ;
        RECT  1.565 0.700 1.635 0.920 ;
        RECT  0.485 0.195 1.580 0.265 ;
        RECT  1.495 0.335 1.565 0.770 ;
        RECT  1.410 0.850 1.450 0.920 ;
        RECT  1.340 0.345 1.410 0.920 ;
        RECT  0.930 0.345 1.340 0.415 ;
        RECT  1.110 0.850 1.340 0.920 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  0.330 0.995 1.220 1.065 ;
        RECT  0.860 0.520 0.915 0.640 ;
        RECT  0.790 0.345 0.860 0.915 ;
        RECT  0.570 0.345 0.790 0.415 ;
        RECT  0.570 0.845 0.790 0.915 ;
        RECT  0.415 0.195 0.485 0.910 ;
        RECT  0.260 0.340 0.330 1.065 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.995 0.260 1.065 ;
        RECT  0.055 0.280 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.065 ;
    END
END DFKSND1BWP

MACRO DFKSND2BWP
    CLASS CORE ;
    FOREIGN DFKSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.720 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 0.355 3.885 0.805 ;
        RECT  3.825 0.185 3.830 0.805 ;
        RECT  3.815 0.185 3.825 1.035 ;
        RECT  3.760 0.185 3.815 0.465 ;
        RECT  3.755 0.735 3.815 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 0.375 3.540 0.805 ;
        RECT  3.350 0.375 3.470 0.445 ;
        RECT  3.465 0.735 3.470 0.805 ;
        RECT  3.395 0.735 3.465 1.050 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.010 0.300 ;
        RECT  0.000 -0.115 3.935 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.895 4.010 1.375 ;
        RECT  3.645 1.145 3.930 1.375 ;
        RECT  3.575 0.895 3.645 1.375 ;
        RECT  3.285 1.145 3.575 1.375 ;
        RECT  3.215 0.895 3.285 1.375 ;
        RECT  2.050 1.145 3.215 1.375 ;
        RECT  1.930 0.845 2.050 1.375 ;
        RECT  0.000 1.145 1.930 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.680 0.545 3.740 0.615 ;
        RECT  3.610 0.210 3.680 0.615 ;
        RECT  2.670 0.210 3.610 0.280 ;
        RECT  3.280 0.545 3.400 0.615 ;
        RECT  3.210 0.365 3.280 0.805 ;
        RECT  2.810 0.365 3.210 0.435 ;
        RECT  3.105 0.735 3.210 0.805 ;
        RECT  3.035 0.735 3.105 1.035 ;
        RECT  2.950 0.545 3.030 0.615 ;
        RECT  2.880 0.545 2.950 1.060 ;
        RECT  2.350 0.990 2.880 1.060 ;
        RECT  2.740 0.365 2.810 0.640 ;
        RECT  2.670 0.780 2.690 0.910 ;
        RECT  2.600 0.185 2.670 0.910 ;
        RECT  2.450 0.195 2.520 0.920 ;
        RECT  2.350 0.195 2.450 0.265 ;
        RECT  2.425 0.800 2.450 0.920 ;
        RECT  2.350 0.350 2.380 0.470 ;
        RECT  2.220 0.185 2.350 0.265 ;
        RECT  2.280 0.350 2.350 1.060 ;
        RECT  1.700 0.195 2.220 0.265 ;
        RECT  2.140 0.360 2.210 1.020 ;
        RECT  1.855 0.360 2.140 0.430 ;
        RECT  2.000 0.510 2.070 0.770 ;
        RECT  1.635 0.700 2.000 0.770 ;
        RECT  1.785 0.360 1.855 0.600 ;
        RECT  1.340 0.995 1.760 1.065 ;
        RECT  1.580 0.185 1.700 0.265 ;
        RECT  1.565 0.700 1.635 0.920 ;
        RECT  0.485 0.195 1.580 0.265 ;
        RECT  1.495 0.335 1.565 0.770 ;
        RECT  1.410 0.850 1.450 0.920 ;
        RECT  1.340 0.345 1.410 0.920 ;
        RECT  0.930 0.345 1.340 0.415 ;
        RECT  1.110 0.850 1.340 0.920 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  0.330 0.995 1.220 1.065 ;
        RECT  0.860 0.520 0.915 0.640 ;
        RECT  0.790 0.345 0.860 0.915 ;
        RECT  0.570 0.345 0.790 0.415 ;
        RECT  0.570 0.845 0.790 0.915 ;
        RECT  0.415 0.195 0.485 0.910 ;
        RECT  0.260 0.340 0.330 1.065 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.995 0.260 1.065 ;
        RECT  0.055 0.280 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.065 ;
    END
END DFKSND2BWP

MACRO DFKSND4BWP
    CLASS CORE ;
    FOREIGN DFKSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.720 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.525 0.465 ;
        RECT  4.515 0.765 4.525 1.065 ;
        RECT  4.455 0.185 4.515 1.065 ;
        RECT  4.305 0.355 4.455 0.905 ;
        RECT  4.165 0.355 4.305 0.465 ;
        RECT  4.165 0.765 4.305 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.800 0.475 ;
        RECT  3.715 0.765 3.785 1.065 ;
        RECT  3.675 0.765 3.715 0.905 ;
        RECT  3.465 0.355 3.675 0.905 ;
        RECT  3.320 0.355 3.465 0.475 ;
        RECT  3.405 0.765 3.465 0.905 ;
        RECT  3.335 0.765 3.405 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.275 ;
        RECT  0.330 -0.115 4.250 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.680 4.710 1.375 ;
        RECT  4.345 1.145 4.630 1.375 ;
        RECT  4.275 0.975 4.345 1.375 ;
        RECT  3.975 1.145 4.275 1.375 ;
        RECT  3.905 0.745 3.975 1.375 ;
        RECT  3.595 1.145 3.905 1.375 ;
        RECT  3.525 0.975 3.595 1.375 ;
        RECT  2.050 1.145 3.525 1.375 ;
        RECT  1.930 0.845 2.050 1.375 ;
        RECT  0.330 1.145 1.930 1.375 ;
        RECT  0.210 1.030 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.355 4.235 0.465 ;
        RECT  4.165 0.765 4.235 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        RECT  3.745 0.355 3.800 0.475 ;
        RECT  3.745 0.765 3.785 1.065 ;
        RECT  3.320 0.355 3.395 0.475 ;
        RECT  3.335 0.765 3.395 1.065 ;
        RECT  3.980 0.545 4.130 0.615 ;
        RECT  3.910 0.215 3.980 0.615 ;
        RECT  2.640 0.215 3.910 0.285 ;
        RECT  3.190 0.545 3.315 0.615 ;
        RECT  3.120 0.370 3.190 1.000 ;
        RECT  2.780 0.370 3.120 0.440 ;
        RECT  2.930 0.930 3.120 1.000 ;
        RECT  2.955 0.520 3.025 0.850 ;
        RECT  2.820 0.780 2.955 0.850 ;
        RECT  2.750 0.780 2.820 1.065 ;
        RECT  2.710 0.370 2.780 0.640 ;
        RECT  2.350 0.995 2.750 1.065 ;
        RECT  2.570 0.200 2.640 0.790 ;
        RECT  2.430 0.195 2.500 0.925 ;
        RECT  2.300 0.195 2.430 0.265 ;
        RECT  2.280 0.350 2.350 1.065 ;
        RECT  2.180 0.185 2.300 0.265 ;
        RECT  2.140 0.360 2.210 1.060 ;
        RECT  1.700 0.195 2.180 0.265 ;
        RECT  1.855 0.360 2.140 0.430 ;
        RECT  2.000 0.510 2.070 0.770 ;
        RECT  1.635 0.700 2.000 0.770 ;
        RECT  1.785 0.360 1.855 0.600 ;
        RECT  1.340 0.995 1.760 1.065 ;
        RECT  1.580 0.185 1.700 0.265 ;
        RECT  1.565 0.700 1.635 0.920 ;
        RECT  0.485 0.195 1.580 0.265 ;
        RECT  1.495 0.335 1.565 0.770 ;
        RECT  1.410 0.850 1.450 0.920 ;
        RECT  1.340 0.345 1.410 0.920 ;
        RECT  0.930 0.345 1.340 0.415 ;
        RECT  1.110 0.850 1.340 0.920 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  0.620 0.995 1.220 1.065 ;
        RECT  0.860 0.520 0.915 0.640 ;
        RECT  0.790 0.345 0.860 0.905 ;
        RECT  0.570 0.345 0.790 0.415 ;
        RECT  0.570 0.835 0.790 0.905 ;
        RECT  0.500 0.995 0.620 1.075 ;
        RECT  0.480 0.995 0.500 1.065 ;
        RECT  0.415 0.185 0.485 0.810 ;
        RECT  0.410 0.890 0.480 1.065 ;
        RECT  0.330 0.890 0.410 0.960 ;
        RECT  0.260 0.340 0.330 0.960 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.890 0.260 0.960 ;
        RECT  0.055 0.270 0.125 0.410 ;
        RECT  0.055 0.890 0.125 1.040 ;
    END
END DFKSND4BWP

MACRO DFNCND1BWP
    CLASS CORE ;
    FOREIGN DFNCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.045 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.520 0.730 3.535 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.415 3.310 0.785 ;
        RECT  3.205 0.415 3.240 0.485 ;
        RECT  3.110 0.715 3.240 0.785 ;
        RECT  3.115 0.205 3.205 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.630 ;
        RECT  2.645 0.510 2.695 0.630 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 -0.115 3.640 0.115 ;
        RECT  3.320 -0.115 3.400 0.335 ;
        RECT  2.615 -0.115 3.320 0.115 ;
        RECT  2.545 -0.115 2.615 0.360 ;
        RECT  1.570 -0.115 2.545 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.145 3.640 1.375 ;
        RECT  3.300 1.010 3.420 1.375 ;
        RECT  0.690 1.145 3.300 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.450 0.520 3.460 0.640 ;
        RECT  3.380 0.520 3.450 0.935 ;
        RECT  2.910 0.865 3.380 0.935 ;
        RECT  3.005 0.555 3.150 0.625 ;
        RECT  2.935 0.230 3.005 0.775 ;
        RECT  2.510 0.705 2.935 0.775 ;
        RECT  2.840 0.845 2.910 0.935 ;
        RECT  2.770 1.005 2.880 1.075 ;
        RECT  2.370 0.845 2.840 0.915 ;
        RECT  2.700 0.985 2.770 1.075 ;
        RECT  2.230 0.985 2.700 1.055 ;
        RECT  2.440 0.520 2.510 0.775 ;
        RECT  2.410 0.520 2.440 0.640 ;
        RECT  2.340 0.375 2.430 0.445 ;
        RECT  2.340 0.700 2.370 0.915 ;
        RECT  2.300 0.375 2.340 0.915 ;
        RECT  1.710 0.200 2.330 0.270 ;
        RECT  2.270 0.375 2.300 0.770 ;
        RECT  2.130 0.375 2.270 0.445 ;
        RECT  2.175 0.830 2.230 1.055 ;
        RECT  2.160 0.660 2.175 1.055 ;
        RECT  2.105 0.660 2.160 0.900 ;
        RECT  2.045 0.660 2.105 0.730 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.350 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.195 1.370 0.430 ;
        RECT  1.160 0.195 1.300 0.265 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.840 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.770 0.845 0.840 1.055 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNCND1BWP

MACRO DFNCND2BWP
    CLASS CORE ;
    FOREIGN DFNCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.355 4.025 0.800 ;
        RECT  3.955 0.185 3.965 1.035 ;
        RECT  3.895 0.185 3.955 0.465 ;
        RECT  3.895 0.730 3.955 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 0.785 ;
        RECT  3.475 0.185 3.535 0.465 ;
        RECT  3.440 0.715 3.535 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0534 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.640 ;
        RECT  2.580 0.510 2.695 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.300 ;
        RECT  3.755 -0.115 4.070 0.115 ;
        RECT  3.685 -0.115 3.755 0.465 ;
        RECT  3.365 -0.115 3.685 0.115 ;
        RECT  3.295 -0.115 3.365 0.420 ;
        RECT  2.605 -0.115 3.295 0.115 ;
        RECT  2.535 -0.115 2.605 0.430 ;
        RECT  1.570 -0.115 2.535 0.115 ;
        RECT  1.500 -0.115 1.570 0.280 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.905 4.150 1.375 ;
        RECT  3.780 1.145 4.070 1.375 ;
        RECT  3.660 1.030 3.780 1.375 ;
        RECT  3.380 1.145 3.660 1.375 ;
        RECT  3.260 1.030 3.380 1.375 ;
        RECT  0.690 1.145 3.260 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.780 0.545 3.880 0.615 ;
        RECT  3.710 0.545 3.780 0.925 ;
        RECT  2.370 0.855 3.710 0.925 ;
        RECT  3.200 0.545 3.460 0.615 ;
        RECT  3.130 0.325 3.200 0.785 ;
        RECT  2.890 0.325 3.130 0.395 ;
        RECT  2.510 0.715 3.130 0.785 ;
        RECT  2.610 1.005 2.840 1.075 ;
        RECT  2.570 0.995 2.610 1.075 ;
        RECT  2.230 0.995 2.570 1.065 ;
        RECT  2.440 0.520 2.510 0.785 ;
        RECT  2.340 0.375 2.450 0.445 ;
        RECT  2.410 0.520 2.440 0.640 ;
        RECT  2.340 0.700 2.370 0.925 ;
        RECT  1.710 0.200 2.340 0.270 ;
        RECT  2.300 0.375 2.340 0.925 ;
        RECT  2.270 0.375 2.300 0.770 ;
        RECT  2.130 0.375 2.270 0.445 ;
        RECT  2.175 0.830 2.230 1.065 ;
        RECT  2.160 0.660 2.175 1.065 ;
        RECT  2.105 0.660 2.160 0.900 ;
        RECT  2.045 0.660 2.105 0.730 ;
        RECT  1.970 0.985 2.090 1.075 ;
        RECT  1.975 0.350 2.045 0.730 ;
        RECT  1.850 0.835 2.010 0.905 ;
        RECT  1.160 0.985 1.970 1.055 ;
        RECT  1.780 0.350 1.850 0.905 ;
        RECT  1.300 0.695 1.780 0.765 ;
        RECT  1.640 0.200 1.710 0.430 ;
        RECT  1.460 0.525 1.700 0.595 ;
        RECT  1.370 0.360 1.640 0.430 ;
        RECT  1.110 0.835 1.590 0.905 ;
        RECT  1.390 0.500 1.460 0.595 ;
        RECT  1.110 0.500 1.390 0.570 ;
        RECT  1.300 0.205 1.370 0.430 ;
        RECT  1.160 0.205 1.300 0.275 ;
        RECT  1.180 0.660 1.300 0.765 ;
        RECT  1.040 0.185 1.160 0.275 ;
        RECT  1.040 0.985 1.160 1.075 ;
        RECT  1.040 0.350 1.110 0.765 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.930 0.350 1.040 0.420 ;
        RECT  1.025 0.695 1.040 0.765 ;
        RECT  0.840 0.985 1.040 1.055 ;
        RECT  0.955 0.695 1.025 0.915 ;
        RECT  0.770 0.845 0.840 1.055 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNCND2BWP

MACRO DFNCND4BWP
    CLASS CORE ;
    FOREIGN DFNCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.665 0.485 ;
        RECT  4.655 0.765 4.665 1.065 ;
        RECT  4.595 0.185 4.655 1.065 ;
        RECT  4.445 0.355 4.595 0.905 ;
        RECT  4.310 0.355 4.445 0.485 ;
        RECT  4.305 0.765 4.445 0.905 ;
        RECT  4.240 0.185 4.310 0.485 ;
        RECT  4.235 0.765 4.305 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.705 3.960 0.785 ;
        RECT  3.855 0.185 3.925 0.475 ;
        RECT  3.815 0.355 3.855 0.475 ;
        RECT  3.605 0.355 3.815 0.785 ;
        RECT  3.545 0.355 3.605 0.475 ;
        RECT  3.440 0.705 3.605 0.785 ;
        RECT  3.475 0.185 3.545 0.475 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.630 ;
        RECT  0.735 0.355 0.805 0.630 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0526 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.640 ;
        RECT  2.615 0.510 2.695 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.115 4.900 0.115 ;
        RECT  4.770 -0.115 4.850 0.465 ;
        RECT  4.510 -0.115 4.770 0.115 ;
        RECT  4.390 -0.115 4.510 0.275 ;
        RECT  4.115 -0.115 4.390 0.115 ;
        RECT  4.045 -0.115 4.115 0.465 ;
        RECT  3.760 -0.115 4.045 0.115 ;
        RECT  3.640 -0.115 3.760 0.275 ;
        RECT  3.365 -0.115 3.640 0.115 ;
        RECT  3.295 -0.115 3.365 0.445 ;
        RECT  2.625 -0.115 3.295 0.115 ;
        RECT  2.555 -0.115 2.625 0.430 ;
        RECT  1.590 -0.115 2.555 0.115 ;
        RECT  1.520 -0.115 1.590 0.280 ;
        RECT  0.000 -0.115 1.520 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.145 4.900 1.375 ;
        RECT  4.770 0.680 4.850 1.375 ;
        RECT  4.485 1.145 4.770 1.375 ;
        RECT  4.415 0.975 4.485 1.375 ;
        RECT  4.140 1.145 4.415 1.375 ;
        RECT  4.020 1.010 4.140 1.375 ;
        RECT  3.760 1.145 4.020 1.375 ;
        RECT  3.640 1.010 3.760 1.375 ;
        RECT  3.390 1.145 3.640 1.375 ;
        RECT  3.270 1.010 3.390 1.375 ;
        RECT  0.685 1.145 3.270 1.375 ;
        RECT  0.615 0.895 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.310 0.355 4.375 0.485 ;
        RECT  4.305 0.765 4.375 0.905 ;
        RECT  4.240 0.185 4.310 0.485 ;
        RECT  4.235 0.765 4.305 1.065 ;
        RECT  3.885 0.705 3.960 0.785 ;
        RECT  3.885 0.185 3.925 0.475 ;
        RECT  3.475 0.185 3.535 0.475 ;
        RECT  3.440 0.705 3.535 0.785 ;
        RECT  4.130 0.545 4.200 0.615 ;
        RECT  4.060 0.545 4.130 0.925 ;
        RECT  2.390 0.855 4.060 0.925 ;
        RECT  3.220 0.545 3.470 0.615 ;
        RECT  3.150 0.325 3.220 0.785 ;
        RECT  2.890 0.325 3.150 0.395 ;
        RECT  2.530 0.715 3.150 0.785 ;
        RECT  2.740 0.995 2.860 1.075 ;
        RECT  2.250 0.995 2.740 1.065 ;
        RECT  2.460 0.520 2.530 0.785 ;
        RECT  2.360 0.375 2.470 0.445 ;
        RECT  2.430 0.520 2.460 0.640 ;
        RECT  2.360 0.700 2.390 0.925 ;
        RECT  1.730 0.200 2.360 0.270 ;
        RECT  2.320 0.375 2.360 0.925 ;
        RECT  2.290 0.375 2.320 0.770 ;
        RECT  2.150 0.375 2.290 0.445 ;
        RECT  2.195 0.830 2.250 1.065 ;
        RECT  2.180 0.660 2.195 1.065 ;
        RECT  2.125 0.660 2.180 0.900 ;
        RECT  2.065 0.660 2.125 0.730 ;
        RECT  1.990 0.985 2.110 1.075 ;
        RECT  1.995 0.350 2.065 0.730 ;
        RECT  1.870 0.835 2.030 0.905 ;
        RECT  1.180 0.985 1.990 1.055 ;
        RECT  1.800 0.350 1.870 0.905 ;
        RECT  1.320 0.695 1.800 0.765 ;
        RECT  1.660 0.200 1.730 0.430 ;
        RECT  1.480 0.525 1.720 0.595 ;
        RECT  1.390 0.360 1.660 0.430 ;
        RECT  1.130 0.835 1.610 0.905 ;
        RECT  1.410 0.500 1.480 0.595 ;
        RECT  1.130 0.500 1.410 0.570 ;
        RECT  1.320 0.210 1.390 0.430 ;
        RECT  1.180 0.210 1.320 0.280 ;
        RECT  1.200 0.660 1.320 0.765 ;
        RECT  1.060 0.185 1.180 0.280 ;
        RECT  1.060 0.985 1.180 1.075 ;
        RECT  1.060 0.350 1.130 0.765 ;
        RECT  0.330 0.210 1.060 0.280 ;
        RECT  0.950 0.350 1.060 0.420 ;
        RECT  1.050 0.695 1.060 0.765 ;
        RECT  0.875 0.985 1.060 1.055 ;
        RECT  0.980 0.695 1.050 0.915 ;
        RECT  0.805 0.735 0.875 1.055 ;
        RECT  0.600 0.735 0.805 0.805 ;
        RECT  0.525 0.350 0.600 0.805 ;
        RECT  0.435 0.350 0.525 0.470 ;
        RECT  0.505 0.735 0.525 0.805 ;
        RECT  0.435 0.735 0.505 1.035 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.210 0.330 0.940 ;
        RECT  0.055 0.210 0.260 0.330 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFNCND4BWP

MACRO DFNCSND1BWP
    CLASS CORE ;
    FOREIGN DFNCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.800 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.740 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0779 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.720 0.775 3.750 1.045 ;
        RECT  3.675 0.350 3.720 1.045 ;
        RECT  3.650 0.350 3.675 0.915 ;
        RECT  3.560 0.350 3.650 0.470 ;
        RECT  3.560 0.775 3.650 0.915 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.495 3.185 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.115 4.060 0.115 ;
        RECT  2.990 -0.115 3.110 0.275 ;
        RECT  1.620 -0.115 2.990 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 4.060 1.375 ;
        RECT  2.600 1.030 2.720 1.375 ;
        RECT  2.010 1.145 2.600 1.375 ;
        RECT  1.890 1.010 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.005 1.650 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.880 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.260 0.210 3.790 0.280 ;
        RECT  3.480 0.545 3.570 0.615 ;
        RECT  3.410 0.355 3.480 1.045 ;
        RECT  3.340 0.355 3.410 0.425 ;
        RECT  2.860 0.975 3.410 1.045 ;
        RECT  3.270 0.520 3.340 0.905 ;
        RECT  2.345 0.835 3.270 0.905 ;
        RECT  3.190 0.210 3.260 0.425 ;
        RECT  2.485 0.355 3.190 0.425 ;
        RECT  2.485 0.695 2.910 0.765 ;
        RECT  1.790 0.200 2.490 0.270 ;
        RECT  2.415 0.355 2.485 0.765 ;
        RECT  2.250 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.905 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.860 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.360 0.860 2.120 0.930 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  0.330 0.195 1.310 0.265 ;
        RECT  0.840 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.770 0.845 0.840 1.050 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNCSND1BWP

MACRO DFNCSND2BWP
    CLASS CORE ;
    FOREIGN DFNCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.790 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.385 0.355 4.445 0.810 ;
        RECT  4.375 0.185 4.385 1.040 ;
        RECT  4.315 0.185 4.375 0.465 ;
        RECT  4.315 0.740 4.375 1.040 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.355 4.025 1.045 ;
        RECT  3.920 0.355 3.955 0.455 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0584 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.690 0.640 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.300 ;
        RECT  3.040 -0.115 4.490 0.115 ;
        RECT  2.970 -0.115 3.040 0.270 ;
        RECT  1.620 -0.115 2.970 0.115 ;
        RECT  1.500 -0.115 1.620 0.200 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.895 4.570 1.375 ;
        RECT  4.195 1.145 4.490 1.375 ;
        RECT  4.125 0.735 4.195 1.375 ;
        RECT  3.840 1.145 4.125 1.375 ;
        RECT  3.720 1.005 3.840 1.375 ;
        RECT  3.470 1.145 3.720 1.375 ;
        RECT  3.350 1.005 3.470 1.375 ;
        RECT  3.100 1.145 3.350 1.375 ;
        RECT  2.980 1.005 3.100 1.375 ;
        RECT  2.730 1.145 2.980 1.375 ;
        RECT  2.610 1.005 2.730 1.375 ;
        RECT  2.010 1.145 2.610 1.375 ;
        RECT  1.890 1.010 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.005 1.650 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.210 0.545 4.300 0.615 ;
        RECT  4.140 0.215 4.210 0.615 ;
        RECT  3.185 0.215 4.140 0.285 ;
        RECT  3.830 0.520 3.880 0.640 ;
        RECT  3.760 0.355 3.830 0.935 ;
        RECT  3.325 0.355 3.760 0.425 ;
        RECT  3.170 0.865 3.760 0.935 ;
        RECT  3.395 0.520 3.465 0.785 ;
        RECT  3.080 0.715 3.395 0.785 ;
        RECT  3.255 0.355 3.325 0.615 ;
        RECT  2.860 0.545 3.255 0.615 ;
        RECT  3.115 0.215 3.185 0.425 ;
        RECT  2.485 0.355 3.115 0.425 ;
        RECT  3.010 0.715 3.080 0.935 ;
        RECT  2.345 0.865 3.010 0.935 ;
        RECT  2.485 0.725 2.910 0.795 ;
        RECT  2.415 0.355 2.485 0.795 ;
        RECT  1.790 0.200 2.450 0.270 ;
        RECT  2.250 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.935 ;
        RECT  2.165 0.570 2.275 0.640 ;
        RECT  1.985 0.710 2.190 0.780 ;
        RECT  2.120 0.860 2.190 1.075 ;
        RECT  2.095 0.350 2.165 0.640 ;
        RECT  1.360 0.860 2.120 0.930 ;
        RECT  1.915 0.350 1.985 0.780 ;
        RECT  1.600 0.710 1.915 0.780 ;
        RECT  1.720 0.200 1.790 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.720 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.195 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  0.330 0.195 1.310 0.265 ;
        RECT  0.840 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.770 0.845 0.840 1.050 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNCSND2BWP

MACRO DFNCSND4BWP
    CLASS CORE ;
    FOREIGN DFNCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0464 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.790 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.185 5.085 0.485 ;
        RECT  5.075 0.765 5.085 1.065 ;
        RECT  5.015 0.185 5.075 1.065 ;
        RECT  4.865 0.355 5.015 0.905 ;
        RECT  4.730 0.355 4.865 0.485 ;
        RECT  4.725 0.765 4.865 0.905 ;
        RECT  4.660 0.185 4.730 0.485 ;
        RECT  4.655 0.765 4.725 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.350 4.370 0.485 ;
        RECT  4.275 0.765 4.345 1.065 ;
        RECT  4.235 0.765 4.275 0.905 ;
        RECT  4.025 0.350 4.235 0.905 ;
        RECT  3.900 0.350 4.025 0.470 ;
        RECT  4.005 0.765 4.025 0.905 ;
        RECT  3.915 0.765 4.005 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.520 0.940 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.690 0.640 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.905 -0.115 5.190 0.115 ;
        RECT  4.835 -0.115 4.905 0.280 ;
        RECT  3.030 -0.115 4.835 0.115 ;
        RECT  2.960 -0.115 3.030 0.270 ;
        RECT  1.640 -0.115 2.960 0.115 ;
        RECT  1.520 -0.115 1.640 0.200 ;
        RECT  0.000 -0.115 1.520 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.675 5.270 1.375 ;
        RECT  4.905 1.145 5.190 1.375 ;
        RECT  4.835 0.975 4.905 1.375 ;
        RECT  4.535 1.145 4.835 1.375 ;
        RECT  4.465 0.745 4.535 1.375 ;
        RECT  4.170 1.145 4.465 1.375 ;
        RECT  4.090 0.975 4.170 1.375 ;
        RECT  3.830 1.145 4.090 1.375 ;
        RECT  3.710 1.005 3.830 1.375 ;
        RECT  3.470 1.145 3.710 1.375 ;
        RECT  3.350 1.005 3.470 1.375 ;
        RECT  3.100 1.145 3.350 1.375 ;
        RECT  2.980 1.005 3.100 1.375 ;
        RECT  2.730 1.145 2.980 1.375 ;
        RECT  2.610 1.005 2.730 1.375 ;
        RECT  2.010 1.145 2.610 1.375 ;
        RECT  1.890 1.000 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.000 1.650 1.375 ;
        RECT  0.665 1.145 1.530 1.375 ;
        RECT  0.595 0.895 0.665 1.375 ;
        RECT  0.330 1.145 0.595 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.355 4.795 0.485 ;
        RECT  4.725 0.765 4.795 0.905 ;
        RECT  4.660 0.185 4.730 0.485 ;
        RECT  4.655 0.765 4.725 1.065 ;
        RECT  4.305 0.350 4.370 0.485 ;
        RECT  4.305 0.765 4.345 1.065 ;
        RECT  3.900 0.350 3.955 0.470 ;
        RECT  3.915 0.765 3.955 1.065 ;
        RECT  4.550 0.545 4.620 0.615 ;
        RECT  4.480 0.210 4.550 0.615 ;
        RECT  3.185 0.210 4.480 0.280 ;
        RECT  3.830 0.545 3.930 0.615 ;
        RECT  3.760 0.355 3.830 0.935 ;
        RECT  3.325 0.355 3.760 0.425 ;
        RECT  3.170 0.865 3.760 0.935 ;
        RECT  3.395 0.520 3.465 0.785 ;
        RECT  3.080 0.715 3.395 0.785 ;
        RECT  3.255 0.355 3.325 0.615 ;
        RECT  2.860 0.545 3.255 0.615 ;
        RECT  3.115 0.210 3.185 0.425 ;
        RECT  2.485 0.355 3.115 0.425 ;
        RECT  3.010 0.715 3.080 0.935 ;
        RECT  2.345 0.865 3.010 0.935 ;
        RECT  2.485 0.725 2.910 0.795 ;
        RECT  1.810 0.200 2.500 0.270 ;
        RECT  2.415 0.355 2.485 0.795 ;
        RECT  2.270 0.385 2.415 0.455 ;
        RECT  2.275 0.570 2.345 0.935 ;
        RECT  2.185 0.570 2.275 0.640 ;
        RECT  2.005 0.710 2.190 0.780 ;
        RECT  2.120 0.860 2.190 1.075 ;
        RECT  2.115 0.350 2.185 0.640 ;
        RECT  1.360 0.860 2.120 0.930 ;
        RECT  1.935 0.350 2.005 0.780 ;
        RECT  1.600 0.710 1.935 0.780 ;
        RECT  1.740 0.200 1.810 0.340 ;
        RECT  1.670 0.410 1.760 0.640 ;
        RECT  1.380 0.270 1.740 0.340 ;
        RECT  1.080 0.410 1.670 0.480 ;
        RECT  1.530 0.550 1.600 0.780 ;
        RECT  1.220 0.550 1.530 0.620 ;
        RECT  1.360 0.690 1.460 0.790 ;
        RECT  1.310 0.210 1.380 0.340 ;
        RECT  1.220 0.720 1.360 0.790 ;
        RECT  1.290 0.860 1.360 1.050 ;
        RECT  1.180 0.210 1.310 0.280 ;
        RECT  0.875 0.980 1.290 1.050 ;
        RECT  1.150 0.720 1.220 0.900 ;
        RECT  1.060 0.195 1.180 0.280 ;
        RECT  1.010 0.355 1.080 0.900 ;
        RECT  0.330 0.210 1.060 0.280 ;
        RECT  0.950 0.355 1.010 0.425 ;
        RECT  0.955 0.780 1.010 0.900 ;
        RECT  0.805 0.735 0.875 1.050 ;
        RECT  0.585 0.735 0.805 0.805 ;
        RECT  0.515 0.350 0.585 0.805 ;
        RECT  0.435 0.350 0.515 0.470 ;
        RECT  0.485 0.735 0.515 0.805 ;
        RECT  0.415 0.735 0.485 1.035 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.210 0.330 0.940 ;
        RECT  0.055 0.210 0.260 0.330 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFNCSND4BWP

MACRO DFND1BWP
    CLASS CORE ;
    FOREIGN DFND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.960 0.195 3.045 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.350 2.425 0.470 ;
        RECT  2.345 0.775 2.405 0.905 ;
        RECT  2.275 0.350 2.345 0.905 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.145 3.080 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.820 0.210 2.890 0.640 ;
        RECT  2.140 0.210 2.820 0.280 ;
        RECT  2.680 0.520 2.750 1.050 ;
        RECT  2.650 0.520 2.680 0.640 ;
        RECT  1.860 0.980 2.680 1.050 ;
        RECT  2.580 0.375 2.640 0.445 ;
        RECT  2.580 0.775 2.605 0.905 ;
        RECT  2.510 0.375 2.580 0.905 ;
        RECT  2.430 0.545 2.510 0.615 ;
        RECT  2.070 0.210 2.140 0.910 ;
        RECT  1.950 0.295 2.070 0.415 ;
        RECT  1.930 0.820 2.070 0.910 ;
        RECT  1.880 0.675 1.980 0.745 ;
        RECT  1.810 0.195 1.880 0.745 ;
        RECT  1.790 0.840 1.860 1.050 ;
        RECT  1.710 0.195 1.810 0.265 ;
        RECT  1.740 0.840 1.790 0.910 ;
        RECT  1.670 0.345 1.740 0.910 ;
        RECT  1.600 0.985 1.720 1.075 ;
        RECT  1.570 0.185 1.710 0.265 ;
        RECT  1.530 0.345 1.600 0.905 ;
        RECT  0.840 0.985 1.600 1.055 ;
        RECT  1.160 0.195 1.570 0.265 ;
        RECT  1.280 0.345 1.530 0.415 ;
        RECT  1.520 0.785 1.530 0.905 ;
        RECT  1.430 0.520 1.460 0.640 ;
        RECT  1.360 0.520 1.430 0.900 ;
        RECT  1.130 0.830 1.360 0.900 ;
        RECT  1.210 0.345 1.280 0.760 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.900 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.930 0.830 1.060 0.900 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.770 0.845 0.840 1.055 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFND1BWP

MACRO DFND2BWP
    CLASS CORE ;
    FOREIGN DFND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 0.355 3.325 0.805 ;
        RECT  3.265 0.185 3.270 0.805 ;
        RECT  3.255 0.185 3.265 1.035 ;
        RECT  3.200 0.185 3.255 0.465 ;
        RECT  3.195 0.735 3.255 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.910 0.785 ;
        RECT  2.790 0.355 2.835 0.425 ;
        RECT  2.790 0.715 2.835 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.300 ;
        RECT  0.000 -0.115 3.370 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.895 3.450 1.375 ;
        RECT  3.100 1.145 3.370 1.375 ;
        RECT  2.980 1.020 3.100 1.375 ;
        RECT  2.720 1.145 2.980 1.375 ;
        RECT  2.600 1.010 2.720 1.375 ;
        RECT  0.690 1.145 2.600 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.110 0.545 3.180 0.615 ;
        RECT  3.040 0.215 3.110 0.940 ;
        RECT  2.090 0.215 3.040 0.285 ;
        RECT  2.520 0.870 3.040 0.940 ;
        RECT  2.700 0.520 2.765 0.640 ;
        RECT  2.630 0.375 2.700 0.800 ;
        RECT  2.230 0.375 2.630 0.445 ;
        RECT  2.440 0.680 2.630 0.800 ;
        RECT  2.450 0.870 2.520 1.050 ;
        RECT  1.990 0.980 2.450 1.050 ;
        RECT  2.370 0.540 2.420 0.610 ;
        RECT  2.300 0.540 2.370 0.910 ;
        RECT  1.810 0.840 2.300 0.910 ;
        RECT  2.160 0.375 2.230 0.615 ;
        RECT  2.090 0.545 2.160 0.615 ;
        RECT  2.020 0.215 2.090 0.355 ;
        RECT  1.950 0.510 1.995 0.770 ;
        RECT  1.925 0.195 1.950 0.770 ;
        RECT  1.880 0.195 1.925 0.580 ;
        RECT  1.760 0.195 1.880 0.265 ;
        RECT  1.740 0.345 1.810 0.910 ;
        RECT  1.650 0.985 1.770 1.075 ;
        RECT  1.610 0.185 1.760 0.265 ;
        RECT  0.840 0.985 1.650 1.055 ;
        RECT  1.570 0.345 1.640 0.905 ;
        RECT  1.160 0.195 1.610 0.265 ;
        RECT  1.280 0.345 1.570 0.415 ;
        RECT  1.560 0.785 1.570 0.905 ;
        RECT  1.470 0.520 1.500 0.640 ;
        RECT  1.400 0.520 1.470 0.900 ;
        RECT  1.130 0.830 1.400 0.900 ;
        RECT  1.210 0.345 1.280 0.760 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.900 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.930 0.830 1.060 0.900 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.770 0.845 0.840 1.055 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFND2BWP

MACRO DFND4BWP
    CLASS CORE ;
    FOREIGN DFND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.765 3.965 1.065 ;
        RECT  3.815 0.355 3.895 0.465 ;
        RECT  3.815 0.765 3.895 0.905 ;
        RECT  3.605 0.355 3.815 0.905 ;
        RECT  3.585 0.355 3.605 0.465 ;
        RECT  3.515 0.765 3.605 1.065 ;
        RECT  3.515 0.185 3.585 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.710 3.250 0.800 ;
        RECT  3.115 0.355 3.230 0.445 ;
        RECT  2.905 0.355 3.115 0.800 ;
        RECT  2.730 0.355 2.905 0.445 ;
        RECT  2.770 0.710 2.905 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.950 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.465 ;
        RECT  3.775 -0.115 4.070 0.115 ;
        RECT  3.705 -0.115 3.775 0.285 ;
        RECT  0.000 -0.115 3.705 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.680 4.150 1.375 ;
        RECT  3.775 1.145 4.070 1.375 ;
        RECT  3.705 0.975 3.775 1.375 ;
        RECT  3.430 1.145 3.705 1.375 ;
        RECT  3.310 1.010 3.430 1.375 ;
        RECT  3.070 1.145 3.310 1.375 ;
        RECT  2.950 1.010 3.070 1.375 ;
        RECT  2.710 1.145 2.950 1.375 ;
        RECT  2.590 1.010 2.710 1.375 ;
        RECT  0.685 1.145 2.590 1.375 ;
        RECT  0.615 0.895 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.765 3.965 1.065 ;
        RECT  3.885 0.355 3.895 0.465 ;
        RECT  3.885 0.765 3.895 0.905 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.515 0.765 3.535 1.065 ;
        RECT  3.185 0.710 3.250 0.800 ;
        RECT  3.185 0.355 3.230 0.445 ;
        RECT  2.730 0.355 2.835 0.445 ;
        RECT  2.770 0.710 2.835 0.800 ;
        RECT  3.390 0.545 3.510 0.615 ;
        RECT  3.320 0.215 3.390 0.940 ;
        RECT  2.070 0.215 3.320 0.285 ;
        RECT  2.500 0.870 3.320 0.940 ;
        RECT  2.620 0.545 2.800 0.615 ;
        RECT  2.550 0.355 2.620 0.800 ;
        RECT  2.210 0.355 2.550 0.425 ;
        RECT  2.420 0.700 2.550 0.800 ;
        RECT  2.430 0.870 2.500 1.030 ;
        RECT  2.350 0.545 2.470 0.615 ;
        RECT  1.970 0.960 2.430 1.030 ;
        RECT  2.280 0.545 2.350 0.890 ;
        RECT  1.780 0.820 2.280 0.890 ;
        RECT  2.140 0.355 2.210 0.615 ;
        RECT  2.090 0.545 2.140 0.615 ;
        RECT  2.000 0.215 2.070 0.440 ;
        RECT  1.930 0.675 2.020 0.745 ;
        RECT  1.860 0.210 1.930 0.745 ;
        RECT  1.720 0.210 1.860 0.280 ;
        RECT  1.710 0.360 1.780 0.890 ;
        RECT  1.650 0.985 1.770 1.075 ;
        RECT  1.600 0.185 1.720 0.280 ;
        RECT  0.875 0.985 1.650 1.055 ;
        RECT  1.570 0.360 1.640 0.905 ;
        RECT  1.180 0.210 1.600 0.280 ;
        RECT  1.320 0.360 1.570 0.430 ;
        RECT  1.560 0.785 1.570 0.905 ;
        RECT  1.470 0.520 1.500 0.640 ;
        RECT  1.400 0.520 1.470 0.900 ;
        RECT  1.150 0.830 1.400 0.900 ;
        RECT  1.250 0.360 1.320 0.760 ;
        RECT  1.060 0.185 1.180 0.280 ;
        RECT  1.080 0.350 1.150 0.900 ;
        RECT  0.950 0.350 1.080 0.420 ;
        RECT  0.950 0.830 1.080 0.900 ;
        RECT  0.330 0.210 1.060 0.280 ;
        RECT  0.805 0.735 0.875 1.055 ;
        RECT  0.600 0.735 0.805 0.805 ;
        RECT  0.525 0.350 0.600 0.805 ;
        RECT  0.435 0.350 0.525 0.470 ;
        RECT  0.505 0.735 0.525 0.805 ;
        RECT  0.435 0.735 0.505 1.035 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.210 0.330 0.940 ;
        RECT  0.055 0.210 0.260 0.330 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFND4BWP

MACRO DFNSND1BWP
    CLASS CORE ;
    FOREIGN DFNSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.045 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.515 0.740 3.535 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.305 0.765 3.330 1.045 ;
        RECT  3.235 0.350 3.305 1.045 ;
        RECT  3.140 0.350 3.235 0.470 ;
        RECT  3.140 0.765 3.235 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.520 0.920 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.640 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.145 3.640 1.375 ;
        RECT  2.370 1.035 2.490 1.375 ;
        RECT  1.770 1.145 2.370 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.690 1.145 1.650 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.445 0.520 3.465 0.640 ;
        RECT  3.375 0.210 3.445 0.640 ;
        RECT  2.405 0.210 3.375 0.280 ;
        RECT  3.060 0.550 3.160 0.620 ;
        RECT  2.990 0.360 3.060 1.045 ;
        RECT  2.920 0.360 2.990 0.430 ;
        RECT  2.610 0.975 2.990 1.045 ;
        RECT  2.845 0.510 2.915 0.905 ;
        RECT  2.500 0.835 2.845 0.905 ;
        RECT  2.330 0.695 2.670 0.765 ;
        RECT  2.430 0.835 2.500 0.925 ;
        RECT  2.105 0.855 2.430 0.925 ;
        RECT  2.335 0.210 2.405 0.455 ;
        RECT  2.250 0.385 2.335 0.455 ;
        RECT  2.250 0.695 2.330 0.785 ;
        RECT  1.160 0.210 2.260 0.280 ;
        RECT  2.180 0.385 2.250 0.785 ;
        RECT  2.050 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.925 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.840 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.770 0.845 0.840 1.050 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNSND1BWP

MACRO DFNSND2BWP
    CLASS CORE ;
    FOREIGN DFNSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.825 0.355 3.885 0.815 ;
        RECT  3.815 0.185 3.825 1.035 ;
        RECT  3.755 0.185 3.815 0.465 ;
        RECT  3.755 0.745 3.815 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.350 3.465 1.045 ;
        RECT  3.375 0.350 3.395 0.470 ;
        RECT  3.375 0.745 3.395 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.520 0.920 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.300 ;
        RECT  0.000 -0.115 3.930 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.905 4.010 1.375 ;
        RECT  3.635 1.145 3.930 1.375 ;
        RECT  3.565 0.735 3.635 1.375 ;
        RECT  3.285 1.145 3.565 1.375 ;
        RECT  3.160 1.010 3.285 1.375 ;
        RECT  2.910 1.145 3.160 1.375 ;
        RECT  2.790 1.010 2.910 1.375 ;
        RECT  2.490 1.145 2.790 1.375 ;
        RECT  2.370 1.035 2.490 1.375 ;
        RECT  1.770 1.145 2.370 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.690 1.145 1.650 1.375 ;
        RECT  0.570 1.005 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.670 0.545 3.740 0.615 ;
        RECT  3.600 0.210 3.670 0.615 ;
        RECT  2.405 0.210 3.600 0.280 ;
        RECT  3.260 0.520 3.325 0.640 ;
        RECT  3.190 0.365 3.260 0.940 ;
        RECT  2.775 0.365 3.190 0.435 ;
        RECT  2.960 0.870 3.190 0.940 ;
        RECT  2.925 0.520 2.995 0.800 ;
        RECT  2.860 0.730 2.925 0.800 ;
        RECT  2.790 0.730 2.860 0.940 ;
        RECT  2.105 0.870 2.790 0.940 ;
        RECT  2.705 0.365 2.775 0.640 ;
        RECT  2.250 0.730 2.670 0.800 ;
        RECT  2.335 0.210 2.405 0.455 ;
        RECT  2.250 0.385 2.335 0.455 ;
        RECT  1.160 0.210 2.260 0.280 ;
        RECT  2.180 0.385 2.250 0.800 ;
        RECT  2.050 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.940 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.840 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.330 0.195 1.040 0.265 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.770 0.845 0.840 1.050 ;
        RECT  0.575 0.845 0.770 0.915 ;
        RECT  0.505 0.340 0.575 0.915 ;
        RECT  0.415 0.340 0.505 0.460 ;
        RECT  0.415 0.795 0.505 0.915 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.195 0.330 0.970 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.850 0.260 0.970 ;
    END
END DFNSND2BWP

MACRO DFNSND4BWP
    CLASS CORE ;
    FOREIGN DFNSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.525 0.465 ;
        RECT  4.515 0.765 4.525 1.065 ;
        RECT  4.455 0.185 4.515 1.065 ;
        RECT  4.305 0.355 4.455 0.905 ;
        RECT  4.165 0.355 4.305 0.465 ;
        RECT  4.165 0.765 4.305 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.820 0.455 ;
        RECT  3.715 0.765 3.785 1.060 ;
        RECT  3.675 0.765 3.715 0.905 ;
        RECT  3.465 0.355 3.675 0.905 ;
        RECT  3.300 0.355 3.465 0.455 ;
        RECT  3.405 0.765 3.465 0.905 ;
        RECT  3.335 0.765 3.405 1.060 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.970 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.275 ;
        RECT  0.000 -0.115 4.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.675 4.710 1.375 ;
        RECT  4.345 1.145 4.630 1.375 ;
        RECT  4.275 0.975 4.345 1.375 ;
        RECT  3.975 1.145 4.275 1.375 ;
        RECT  3.905 0.735 3.975 1.375 ;
        RECT  3.610 1.145 3.905 1.375 ;
        RECT  3.510 0.985 3.610 1.375 ;
        RECT  3.240 1.145 3.510 1.375 ;
        RECT  3.120 1.010 3.240 1.375 ;
        RECT  2.870 1.145 3.120 1.375 ;
        RECT  2.750 1.010 2.870 1.375 ;
        RECT  2.510 1.145 2.750 1.375 ;
        RECT  2.390 0.990 2.510 1.375 ;
        RECT  1.790 1.145 2.390 1.375 ;
        RECT  1.670 0.990 1.790 1.375 ;
        RECT  0.685 1.145 1.670 1.375 ;
        RECT  0.615 0.895 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.355 4.235 0.465 ;
        RECT  4.165 0.765 4.235 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        RECT  3.745 0.355 3.820 0.455 ;
        RECT  3.745 0.765 3.785 1.060 ;
        RECT  3.300 0.355 3.395 0.455 ;
        RECT  3.335 0.765 3.395 1.060 ;
        RECT  3.990 0.545 4.130 0.615 ;
        RECT  3.920 0.215 3.990 0.615 ;
        RECT  2.405 0.215 3.920 0.285 ;
        RECT  3.220 0.545 3.370 0.615 ;
        RECT  3.150 0.355 3.220 0.940 ;
        RECT  2.775 0.355 3.150 0.425 ;
        RECT  2.920 0.870 3.150 0.940 ;
        RECT  2.955 0.520 3.025 0.800 ;
        RECT  2.840 0.730 2.955 0.800 ;
        RECT  2.770 0.730 2.840 0.920 ;
        RECT  2.705 0.355 2.775 0.640 ;
        RECT  2.125 0.850 2.770 0.920 ;
        RECT  2.280 0.710 2.690 0.780 ;
        RECT  2.335 0.215 2.405 0.455 ;
        RECT  2.280 0.385 2.335 0.455 ;
        RECT  2.210 0.385 2.280 0.780 ;
        RECT  1.180 0.210 2.250 0.280 ;
        RECT  2.050 0.385 2.210 0.455 ;
        RECT  2.055 0.570 2.125 0.920 ;
        RECT  1.965 0.570 2.055 0.640 ;
        RECT  1.785 0.710 1.970 0.780 ;
        RECT  1.900 0.850 1.970 1.075 ;
        RECT  1.895 0.360 1.965 0.640 ;
        RECT  1.290 0.850 1.900 0.920 ;
        RECT  1.710 0.360 1.785 0.780 ;
        RECT  1.295 0.710 1.710 0.780 ;
        RECT  1.425 0.355 1.495 0.640 ;
        RECT  1.140 0.355 1.425 0.425 ;
        RECT  1.225 0.520 1.295 0.780 ;
        RECT  1.220 0.850 1.290 1.050 ;
        RECT  0.875 0.980 1.220 1.050 ;
        RECT  1.060 0.195 1.180 0.280 ;
        RECT  1.070 0.355 1.140 0.890 ;
        RECT  0.950 0.355 1.070 0.425 ;
        RECT  0.950 0.820 1.070 0.890 ;
        RECT  0.330 0.210 1.060 0.280 ;
        RECT  0.805 0.735 0.875 1.050 ;
        RECT  0.600 0.735 0.805 0.805 ;
        RECT  0.525 0.350 0.600 0.805 ;
        RECT  0.435 0.350 0.525 0.470 ;
        RECT  0.505 0.735 0.525 0.805 ;
        RECT  0.435 0.735 0.505 1.035 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.210 0.330 0.940 ;
        RECT  0.055 0.210 0.260 0.330 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFNSND4BWP

MACRO DFQD1BWP
    CLASS CORE ;
    FOREIGN DFQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.675 0.195 2.765 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.565 -0.115 2.800 0.115 ;
        RECT  2.495 -0.115 2.565 0.325 ;
        RECT  2.205 -0.115 2.495 0.115 ;
        RECT  2.135 -0.115 2.205 0.325 ;
        RECT  0.665 -0.115 2.135 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.565 1.145 2.800 1.375 ;
        RECT  2.495 0.910 2.565 1.375 ;
        RECT  0.000 1.145 2.495 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.455 0.405 2.525 0.815 ;
        RECT  2.385 0.405 2.455 0.475 ;
        RECT  2.385 0.745 2.455 0.815 ;
        RECT  2.315 0.195 2.385 0.475 ;
        RECT  2.315 0.745 2.385 1.030 ;
        RECT  2.085 0.405 2.315 0.475 ;
        RECT  2.245 0.545 2.300 0.615 ;
        RECT  2.175 0.545 2.245 0.910 ;
        RECT  1.740 0.840 2.175 0.910 ;
        RECT  2.015 0.405 2.085 0.580 ;
        RECT  1.880 0.685 1.980 0.755 ;
        RECT  1.810 0.195 1.880 0.755 ;
        RECT  1.710 0.195 1.810 0.265 ;
        RECT  1.670 0.345 1.740 0.910 ;
        RECT  1.600 0.985 1.720 1.075 ;
        RECT  1.570 0.185 1.710 0.265 ;
        RECT  1.530 0.345 1.600 0.905 ;
        RECT  0.330 0.985 1.600 1.055 ;
        RECT  1.160 0.195 1.570 0.265 ;
        RECT  1.280 0.345 1.530 0.415 ;
        RECT  1.520 0.785 1.530 0.905 ;
        RECT  1.430 0.520 1.460 0.640 ;
        RECT  1.360 0.520 1.430 0.905 ;
        RECT  1.130 0.835 1.360 0.905 ;
        RECT  1.210 0.345 1.280 0.760 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.910 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFQD1BWP

MACRO DFQD2BWP
    CLASS CORE ;
    FOREIGN DFQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.355 2.905 0.830 ;
        RECT  2.835 0.195 2.845 1.045 ;
        RECT  2.775 0.195 2.835 0.475 ;
        RECT  2.775 0.740 2.835 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.300 ;
        RECT  2.665 -0.115 2.950 0.115 ;
        RECT  2.595 -0.115 2.665 0.325 ;
        RECT  2.285 -0.115 2.595 0.115 ;
        RECT  2.215 -0.115 2.285 0.325 ;
        RECT  0.665 -0.115 2.215 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.910 3.030 1.375 ;
        RECT  2.665 1.145 2.950 1.375 ;
        RECT  2.595 0.910 2.665 1.375 ;
        RECT  2.285 1.145 2.595 1.375 ;
        RECT  2.215 0.980 2.285 1.375 ;
        RECT  0.000 1.145 2.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.635 0.545 2.740 0.615 ;
        RECT  2.565 0.405 2.635 0.815 ;
        RECT  2.465 0.405 2.565 0.475 ;
        RECT  2.465 0.745 2.565 0.815 ;
        RECT  2.395 0.195 2.465 0.475 ;
        RECT  2.395 0.745 2.465 1.030 ;
        RECT  2.155 0.405 2.395 0.475 ;
        RECT  2.325 0.545 2.380 0.615 ;
        RECT  2.255 0.545 2.325 0.910 ;
        RECT  1.780 0.840 2.255 0.910 ;
        RECT  2.085 0.405 2.155 0.580 ;
        RECT  1.920 0.685 2.020 0.755 ;
        RECT  1.850 0.195 1.920 0.755 ;
        RECT  1.750 0.195 1.850 0.265 ;
        RECT  1.710 0.345 1.780 0.910 ;
        RECT  1.640 0.985 1.760 1.075 ;
        RECT  1.610 0.185 1.750 0.265 ;
        RECT  1.570 0.345 1.640 0.905 ;
        RECT  0.330 0.985 1.640 1.055 ;
        RECT  1.160 0.195 1.610 0.265 ;
        RECT  1.295 0.345 1.570 0.415 ;
        RECT  1.560 0.785 1.570 0.905 ;
        RECT  1.470 0.520 1.500 0.640 ;
        RECT  1.400 0.520 1.470 0.905 ;
        RECT  1.130 0.835 1.400 0.905 ;
        RECT  1.225 0.345 1.295 0.640 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.910 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.055 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFQD2BWP

MACRO DFQD4BWP
    CLASS CORE ;
    FOREIGN DFQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  3.055 0.765 3.125 1.065 ;
        RECT  2.975 0.355 3.055 0.465 ;
        RECT  2.975 0.765 3.055 0.905 ;
        RECT  2.765 0.355 2.975 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.765 2.765 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.495 0.950 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.465 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.275 ;
        RECT  2.585 -0.115 2.850 0.115 ;
        RECT  2.515 -0.115 2.585 0.315 ;
        RECT  2.225 -0.115 2.515 0.115 ;
        RECT  2.155 -0.115 2.225 0.315 ;
        RECT  0.665 -0.115 2.155 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.675 3.310 1.375 ;
        RECT  2.945 1.145 3.230 1.375 ;
        RECT  2.875 0.975 2.945 1.375 ;
        RECT  2.610 1.145 2.875 1.375 ;
        RECT  2.490 1.010 2.610 1.375 ;
        RECT  0.690 1.145 2.490 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.055 0.185 3.125 0.465 ;
        RECT  3.055 0.765 3.125 1.065 ;
        RECT  3.045 0.355 3.055 0.465 ;
        RECT  3.045 0.765 3.055 0.905 ;
        RECT  2.540 0.520 2.650 0.640 ;
        RECT  2.470 0.395 2.540 0.940 ;
        RECT  2.405 0.395 2.470 0.465 ;
        RECT  2.300 0.870 2.470 0.940 ;
        RECT  2.335 0.185 2.405 0.465 ;
        RECT  2.310 0.545 2.360 0.615 ;
        RECT  2.155 0.395 2.335 0.465 ;
        RECT  2.240 0.545 2.310 0.800 ;
        RECT  2.180 0.730 2.240 0.800 ;
        RECT  2.110 0.730 2.180 0.890 ;
        RECT  2.085 0.395 2.155 0.640 ;
        RECT  1.790 0.820 2.110 0.890 ;
        RECT  1.930 0.675 2.000 0.745 ;
        RECT  1.860 0.195 1.930 0.745 ;
        RECT  1.740 0.195 1.860 0.265 ;
        RECT  1.720 0.345 1.790 0.890 ;
        RECT  1.630 0.985 1.750 1.075 ;
        RECT  1.590 0.185 1.740 0.265 ;
        RECT  0.850 0.985 1.630 1.055 ;
        RECT  1.550 0.345 1.620 0.905 ;
        RECT  1.160 0.195 1.590 0.265 ;
        RECT  1.295 0.345 1.550 0.415 ;
        RECT  1.540 0.785 1.550 0.905 ;
        RECT  1.450 0.520 1.480 0.640 ;
        RECT  1.380 0.520 1.450 0.905 ;
        RECT  1.130 0.835 1.380 0.905 ;
        RECT  1.225 0.345 1.295 0.640 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.060 0.350 1.130 0.905 ;
        RECT  0.930 0.350 1.060 0.420 ;
        RECT  0.930 0.835 1.060 0.905 ;
        RECT  0.830 0.195 1.040 0.265 ;
        RECT  0.780 0.870 0.850 1.055 ;
        RECT  0.760 0.195 0.830 0.410 ;
        RECT  0.330 0.870 0.780 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.475 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.475 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFQD4BWP

MACRO DFSND1BWP
    CLASS CORE ;
    FOREIGN DFSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.605 1.045 ;
        RECT  3.515 0.185 3.535 0.465 ;
        RECT  3.515 0.740 3.535 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.305 0.765 3.330 1.045 ;
        RECT  3.235 0.350 3.305 1.045 ;
        RECT  3.140 0.350 3.235 0.470 ;
        RECT  3.140 0.765 3.235 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.665 -0.115 3.640 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 3.640 1.375 ;
        RECT  2.360 1.010 2.480 1.375 ;
        RECT  1.770 1.145 2.360 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.000 1.145 1.650 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.445 0.520 3.465 0.640 ;
        RECT  3.375 0.210 3.445 0.640 ;
        RECT  2.405 0.210 3.375 0.280 ;
        RECT  3.060 0.550 3.160 0.620 ;
        RECT  2.990 0.360 3.060 1.045 ;
        RECT  2.920 0.360 2.990 0.430 ;
        RECT  2.610 0.975 2.990 1.045 ;
        RECT  2.845 0.510 2.915 0.905 ;
        RECT  2.500 0.835 2.845 0.905 ;
        RECT  2.330 0.695 2.670 0.765 ;
        RECT  2.430 0.835 2.500 0.925 ;
        RECT  2.105 0.855 2.430 0.925 ;
        RECT  2.335 0.210 2.405 0.455 ;
        RECT  2.250 0.385 2.335 0.455 ;
        RECT  2.250 0.695 2.330 0.785 ;
        RECT  1.160 0.210 2.260 0.280 ;
        RECT  2.180 0.385 2.250 0.785 ;
        RECT  2.050 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.925 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.330 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFSND1BWP

MACRO DFSND2BWP
    CLASS CORE ;
    FOREIGN DFSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0460 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.825 0.355 3.885 0.815 ;
        RECT  3.815 0.185 3.825 1.035 ;
        RECT  3.755 0.185 3.815 0.465 ;
        RECT  3.755 0.745 3.815 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.350 3.465 1.045 ;
        RECT  3.375 0.350 3.395 0.470 ;
        RECT  3.375 0.745 3.395 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.300 ;
        RECT  0.665 -0.115 3.930 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.905 4.010 1.375 ;
        RECT  3.635 1.145 3.930 1.375 ;
        RECT  3.565 0.735 3.635 1.375 ;
        RECT  2.910 1.145 3.565 1.375 ;
        RECT  2.790 1.010 2.910 1.375 ;
        RECT  2.490 1.145 2.790 1.375 ;
        RECT  2.370 1.035 2.490 1.375 ;
        RECT  1.770 1.145 2.370 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.000 1.145 1.650 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.670 0.545 3.740 0.615 ;
        RECT  3.600 0.210 3.670 0.615 ;
        RECT  2.405 0.210 3.600 0.280 ;
        RECT  3.260 0.520 3.325 0.640 ;
        RECT  3.190 0.365 3.260 0.940 ;
        RECT  2.775 0.365 3.190 0.435 ;
        RECT  2.960 0.870 3.190 0.940 ;
        RECT  2.925 0.520 2.995 0.800 ;
        RECT  2.860 0.730 2.925 0.800 ;
        RECT  2.790 0.730 2.860 0.940 ;
        RECT  2.105 0.870 2.790 0.940 ;
        RECT  2.705 0.365 2.775 0.640 ;
        RECT  2.250 0.730 2.670 0.800 ;
        RECT  2.335 0.210 2.405 0.455 ;
        RECT  2.250 0.385 2.335 0.455 ;
        RECT  1.160 0.210 2.260 0.280 ;
        RECT  2.180 0.385 2.250 0.800 ;
        RECT  2.050 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.940 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.330 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFSND2BWP

MACRO DFSND4BWP
    CLASS CORE ;
    FOREIGN DFSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.625 ;
        RECT  2.430 0.540 2.555 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.525 0.465 ;
        RECT  4.515 0.765 4.525 1.065 ;
        RECT  4.455 0.185 4.515 1.065 ;
        RECT  4.305 0.355 4.455 0.905 ;
        RECT  4.165 0.355 4.305 0.465 ;
        RECT  4.165 0.765 4.305 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.820 0.455 ;
        RECT  3.715 0.765 3.785 1.060 ;
        RECT  3.675 0.765 3.715 0.905 ;
        RECT  3.465 0.355 3.675 0.905 ;
        RECT  3.300 0.355 3.465 0.455 ;
        RECT  3.405 0.765 3.465 0.905 ;
        RECT  3.335 0.765 3.405 1.060 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.275 ;
        RECT  0.665 -0.115 4.250 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.675 4.710 1.375 ;
        RECT  4.345 1.145 4.630 1.375 ;
        RECT  4.275 0.975 4.345 1.375 ;
        RECT  3.975 1.145 4.275 1.375 ;
        RECT  3.905 0.735 3.975 1.375 ;
        RECT  3.610 1.145 3.905 1.375 ;
        RECT  3.510 0.985 3.610 1.375 ;
        RECT  3.240 1.145 3.510 1.375 ;
        RECT  3.120 1.010 3.240 1.375 ;
        RECT  2.870 1.145 3.120 1.375 ;
        RECT  2.750 1.010 2.870 1.375 ;
        RECT  2.510 1.145 2.750 1.375 ;
        RECT  2.390 0.990 2.510 1.375 ;
        RECT  1.770 1.145 2.390 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.690 1.145 1.650 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.355 4.235 0.465 ;
        RECT  4.165 0.765 4.235 0.905 ;
        RECT  4.095 0.185 4.165 0.465 ;
        RECT  4.095 0.765 4.165 1.065 ;
        RECT  3.745 0.355 3.820 0.455 ;
        RECT  3.745 0.765 3.785 1.060 ;
        RECT  3.300 0.355 3.395 0.455 ;
        RECT  3.335 0.765 3.395 1.060 ;
        RECT  3.990 0.545 4.130 0.615 ;
        RECT  3.920 0.215 3.990 0.615 ;
        RECT  2.405 0.215 3.920 0.285 ;
        RECT  3.220 0.545 3.370 0.615 ;
        RECT  3.150 0.355 3.220 0.940 ;
        RECT  2.775 0.355 3.150 0.425 ;
        RECT  2.920 0.870 3.150 0.940 ;
        RECT  2.955 0.520 3.025 0.800 ;
        RECT  2.840 0.730 2.955 0.800 ;
        RECT  2.770 0.730 2.840 0.920 ;
        RECT  2.705 0.355 2.775 0.640 ;
        RECT  2.105 0.850 2.770 0.920 ;
        RECT  2.250 0.710 2.690 0.780 ;
        RECT  2.335 0.215 2.405 0.455 ;
        RECT  2.250 0.385 2.335 0.455 ;
        RECT  2.180 0.385 2.250 0.780 ;
        RECT  1.160 0.210 2.240 0.280 ;
        RECT  2.050 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.920 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.860 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.790 0.870 0.860 1.050 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.330 0.870 0.790 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.475 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.475 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFSND4BWP

MACRO DFSNQD1BWP
    CLASS CORE ;
    FOREIGN DFSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.485 0.630 ;
        RECT  2.320 0.530 2.415 0.630 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.185 3.325 1.045 ;
        RECT  3.235 0.185 3.255 0.465 ;
        RECT  3.235 0.740 3.255 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.115 3.360 0.115 ;
        RECT  3.020 -0.115 3.140 0.270 ;
        RECT  0.665 -0.115 3.020 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 1.145 3.360 1.375 ;
        RECT  3.020 1.120 3.140 1.375 ;
        RECT  1.770 1.145 3.020 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.000 1.145 1.650 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.135 0.520 3.180 0.640 ;
        RECT  3.065 0.370 3.135 1.050 ;
        RECT  2.925 0.370 3.065 0.440 ;
        RECT  2.830 0.980 3.065 1.050 ;
        RECT  2.925 0.520 2.995 0.910 ;
        RECT  2.855 0.185 2.925 0.440 ;
        RECT  2.105 0.840 2.925 0.910 ;
        RECT  2.645 0.370 2.855 0.440 ;
        RECT  2.245 0.700 2.690 0.770 ;
        RECT  2.575 0.370 2.645 0.615 ;
        RECT  2.245 0.365 2.330 0.435 ;
        RECT  2.175 0.365 2.245 0.770 ;
        RECT  1.160 0.210 2.220 0.280 ;
        RECT  2.030 0.385 2.175 0.455 ;
        RECT  2.035 0.570 2.105 0.910 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.330 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFSNQD1BWP

MACRO DFSNQD2BWP
    CLASS CORE ;
    FOREIGN DFSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.485 0.640 ;
        RECT  2.320 0.545 2.415 0.640 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.265 0.355 3.325 0.815 ;
        RECT  3.255 0.185 3.265 1.030 ;
        RECT  3.195 0.185 3.255 0.465 ;
        RECT  3.195 0.735 3.255 1.030 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.300 ;
        RECT  3.110 -0.115 3.370 0.115 ;
        RECT  2.990 -0.115 3.110 0.280 ;
        RECT  2.750 -0.115 2.990 0.115 ;
        RECT  2.630 -0.115 2.750 0.280 ;
        RECT  0.665 -0.115 2.630 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.905 3.450 1.375 ;
        RECT  3.110 1.145 3.370 1.375 ;
        RECT  2.990 1.010 3.110 1.375 ;
        RECT  2.740 1.145 2.990 1.375 ;
        RECT  2.620 1.005 2.740 1.375 ;
        RECT  2.310 1.145 2.620 1.375 ;
        RECT  2.190 0.995 2.310 1.375 ;
        RECT  1.770 1.145 2.190 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.000 1.145 1.650 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.100 0.520 3.150 0.640 ;
        RECT  3.030 0.370 3.100 0.940 ;
        RECT  2.905 0.370 3.030 0.440 ;
        RECT  2.800 0.870 3.030 0.940 ;
        RECT  2.835 0.185 2.905 0.440 ;
        RECT  2.635 0.370 2.835 0.440 ;
        RECT  2.765 0.520 2.835 0.800 ;
        RECT  2.710 0.730 2.765 0.800 ;
        RECT  2.640 0.730 2.710 0.925 ;
        RECT  2.105 0.855 2.640 0.925 ;
        RECT  2.565 0.370 2.635 0.640 ;
        RECT  2.250 0.715 2.530 0.785 ;
        RECT  2.250 0.360 2.340 0.460 ;
        RECT  2.180 0.360 2.250 0.785 ;
        RECT  1.160 0.210 2.220 0.280 ;
        RECT  2.030 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.925 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.330 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.890 ;
        RECT  0.415 0.340 0.515 0.460 ;
        RECT  0.415 0.770 0.515 0.890 ;
        RECT  0.330 0.520 0.375 0.640 ;
        RECT  0.260 0.275 0.330 1.050 ;
        RECT  0.055 0.275 0.260 0.395 ;
        RECT  0.055 0.865 0.260 0.985 ;
    END
END DFSNQD2BWP

MACRO DFSNQD4BWP
    CLASS CORE ;
    FOREIGN DFSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.485 0.640 ;
        RECT  2.340 0.545 2.415 0.640 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.185 3.685 0.465 ;
        RECT  3.675 0.765 3.685 1.060 ;
        RECT  3.615 0.185 3.675 1.060 ;
        RECT  3.465 0.355 3.615 0.905 ;
        RECT  3.325 0.355 3.465 0.465 ;
        RECT  3.325 0.765 3.465 0.905 ;
        RECT  3.255 0.185 3.325 0.465 ;
        RECT  3.255 0.765 3.325 1.060 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.925 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.490 0.190 0.640 ;
        RECT  0.035 0.490 0.105 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.465 ;
        RECT  3.530 -0.115 3.790 0.115 ;
        RECT  3.410 -0.115 3.530 0.275 ;
        RECT  3.170 -0.115 3.410 0.115 ;
        RECT  3.050 -0.115 3.170 0.280 ;
        RECT  2.810 -0.115 3.050 0.115 ;
        RECT  2.690 -0.115 2.810 0.280 ;
        RECT  0.665 -0.115 2.690 0.115 ;
        RECT  0.595 -0.115 0.665 0.270 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.675 3.870 1.375 ;
        RECT  3.520 1.145 3.790 1.375 ;
        RECT  3.420 0.985 3.520 1.375 ;
        RECT  3.170 1.145 3.420 1.375 ;
        RECT  3.050 1.010 3.170 1.375 ;
        RECT  2.780 1.145 3.050 1.375 ;
        RECT  2.660 1.005 2.780 1.375 ;
        RECT  2.330 1.145 2.660 1.375 ;
        RECT  2.210 0.995 2.330 1.375 ;
        RECT  1.770 1.145 2.210 1.375 ;
        RECT  1.650 0.990 1.770 1.375 ;
        RECT  0.690 1.145 1.650 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.325 0.355 3.395 0.465 ;
        RECT  3.325 0.765 3.395 0.905 ;
        RECT  3.255 0.185 3.325 0.465 ;
        RECT  3.255 0.765 3.325 1.060 ;
        RECT  3.160 0.545 3.265 0.615 ;
        RECT  3.090 0.370 3.160 0.940 ;
        RECT  2.965 0.370 3.090 0.440 ;
        RECT  2.860 0.870 3.090 0.940 ;
        RECT  2.895 0.185 2.965 0.440 ;
        RECT  2.835 0.520 2.905 0.800 ;
        RECT  2.655 0.370 2.895 0.440 ;
        RECT  2.730 0.730 2.835 0.800 ;
        RECT  2.660 0.730 2.730 0.925 ;
        RECT  2.105 0.855 2.660 0.925 ;
        RECT  2.585 0.370 2.655 0.640 ;
        RECT  2.250 0.715 2.550 0.785 ;
        RECT  2.250 0.350 2.345 0.470 ;
        RECT  2.180 0.350 2.250 0.785 ;
        RECT  1.160 0.210 2.240 0.280 ;
        RECT  2.030 0.385 2.180 0.455 ;
        RECT  2.035 0.570 2.105 0.925 ;
        RECT  1.945 0.570 2.035 0.640 ;
        RECT  1.765 0.710 1.950 0.780 ;
        RECT  1.880 0.850 1.950 1.075 ;
        RECT  1.875 0.360 1.945 0.640 ;
        RECT  1.270 0.850 1.880 0.920 ;
        RECT  1.695 0.360 1.765 0.780 ;
        RECT  1.275 0.710 1.695 0.780 ;
        RECT  1.405 0.355 1.475 0.640 ;
        RECT  1.080 0.355 1.405 0.425 ;
        RECT  1.205 0.520 1.275 0.780 ;
        RECT  1.200 0.850 1.270 1.050 ;
        RECT  0.860 0.980 1.200 1.050 ;
        RECT  1.040 0.195 1.160 0.280 ;
        RECT  1.010 0.355 1.080 0.885 ;
        RECT  0.830 0.210 1.040 0.280 ;
        RECT  0.930 0.355 1.010 0.425 ;
        RECT  0.930 0.815 1.010 0.885 ;
        RECT  0.790 0.870 0.860 1.050 ;
        RECT  0.760 0.210 0.830 0.410 ;
        RECT  0.330 0.870 0.790 0.940 ;
        RECT  0.585 0.340 0.760 0.410 ;
        RECT  0.515 0.340 0.585 0.800 ;
        RECT  0.485 0.340 0.515 0.475 ;
        RECT  0.400 0.700 0.515 0.800 ;
        RECT  0.415 0.185 0.485 0.475 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.340 0.330 0.940 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.125 0.870 0.260 0.940 ;
        RECT  0.055 0.250 0.125 0.410 ;
        RECT  0.055 0.870 0.125 1.040 ;
    END
END DFSNQD4BWP

MACRO DFXD1BWP
    CLASS CORE ;
    FOREIGN DFXD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.740 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.645 0.340 3.715 0.810 ;
        RECT  3.520 0.340 3.645 0.460 ;
        RECT  3.605 0.730 3.645 0.810 ;
        RECT  3.520 0.730 3.605 1.045 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 -0.115 4.060 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.795 1.145 4.060 1.375 ;
        RECT  3.725 0.890 3.795 1.375 ;
        RECT  2.380 1.145 3.725 1.375 ;
        RECT  2.260 0.865 2.380 1.375 ;
        RECT  0.330 1.145 2.260 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.855 0.520 3.880 0.640 ;
        RECT  3.785 0.195 3.855 0.640 ;
        RECT  3.000 0.195 3.785 0.265 ;
        RECT  3.450 0.545 3.575 0.615 ;
        RECT  3.380 0.365 3.450 0.975 ;
        RECT  3.140 0.365 3.380 0.435 ;
        RECT  3.310 0.905 3.380 0.975 ;
        RECT  3.240 0.520 3.310 0.800 ;
        RECT  3.210 0.730 3.240 0.800 ;
        RECT  3.140 0.730 3.210 1.050 ;
        RECT  3.070 0.365 3.140 0.640 ;
        RECT  2.710 0.980 3.140 1.050 ;
        RECT  3.000 0.805 3.060 0.875 ;
        RECT  2.930 0.195 3.000 0.875 ;
        RECT  2.790 0.195 2.860 0.900 ;
        RECT  2.680 0.195 2.790 0.265 ;
        RECT  2.780 0.780 2.790 0.900 ;
        RECT  2.710 0.350 2.720 0.470 ;
        RECT  2.640 0.350 2.710 1.050 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.545 0.340 2.570 0.790 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.500 0.340 2.545 1.020 ;
        RECT  2.480 0.340 2.500 0.460 ;
        RECT  2.475 0.720 2.500 1.020 ;
        RECT  2.255 0.720 2.475 0.790 ;
        RECT  2.405 0.510 2.430 0.630 ;
        RECT  2.335 0.375 2.405 0.630 ;
        RECT  2.060 0.375 2.335 0.445 ;
        RECT  2.185 0.520 2.255 0.790 ;
        RECT  1.990 0.375 2.060 0.795 ;
        RECT  1.910 0.375 1.990 0.445 ;
        RECT  1.965 0.725 1.990 0.795 ;
        RECT  1.895 0.725 1.965 0.970 ;
        RECT  1.790 0.575 1.910 0.645 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.570 0.865 1.810 0.935 ;
        RECT  1.720 0.350 1.790 0.795 ;
        RECT  1.520 0.350 1.720 0.420 ;
        RECT  1.500 0.725 1.720 0.795 ;
        RECT  1.500 0.865 1.570 1.055 ;
        RECT  1.410 0.545 1.540 0.615 ;
        RECT  0.685 0.985 1.500 1.055 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.140 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.755 0.350 0.830 0.915 ;
        RECT  0.615 0.810 0.685 1.055 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXD1BWP

MACRO DFXD2BWP
    CLASS CORE ;
    FOREIGN DFXD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.805 ;
        RECT  4.235 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.235 0.465 ;
        RECT  4.175 0.735 4.235 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.350 3.885 1.045 ;
        RECT  3.795 0.350 3.815 0.470 ;
        RECT  3.795 0.735 3.815 1.045 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.300 ;
        RECT  0.330 -0.115 4.350 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.895 4.430 1.375 ;
        RECT  4.055 1.145 4.350 1.375 ;
        RECT  3.985 0.735 4.055 1.375 ;
        RECT  2.420 1.145 3.985 1.375 ;
        RECT  2.300 0.865 2.420 1.375 ;
        RECT  0.330 1.145 2.300 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.080 0.545 4.160 0.615 ;
        RECT  4.010 0.210 4.080 0.615 ;
        RECT  3.100 0.210 4.010 0.280 ;
        RECT  3.660 0.520 3.745 0.640 ;
        RECT  3.590 0.365 3.660 1.000 ;
        RECT  3.240 0.365 3.590 0.435 ;
        RECT  3.390 0.930 3.590 1.000 ;
        RECT  3.345 0.520 3.415 0.790 ;
        RECT  3.310 0.720 3.345 0.790 ;
        RECT  3.240 0.720 3.310 1.050 ;
        RECT  3.170 0.365 3.240 0.640 ;
        RECT  2.790 0.980 3.240 1.050 ;
        RECT  3.030 0.185 3.100 0.820 ;
        RECT  2.870 0.195 2.940 0.910 ;
        RECT  2.760 0.195 2.870 0.265 ;
        RECT  2.790 0.350 2.800 0.470 ;
        RECT  2.720 0.350 2.790 1.050 ;
        RECT  2.640 0.185 2.760 0.265 ;
        RECT  2.625 0.340 2.650 0.790 ;
        RECT  2.030 0.195 2.640 0.265 ;
        RECT  2.580 0.340 2.625 1.020 ;
        RECT  2.560 0.340 2.580 0.460 ;
        RECT  2.555 0.720 2.580 1.020 ;
        RECT  2.275 0.720 2.555 0.790 ;
        RECT  2.485 0.510 2.510 0.630 ;
        RECT  2.415 0.375 2.485 0.630 ;
        RECT  2.125 0.375 2.415 0.445 ;
        RECT  2.205 0.520 2.275 0.790 ;
        RECT  2.055 0.375 2.125 0.795 ;
        RECT  1.930 0.375 2.055 0.445 ;
        RECT  1.985 0.725 2.055 0.795 ;
        RECT  1.915 0.725 1.985 0.970 ;
        RECT  1.810 0.575 1.950 0.645 ;
        RECT  0.610 0.195 1.860 0.265 ;
        RECT  1.590 0.865 1.830 0.935 ;
        RECT  1.740 0.350 1.810 0.795 ;
        RECT  1.540 0.350 1.740 0.420 ;
        RECT  1.520 0.725 1.740 0.795 ;
        RECT  1.520 0.865 1.590 1.055 ;
        RECT  1.410 0.545 1.560 0.615 ;
        RECT  0.685 0.985 1.520 1.055 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.140 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.755 0.350 0.830 0.915 ;
        RECT  0.615 0.810 0.685 1.055 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXD2BWP

MACRO DFXD4BWP
    CLASS CORE ;
    FOREIGN DFXD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 4.945 0.465 ;
        RECT  4.935 0.765 4.945 1.065 ;
        RECT  4.875 0.185 4.935 1.065 ;
        RECT  4.725 0.355 4.875 0.905 ;
        RECT  4.585 0.355 4.725 0.465 ;
        RECT  4.585 0.765 4.725 0.905 ;
        RECT  4.515 0.185 4.585 0.465 ;
        RECT  4.515 0.765 4.585 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.355 4.230 0.455 ;
        RECT  4.135 0.765 4.205 1.065 ;
        RECT  4.095 0.765 4.135 0.905 ;
        RECT  3.885 0.355 4.095 0.905 ;
        RECT  3.730 0.355 3.885 0.455 ;
        RECT  3.825 0.765 3.885 0.905 ;
        RECT  3.755 0.765 3.825 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.465 ;
        RECT  4.790 -0.115 5.050 0.115 ;
        RECT  4.670 -0.115 4.790 0.275 ;
        RECT  0.330 -0.115 4.670 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.145 5.180 1.375 ;
        RECT  5.050 0.675 5.130 1.375 ;
        RECT  4.765 1.145 5.050 1.375 ;
        RECT  4.695 0.975 4.765 1.375 ;
        RECT  4.395 1.145 4.695 1.375 ;
        RECT  4.325 0.735 4.395 1.375 ;
        RECT  4.030 1.145 4.325 1.375 ;
        RECT  3.930 0.985 4.030 1.375 ;
        RECT  3.660 1.145 3.930 1.375 ;
        RECT  3.540 1.030 3.660 1.375 ;
        RECT  3.280 1.145 3.540 1.375 ;
        RECT  3.160 1.010 3.280 1.375 ;
        RECT  2.400 1.145 3.160 1.375 ;
        RECT  2.280 0.865 2.400 1.375 ;
        RECT  0.330 1.145 2.280 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.355 4.655 0.465 ;
        RECT  4.585 0.765 4.655 0.905 ;
        RECT  4.515 0.185 4.585 0.465 ;
        RECT  4.515 0.765 4.585 1.065 ;
        RECT  4.165 0.355 4.230 0.455 ;
        RECT  4.165 0.765 4.205 1.065 ;
        RECT  3.730 0.355 3.815 0.455 ;
        RECT  3.755 0.765 3.815 1.065 ;
        RECT  4.400 0.545 4.560 0.615 ;
        RECT  4.330 0.215 4.400 0.615 ;
        RECT  3.055 0.215 4.330 0.285 ;
        RECT  3.630 0.545 3.760 0.615 ;
        RECT  3.560 0.355 3.630 0.960 ;
        RECT  3.195 0.355 3.560 0.425 ;
        RECT  3.350 0.890 3.560 0.960 ;
        RECT  3.375 0.520 3.445 0.815 ;
        RECT  3.270 0.745 3.375 0.815 ;
        RECT  3.200 0.745 3.270 0.940 ;
        RECT  3.080 0.870 3.200 0.940 ;
        RECT  3.125 0.355 3.195 0.640 ;
        RECT  3.010 0.870 3.080 1.060 ;
        RECT  2.985 0.185 3.055 0.800 ;
        RECT  2.750 0.990 3.010 1.060 ;
        RECT  2.830 0.195 2.900 0.910 ;
        RECT  2.720 0.195 2.830 0.265 ;
        RECT  2.820 0.790 2.830 0.910 ;
        RECT  2.750 0.350 2.760 0.470 ;
        RECT  2.680 0.350 2.750 1.060 ;
        RECT  2.600 0.185 2.720 0.265 ;
        RECT  2.575 0.340 2.610 0.790 ;
        RECT  2.030 0.195 2.600 0.265 ;
        RECT  2.540 0.340 2.575 1.020 ;
        RECT  2.520 0.340 2.540 0.460 ;
        RECT  2.505 0.720 2.540 1.020 ;
        RECT  2.275 0.720 2.505 0.790 ;
        RECT  2.445 0.510 2.470 0.630 ;
        RECT  2.375 0.375 2.445 0.630 ;
        RECT  2.125 0.375 2.375 0.445 ;
        RECT  2.205 0.520 2.275 0.790 ;
        RECT  2.055 0.375 2.125 0.795 ;
        RECT  1.930 0.375 2.055 0.445 ;
        RECT  2.005 0.725 2.055 0.795 ;
        RECT  1.935 0.725 2.005 0.970 ;
        RECT  1.810 0.575 1.970 0.645 ;
        RECT  0.610 0.210 1.860 0.280 ;
        RECT  1.590 0.865 1.850 0.935 ;
        RECT  1.740 0.350 1.810 0.795 ;
        RECT  1.540 0.350 1.740 0.420 ;
        RECT  1.540 0.725 1.740 0.795 ;
        RECT  1.520 0.865 1.590 1.045 ;
        RECT  1.410 0.545 1.560 0.615 ;
        RECT  0.685 0.975 1.520 1.045 ;
        RECT  1.340 0.350 1.410 0.905 ;
        RECT  1.170 0.350 1.340 0.420 ;
        RECT  1.140 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.835 0.900 0.905 ;
        RECT  0.755 0.350 0.830 0.905 ;
        RECT  0.615 0.810 0.685 1.045 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXD4BWP

MACRO DFXQD1BWP
    CLASS CORE ;
    FOREIGN DFXQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.185 3.745 1.045 ;
        RECT  3.655 0.185 3.675 0.465 ;
        RECT  3.655 0.740 3.675 1.045 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 -0.115 3.780 0.115 ;
        RECT  3.440 -0.115 3.560 0.275 ;
        RECT  0.330 -0.115 3.440 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 1.145 3.780 1.375 ;
        RECT  3.095 0.940 3.165 1.375 ;
        RECT  2.380 1.145 3.095 1.375 ;
        RECT  2.260 0.865 2.380 1.375 ;
        RECT  0.330 1.145 2.260 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.585 0.520 3.600 0.640 ;
        RECT  3.515 0.370 3.585 0.995 ;
        RECT  3.345 0.370 3.515 0.440 ;
        RECT  3.250 0.925 3.515 0.995 ;
        RECT  3.345 0.520 3.415 0.830 ;
        RECT  3.275 0.185 3.345 0.440 ;
        RECT  3.010 0.760 3.345 0.830 ;
        RECT  3.055 0.370 3.275 0.440 ;
        RECT  2.985 0.370 3.055 0.640 ;
        RECT  2.940 0.760 3.010 1.050 ;
        RECT  2.720 0.980 2.940 1.050 ;
        RECT  2.790 0.195 2.860 0.900 ;
        RECT  2.680 0.195 2.790 0.265 ;
        RECT  2.650 0.350 2.720 1.050 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.545 0.340 2.570 0.790 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.500 0.340 2.545 1.020 ;
        RECT  2.480 0.340 2.500 0.460 ;
        RECT  2.475 0.720 2.500 1.020 ;
        RECT  2.255 0.720 2.475 0.790 ;
        RECT  2.405 0.510 2.430 0.630 ;
        RECT  2.335 0.375 2.405 0.630 ;
        RECT  2.060 0.375 2.335 0.445 ;
        RECT  2.185 0.520 2.255 0.790 ;
        RECT  1.990 0.375 2.060 0.795 ;
        RECT  1.910 0.375 1.990 0.445 ;
        RECT  1.965 0.725 1.990 0.795 ;
        RECT  1.895 0.725 1.965 0.970 ;
        RECT  1.790 0.575 1.910 0.645 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.570 0.865 1.810 0.935 ;
        RECT  1.720 0.350 1.790 0.795 ;
        RECT  1.520 0.350 1.720 0.420 ;
        RECT  1.500 0.725 1.720 0.795 ;
        RECT  1.500 0.865 1.570 1.055 ;
        RECT  1.410 0.545 1.540 0.615 ;
        RECT  0.685 0.985 1.500 1.055 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.140 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.755 0.350 0.830 0.915 ;
        RECT  0.615 0.810 0.685 1.055 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXQD1BWP

MACRO DFXQD2BWP
    CLASS CORE ;
    FOREIGN DFXQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.685 0.355 3.745 0.805 ;
        RECT  3.675 0.185 3.685 1.035 ;
        RECT  3.615 0.185 3.675 0.465 ;
        RECT  3.615 0.735 3.675 1.035 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.300 ;
        RECT  3.530 -0.115 3.790 0.115 ;
        RECT  3.410 -0.115 3.530 0.270 ;
        RECT  3.170 -0.115 3.410 0.115 ;
        RECT  3.050 -0.115 3.170 0.280 ;
        RECT  0.330 -0.115 3.050 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.895 3.870 1.375 ;
        RECT  3.150 1.145 3.790 1.375 ;
        RECT  3.080 0.945 3.150 1.375 ;
        RECT  2.380 1.145 3.080 1.375 ;
        RECT  2.260 0.865 2.380 1.375 ;
        RECT  0.330 1.145 2.260 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.480 0.520 3.570 0.640 ;
        RECT  3.410 0.370 3.480 0.930 ;
        RECT  3.325 0.370 3.410 0.440 ;
        RECT  3.230 0.860 3.410 0.930 ;
        RECT  3.255 0.185 3.325 0.440 ;
        RECT  3.035 0.370 3.255 0.440 ;
        RECT  3.185 0.520 3.255 0.780 ;
        RECT  3.010 0.710 3.185 0.780 ;
        RECT  2.965 0.370 3.035 0.640 ;
        RECT  2.940 0.710 3.010 1.050 ;
        RECT  2.720 0.980 2.940 1.050 ;
        RECT  2.790 0.195 2.860 0.900 ;
        RECT  2.680 0.195 2.790 0.265 ;
        RECT  2.650 0.350 2.720 1.050 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.545 0.340 2.570 0.790 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.500 0.340 2.545 1.020 ;
        RECT  2.480 0.340 2.500 0.460 ;
        RECT  2.475 0.720 2.500 1.020 ;
        RECT  2.255 0.720 2.475 0.790 ;
        RECT  2.405 0.510 2.430 0.630 ;
        RECT  2.335 0.375 2.405 0.630 ;
        RECT  2.060 0.375 2.335 0.445 ;
        RECT  2.185 0.520 2.255 0.790 ;
        RECT  1.990 0.375 2.060 0.795 ;
        RECT  1.910 0.375 1.990 0.445 ;
        RECT  1.965 0.725 1.990 0.795 ;
        RECT  1.895 0.725 1.965 0.970 ;
        RECT  1.790 0.585 1.910 0.655 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.570 0.865 1.810 0.935 ;
        RECT  1.720 0.350 1.790 0.795 ;
        RECT  1.520 0.350 1.720 0.420 ;
        RECT  1.500 0.725 1.720 0.795 ;
        RECT  1.500 0.865 1.570 1.055 ;
        RECT  1.410 0.545 1.540 0.615 ;
        RECT  0.685 0.985 1.500 1.055 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.140 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.755 0.350 0.830 0.915 ;
        RECT  0.615 0.810 0.685 1.055 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXQD2BWP

MACRO DFXQD4BWP
    CLASS CORE ;
    FOREIGN DFXQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.105 0.465 ;
        RECT  4.095 0.765 4.105 1.065 ;
        RECT  4.035 0.185 4.095 1.065 ;
        RECT  3.885 0.355 4.035 0.905 ;
        RECT  3.745 0.355 3.885 0.465 ;
        RECT  3.745 0.765 3.885 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.920 0.520 1.015 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.465 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.590 -0.115 3.830 0.115 ;
        RECT  3.470 -0.115 3.590 0.275 ;
        RECT  3.230 -0.115 3.470 0.115 ;
        RECT  3.110 -0.115 3.230 0.275 ;
        RECT  0.330 -0.115 3.110 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.675 4.290 1.375 ;
        RECT  3.940 1.145 4.210 1.375 ;
        RECT  3.840 0.985 3.940 1.375 ;
        RECT  3.565 1.145 3.840 1.375 ;
        RECT  3.495 0.905 3.565 1.375 ;
        RECT  3.205 1.145 3.495 1.375 ;
        RECT  3.135 0.960 3.205 1.375 ;
        RECT  2.390 1.145 3.135 1.375 ;
        RECT  2.270 0.865 2.390 1.375 ;
        RECT  0.330 1.145 2.270 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.355 3.815 0.465 ;
        RECT  3.745 0.765 3.815 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        RECT  3.570 0.545 3.680 0.615 ;
        RECT  3.500 0.370 3.570 0.805 ;
        RECT  3.385 0.370 3.500 0.440 ;
        RECT  3.385 0.735 3.500 0.805 ;
        RECT  3.315 0.185 3.385 0.440 ;
        RECT  3.315 0.735 3.385 1.035 ;
        RECT  3.230 0.545 3.350 0.615 ;
        RECT  3.075 0.370 3.315 0.440 ;
        RECT  3.160 0.545 3.230 0.860 ;
        RECT  3.040 0.790 3.160 0.860 ;
        RECT  3.005 0.370 3.075 0.640 ;
        RECT  2.970 0.790 3.040 1.060 ;
        RECT  2.730 0.990 2.970 1.060 ;
        RECT  2.810 0.195 2.880 0.910 ;
        RECT  2.700 0.195 2.810 0.265 ;
        RECT  2.800 0.790 2.810 0.910 ;
        RECT  2.730 0.350 2.740 0.470 ;
        RECT  2.660 0.350 2.730 1.060 ;
        RECT  2.580 0.185 2.700 0.265 ;
        RECT  2.555 0.350 2.590 0.790 ;
        RECT  2.030 0.195 2.580 0.265 ;
        RECT  2.520 0.350 2.555 1.040 ;
        RECT  2.500 0.350 2.520 0.470 ;
        RECT  2.485 0.720 2.520 1.040 ;
        RECT  2.275 0.720 2.485 0.790 ;
        RECT  2.425 0.520 2.450 0.640 ;
        RECT  2.355 0.375 2.425 0.640 ;
        RECT  2.125 0.375 2.355 0.445 ;
        RECT  2.205 0.520 2.275 0.790 ;
        RECT  2.055 0.375 2.125 0.795 ;
        RECT  1.930 0.375 2.055 0.445 ;
        RECT  2.005 0.725 2.055 0.795 ;
        RECT  1.935 0.725 2.005 0.970 ;
        RECT  1.810 0.575 1.970 0.645 ;
        RECT  0.610 0.210 1.860 0.280 ;
        RECT  1.590 0.865 1.850 0.935 ;
        RECT  1.740 0.350 1.810 0.795 ;
        RECT  1.540 0.350 1.740 0.420 ;
        RECT  1.540 0.725 1.740 0.795 ;
        RECT  1.520 0.865 1.590 1.045 ;
        RECT  1.410 0.545 1.560 0.615 ;
        RECT  0.685 0.975 1.520 1.045 ;
        RECT  1.340 0.350 1.410 0.905 ;
        RECT  1.170 0.350 1.340 0.420 ;
        RECT  1.140 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.930 0.420 ;
        RECT  0.830 0.835 0.900 0.905 ;
        RECT  0.755 0.350 0.830 0.905 ;
        RECT  0.615 0.810 0.685 1.045 ;
        RECT  0.525 0.565 0.620 0.635 ;
        RECT  0.455 0.350 0.525 0.915 ;
        RECT  0.125 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END DFXQD4BWP

MACRO EDFCND1BWP
    CLASS CORE ;
    FOREIGN EDFCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.585 1.050 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.730 4.515 1.050 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.350 4.285 0.905 ;
        RECT  4.185 0.350 4.215 0.485 ;
        RECT  4.095 0.775 4.215 0.905 ;
        RECT  4.095 0.185 4.185 0.485 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.350 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0352 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.495 3.745 0.770 ;
        RECT  3.625 0.600 3.655 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.280 ;
        RECT  3.650 -0.115 4.280 0.115 ;
        RECT  3.530 -0.115 3.650 0.255 ;
        RECT  2.570 -0.115 3.530 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.475 -0.115 2.500 0.115 ;
        RECT  1.355 -0.115 1.475 0.125 ;
        RECT  1.140 -0.115 1.355 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 1.120 4.400 1.375 ;
        RECT  4.040 1.145 4.280 1.375 ;
        RECT  3.920 1.120 4.040 1.375 ;
        RECT  3.620 1.145 3.920 1.375 ;
        RECT  3.500 1.130 3.620 1.375 ;
        RECT  2.610 1.145 3.500 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  1.120 1.145 1.360 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.640 ;
        RECT  4.355 0.520 4.425 1.050 ;
        RECT  3.360 0.980 4.355 1.050 ;
        RECT  4.025 0.555 4.100 0.625 ;
        RECT  3.955 0.185 4.025 0.910 ;
        RECT  3.920 0.185 3.955 0.285 ;
        RECT  3.500 0.840 3.955 0.910 ;
        RECT  3.815 0.355 3.885 0.720 ;
        RECT  3.660 0.355 3.815 0.425 ;
        RECT  3.590 0.345 3.660 0.425 ;
        RECT  3.045 0.345 3.590 0.415 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.485 3.450 0.555 ;
        RECT  2.720 0.205 3.360 0.275 ;
        RECT  3.290 0.485 3.360 1.050 ;
        RECT  3.150 0.485 3.290 0.555 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  2.975 0.345 3.045 0.705 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.205 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.620 0.195 1.860 0.265 ;
        RECT  1.730 0.995 1.860 1.075 ;
        RECT  1.715 0.345 1.785 0.770 ;
        RECT  0.610 0.995 1.730 1.065 ;
        RECT  1.575 0.345 1.715 0.465 ;
        RECT  1.570 0.700 1.715 0.770 ;
        RECT  1.490 0.545 1.590 0.615 ;
        RECT  1.420 0.335 1.490 0.780 ;
        RECT  1.170 0.335 1.420 0.405 ;
        RECT  1.150 0.710 1.420 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCND1BWP

MACRO EDFCND2BWP
    CLASS CORE ;
    FOREIGN EDFCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.355 5.005 0.905 ;
        RECT  4.935 0.185 4.945 1.035 ;
        RECT  4.875 0.185 4.935 0.465 ;
        RECT  4.875 0.735 4.935 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.195 4.585 0.905 ;
        RECT  4.495 0.195 4.515 0.475 ;
        RECT  4.495 0.775 4.515 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.350 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0608 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.255 0.640 ;
        RECT  4.095 0.355 4.165 0.770 ;
        RECT  3.745 0.700 4.095 0.770 ;
        RECT  3.665 0.495 3.745 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.055 -0.115 5.125 0.300 ;
        RECT  4.755 -0.115 5.055 0.115 ;
        RECT  4.685 -0.115 4.755 0.445 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  3.650 -0.115 4.280 0.115 ;
        RECT  3.530 -0.115 3.650 0.275 ;
        RECT  2.570 -0.115 3.530 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.475 -0.115 2.500 0.115 ;
        RECT  1.355 -0.115 1.475 0.125 ;
        RECT  1.140 -0.115 1.355 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.140 1.145 5.180 1.375 ;
        RECT  5.040 0.970 5.140 1.375 ;
        RECT  4.780 1.145 5.040 1.375 ;
        RECT  4.660 1.120 4.780 1.375 ;
        RECT  4.400 1.145 4.660 1.375 ;
        RECT  4.280 1.120 4.400 1.375 ;
        RECT  4.020 1.145 4.280 1.375 ;
        RECT  3.900 1.120 4.020 1.375 ;
        RECT  3.620 1.145 3.900 1.375 ;
        RECT  3.500 1.130 3.620 1.375 ;
        RECT  2.610 1.145 3.500 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  1.120 1.145 1.360 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.770 0.545 4.860 0.615 ;
        RECT  4.700 0.545 4.770 1.050 ;
        RECT  3.360 0.980 4.700 1.050 ;
        RECT  4.405 0.520 4.440 0.640 ;
        RECT  4.335 0.210 4.405 0.910 ;
        RECT  3.910 0.210 4.335 0.280 ;
        RECT  3.500 0.840 4.335 0.910 ;
        RECT  3.875 0.355 4.005 0.615 ;
        RECT  3.660 0.355 3.875 0.425 ;
        RECT  3.590 0.345 3.660 0.425 ;
        RECT  3.045 0.345 3.590 0.415 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.485 3.450 0.555 ;
        RECT  2.720 0.205 3.360 0.275 ;
        RECT  3.290 0.485 3.360 1.050 ;
        RECT  3.150 0.485 3.290 0.555 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  2.975 0.345 3.045 0.705 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.205 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.620 0.195 1.860 0.265 ;
        RECT  1.730 0.995 1.860 1.075 ;
        RECT  1.715 0.345 1.785 0.770 ;
        RECT  0.610 0.995 1.730 1.065 ;
        RECT  1.575 0.345 1.715 0.465 ;
        RECT  1.570 0.700 1.715 0.770 ;
        RECT  1.490 0.545 1.590 0.615 ;
        RECT  1.420 0.335 1.490 0.780 ;
        RECT  1.170 0.335 1.420 0.405 ;
        RECT  1.150 0.710 1.420 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCND2BWP

MACRO EDFCND4BWP
    CLASS CORE ;
    FOREIGN EDFCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.185 6.065 0.465 ;
        RECT  6.055 0.735 6.065 1.075 ;
        RECT  5.995 0.185 6.055 1.075 ;
        RECT  5.845 0.355 5.995 0.905 ;
        RECT  5.705 0.355 5.845 0.465 ;
        RECT  5.705 0.735 5.845 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.735 5.705 1.075 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.710 5.340 0.810 ;
        RECT  5.255 0.185 5.325 0.465 ;
        RECT  5.215 0.355 5.255 0.465 ;
        RECT  5.005 0.355 5.215 0.810 ;
        RECT  4.965 0.355 5.005 0.465 ;
        RECT  4.880 0.710 5.005 0.810 ;
        RECT  4.895 0.185 4.965 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.530 1.225 0.630 ;
        RECT  1.015 0.355 1.085 0.630 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.255 0.640 ;
        RECT  4.095 0.355 4.165 0.770 ;
        RECT  3.745 0.700 4.095 0.770 ;
        RECT  3.665 0.495 3.745 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 -0.115 6.300 0.115 ;
        RECT  6.175 -0.115 6.245 0.465 ;
        RECT  5.910 -0.115 6.175 0.115 ;
        RECT  5.790 -0.115 5.910 0.275 ;
        RECT  5.515 -0.115 5.790 0.115 ;
        RECT  5.445 -0.115 5.515 0.465 ;
        RECT  5.170 -0.115 5.445 0.115 ;
        RECT  5.050 -0.115 5.170 0.275 ;
        RECT  4.780 -0.115 5.050 0.115 ;
        RECT  4.660 -0.115 4.780 0.125 ;
        RECT  4.400 -0.115 4.660 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  3.640 -0.115 4.280 0.115 ;
        RECT  3.520 -0.115 3.640 0.220 ;
        RECT  2.570 -0.115 3.520 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.480 -0.115 2.500 0.115 ;
        RECT  1.360 -0.115 1.480 0.140 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.140 ;
        RECT  0.305 -0.115 1.000 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 1.145 6.300 1.375 ;
        RECT  6.175 0.680 6.245 1.375 ;
        RECT  5.885 1.145 6.175 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  5.540 1.145 5.815 1.375 ;
        RECT  5.420 1.020 5.540 1.375 ;
        RECT  5.170 1.145 5.420 1.375 ;
        RECT  5.050 1.020 5.170 1.375 ;
        RECT  4.810 1.145 5.050 1.375 ;
        RECT  4.690 1.020 4.810 1.375 ;
        RECT  4.400 1.145 4.690 1.375 ;
        RECT  4.280 1.120 4.400 1.375 ;
        RECT  4.020 1.145 4.280 1.375 ;
        RECT  3.900 1.120 4.020 1.375 ;
        RECT  3.620 1.145 3.900 1.375 ;
        RECT  3.500 1.130 3.620 1.375 ;
        RECT  2.610 1.145 3.500 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.130 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.355 5.775 0.465 ;
        RECT  5.705 0.735 5.775 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.735 5.705 1.075 ;
        RECT  5.285 0.710 5.340 0.810 ;
        RECT  5.285 0.185 5.325 0.465 ;
        RECT  4.895 0.185 4.935 0.465 ;
        RECT  4.880 0.710 4.935 0.810 ;
        RECT  5.520 0.545 5.670 0.615 ;
        RECT  5.450 0.545 5.520 0.950 ;
        RECT  4.545 0.880 5.450 0.950 ;
        RECT  4.695 0.210 4.765 0.650 ;
        RECT  4.395 0.210 4.695 0.280 ;
        RECT  4.475 0.360 4.545 1.050 ;
        RECT  3.360 0.980 4.475 1.050 ;
        RECT  4.325 0.210 4.395 0.910 ;
        RECT  3.910 0.210 4.325 0.280 ;
        RECT  3.500 0.840 4.325 0.910 ;
        RECT  3.875 0.350 4.005 0.615 ;
        RECT  3.660 0.350 3.875 0.420 ;
        RECT  3.590 0.290 3.660 0.420 ;
        RECT  3.160 0.290 3.590 0.360 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.430 3.450 0.500 ;
        RECT  3.290 0.430 3.360 1.050 ;
        RECT  3.150 0.480 3.290 0.550 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.090 0.290 3.160 0.410 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  3.045 0.340 3.090 0.410 ;
        RECT  2.975 0.340 3.045 0.705 ;
        RECT  2.720 0.200 2.990 0.270 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.200 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.920 0.210 1.860 0.280 ;
        RECT  1.720 0.990 1.850 1.075 ;
        RECT  1.715 0.350 1.785 0.780 ;
        RECT  0.920 0.990 1.720 1.060 ;
        RECT  1.550 0.350 1.715 0.420 ;
        RECT  1.550 0.710 1.715 0.780 ;
        RECT  1.460 0.545 1.570 0.615 ;
        RECT  1.390 0.350 1.460 0.780 ;
        RECT  1.170 0.350 1.390 0.420 ;
        RECT  1.170 0.710 1.390 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.850 0.195 0.920 0.280 ;
        RECT  0.850 0.990 0.920 1.065 ;
        RECT  0.620 0.195 0.850 0.265 ;
        RECT  0.610 0.995 0.850 1.065 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCND4BWP

MACRO EDFCNQD1BWP
    CLASS CORE ;
    FOREIGN EDFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.355 0.185 4.445 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.350 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0360 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.495 3.745 0.770 ;
        RECT  3.625 0.600 3.655 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.235 -0.115 4.480 0.115 ;
        RECT  4.165 -0.115 4.235 0.465 ;
        RECT  3.650 -0.115 4.165 0.115 ;
        RECT  3.530 -0.115 3.650 0.270 ;
        RECT  2.570 -0.115 3.530 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.475 -0.115 2.500 0.115 ;
        RECT  1.355 -0.115 1.475 0.125 ;
        RECT  1.140 -0.115 1.355 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 1.145 4.480 1.375 ;
        RECT  4.175 0.700 4.245 1.375 ;
        RECT  3.985 1.145 4.175 1.375 ;
        RECT  3.915 0.980 3.985 1.375 ;
        RECT  3.595 1.145 3.915 1.375 ;
        RECT  3.525 0.980 3.595 1.375 ;
        RECT  2.610 1.145 3.525 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  1.120 1.145 1.360 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.035 0.545 4.260 0.615 ;
        RECT  3.965 0.205 4.035 0.910 ;
        RECT  3.890 0.205 3.965 0.275 ;
        RECT  3.805 0.840 3.965 0.910 ;
        RECT  3.825 0.355 3.895 0.720 ;
        RECT  3.660 0.355 3.825 0.425 ;
        RECT  3.735 0.840 3.805 1.075 ;
        RECT  3.500 0.840 3.735 0.910 ;
        RECT  3.590 0.345 3.660 0.425 ;
        RECT  3.045 0.345 3.590 0.415 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.485 3.450 0.555 ;
        RECT  2.720 0.205 3.360 0.275 ;
        RECT  3.290 0.485 3.360 1.050 ;
        RECT  3.150 0.485 3.290 0.555 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  2.975 0.345 3.045 0.705 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.205 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.620 0.195 1.860 0.265 ;
        RECT  1.730 0.995 1.860 1.075 ;
        RECT  1.715 0.345 1.785 0.770 ;
        RECT  0.610 0.995 1.730 1.065 ;
        RECT  1.575 0.345 1.715 0.465 ;
        RECT  1.570 0.700 1.715 0.770 ;
        RECT  1.490 0.545 1.590 0.615 ;
        RECT  1.420 0.335 1.490 0.780 ;
        RECT  1.170 0.335 1.420 0.405 ;
        RECT  1.150 0.710 1.420 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCNQD1BWP

MACRO EDFCNQD2BWP
    CLASS CORE ;
    FOREIGN EDFCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 0.355 4.585 0.905 ;
        RECT  4.515 0.185 4.525 1.035 ;
        RECT  4.455 0.185 4.515 0.465 ;
        RECT  4.455 0.735 4.515 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.350 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0624 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.235 0.640 ;
        RECT  4.095 0.495 4.165 0.770 ;
        RECT  3.745 0.700 4.095 0.770 ;
        RECT  3.665 0.495 3.745 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 -0.115 4.760 0.115 ;
        RECT  4.635 -0.115 4.705 0.300 ;
        RECT  4.370 -0.115 4.635 0.115 ;
        RECT  4.250 -0.115 4.370 0.275 ;
        RECT  3.650 -0.115 4.250 0.115 ;
        RECT  3.530 -0.115 3.650 0.270 ;
        RECT  2.570 -0.115 3.530 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.475 -0.115 2.500 0.115 ;
        RECT  1.355 -0.115 1.475 0.125 ;
        RECT  1.140 -0.115 1.355 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 1.145 4.760 1.375 ;
        RECT  4.635 0.960 4.705 1.375 ;
        RECT  4.345 1.145 4.635 1.375 ;
        RECT  4.275 0.980 4.345 1.375 ;
        RECT  3.985 1.145 4.275 1.375 ;
        RECT  3.915 0.980 3.985 1.375 ;
        RECT  3.595 1.145 3.915 1.375 ;
        RECT  3.525 0.980 3.595 1.375 ;
        RECT  2.610 1.145 3.525 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  1.120 1.145 1.360 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.385 0.520 4.410 0.640 ;
        RECT  4.315 0.345 4.385 0.910 ;
        RECT  4.165 0.345 4.315 0.415 ;
        RECT  4.165 0.840 4.315 0.910 ;
        RECT  4.095 0.195 4.165 0.415 ;
        RECT  4.095 0.840 4.165 1.075 ;
        RECT  3.890 0.195 4.095 0.265 ;
        RECT  3.805 0.840 4.095 0.910 ;
        RECT  3.880 0.345 4.000 0.615 ;
        RECT  3.045 0.345 3.880 0.415 ;
        RECT  3.735 0.840 3.805 1.075 ;
        RECT  3.500 0.840 3.735 0.910 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.485 3.450 0.555 ;
        RECT  2.720 0.205 3.360 0.275 ;
        RECT  3.290 0.485 3.360 1.050 ;
        RECT  3.150 0.485 3.290 0.555 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  2.975 0.345 3.045 0.705 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.205 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.620 0.195 1.860 0.265 ;
        RECT  1.730 0.995 1.860 1.075 ;
        RECT  1.715 0.345 1.785 0.770 ;
        RECT  0.610 0.995 1.730 1.065 ;
        RECT  1.575 0.345 1.715 0.465 ;
        RECT  1.570 0.700 1.715 0.770 ;
        RECT  1.490 0.545 1.590 0.615 ;
        RECT  1.420 0.335 1.490 0.780 ;
        RECT  1.170 0.335 1.420 0.405 ;
        RECT  1.150 0.710 1.420 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCNQD2BWP

MACRO EDFCNQD4BWP
    CLASS CORE ;
    FOREIGN EDFCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 4.945 0.465 ;
        RECT  4.935 0.735 4.945 1.075 ;
        RECT  4.875 0.185 4.935 1.075 ;
        RECT  4.725 0.355 4.875 0.905 ;
        RECT  4.565 0.355 4.725 0.465 ;
        RECT  4.565 0.735 4.725 0.905 ;
        RECT  4.495 0.185 4.565 0.465 ;
        RECT  4.495 0.735 4.565 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.530 1.225 0.630 ;
        RECT  1.015 0.355 1.085 0.630 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 0.495 4.255 0.640 ;
        RECT  4.165 0.355 4.185 0.640 ;
        RECT  4.095 0.355 4.165 0.770 ;
        RECT  3.745 0.700 4.095 0.770 ;
        RECT  3.665 0.495 3.745 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.055 -0.115 5.125 0.465 ;
        RECT  4.780 -0.115 5.055 0.115 ;
        RECT  4.660 -0.115 4.780 0.275 ;
        RECT  4.400 -0.115 4.660 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  3.640 -0.115 4.280 0.115 ;
        RECT  3.520 -0.115 3.640 0.220 ;
        RECT  2.570 -0.115 3.520 0.115 ;
        RECT  2.500 -0.115 2.570 0.265 ;
        RECT  1.480 -0.115 2.500 0.115 ;
        RECT  1.360 -0.115 1.480 0.140 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.140 ;
        RECT  0.305 -0.115 1.000 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.055 0.680 5.125 1.375 ;
        RECT  4.755 1.145 5.055 1.375 ;
        RECT  4.685 0.975 4.755 1.375 ;
        RECT  4.375 1.145 4.685 1.375 ;
        RECT  4.305 0.980 4.375 1.375 ;
        RECT  3.995 1.145 4.305 1.375 ;
        RECT  3.925 0.980 3.995 1.375 ;
        RECT  3.595 1.145 3.925 1.375 ;
        RECT  3.525 0.980 3.595 1.375 ;
        RECT  2.610 1.145 3.525 1.375 ;
        RECT  2.490 1.060 2.610 1.375 ;
        RECT  1.480 1.145 2.490 1.375 ;
        RECT  1.360 1.130 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.355 4.655 0.465 ;
        RECT  4.565 0.735 4.655 0.905 ;
        RECT  4.495 0.185 4.565 0.465 ;
        RECT  4.495 0.735 4.565 1.075 ;
        RECT  4.395 0.545 4.590 0.615 ;
        RECT  4.325 0.210 4.395 0.910 ;
        RECT  3.910 0.210 4.325 0.280 ;
        RECT  4.185 0.840 4.325 0.910 ;
        RECT  4.115 0.840 4.185 1.075 ;
        RECT  3.805 0.840 4.115 0.910 ;
        RECT  3.875 0.350 4.005 0.615 ;
        RECT  3.660 0.350 3.875 0.420 ;
        RECT  3.735 0.840 3.805 1.075 ;
        RECT  3.500 0.840 3.735 0.910 ;
        RECT  3.590 0.290 3.660 0.420 ;
        RECT  3.160 0.290 3.590 0.360 ;
        RECT  3.430 0.650 3.500 0.910 ;
        RECT  3.360 0.430 3.450 0.500 ;
        RECT  3.290 0.430 3.360 1.050 ;
        RECT  3.150 0.480 3.290 0.550 ;
        RECT  2.750 0.980 3.290 1.050 ;
        RECT  3.095 0.635 3.165 0.910 ;
        RECT  3.090 0.290 3.160 0.410 ;
        RECT  3.045 0.635 3.095 0.705 ;
        RECT  3.045 0.340 3.090 0.410 ;
        RECT  2.975 0.340 3.045 0.705 ;
        RECT  2.720 0.200 2.990 0.270 ;
        RECT  2.870 0.785 2.990 0.855 ;
        RECT  2.800 0.350 2.870 0.855 ;
        RECT  2.310 0.475 2.800 0.545 ;
        RECT  2.680 0.920 2.750 1.050 ;
        RECT  2.650 0.200 2.720 0.405 ;
        RECT  2.085 0.630 2.720 0.700 ;
        RECT  2.375 0.920 2.680 0.990 ;
        RECT  2.300 0.335 2.650 0.405 ;
        RECT  2.225 0.770 2.610 0.850 ;
        RECT  2.305 0.920 2.375 1.045 ;
        RECT  2.190 0.475 2.310 0.560 ;
        RECT  2.010 0.975 2.305 1.045 ;
        RECT  2.230 0.195 2.300 0.405 ;
        RECT  2.160 0.195 2.230 0.265 ;
        RECT  2.155 0.770 2.225 0.900 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.015 0.345 2.085 0.780 ;
        RECT  1.930 0.345 2.015 0.415 ;
        RECT  1.940 0.710 2.015 0.780 ;
        RECT  1.940 0.850 2.010 1.045 ;
        RECT  1.020 0.850 1.940 0.920 ;
        RECT  1.785 0.555 1.930 0.625 ;
        RECT  0.920 0.210 1.860 0.280 ;
        RECT  1.720 0.990 1.850 1.075 ;
        RECT  1.715 0.350 1.785 0.780 ;
        RECT  0.920 0.990 1.720 1.060 ;
        RECT  1.550 0.350 1.715 0.420 ;
        RECT  1.550 0.710 1.715 0.780 ;
        RECT  1.460 0.545 1.570 0.615 ;
        RECT  1.390 0.350 1.460 0.780 ;
        RECT  1.170 0.350 1.390 0.420 ;
        RECT  1.170 0.710 1.390 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.850 0.195 0.920 0.280 ;
        RECT  0.850 0.990 0.920 1.065 ;
        RECT  0.620 0.195 0.850 0.265 ;
        RECT  0.610 0.995 0.850 1.065 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFCNQD4BWP

MACRO EDFD1BWP
    CLASS CORE ;
    FOREIGN EDFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.350 3.625 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.550 1.225 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 -0.115 4.060 0.115 ;
        RECT  3.720 -0.115 3.840 0.140 ;
        RECT  3.220 -0.115 3.720 0.115 ;
        RECT  3.100 -0.115 3.220 0.140 ;
        RECT  2.375 -0.115 3.100 0.115 ;
        RECT  2.305 -0.115 2.375 0.420 ;
        RECT  1.440 -0.115 2.305 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.145 4.060 1.375 ;
        RECT  3.720 1.130 3.840 1.375 ;
        RECT  3.220 1.145 3.720 1.375 ;
        RECT  3.100 1.130 3.220 1.375 ;
        RECT  2.380 1.145 3.100 1.375 ;
        RECT  2.255 1.020 2.380 1.375 ;
        RECT  1.420 1.145 2.255 1.375 ;
        RECT  1.300 1.135 1.420 1.375 ;
        RECT  1.120 1.145 1.300 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 0.520 3.875 0.640 ;
        RECT  3.740 0.210 3.810 1.060 ;
        RECT  3.000 0.210 3.740 0.280 ;
        RECT  2.540 0.990 3.740 1.060 ;
        RECT  3.395 0.375 3.465 0.870 ;
        RECT  3.150 0.375 3.395 0.445 ;
        RECT  3.280 0.800 3.395 0.870 ;
        RECT  3.190 0.545 3.310 0.640 ;
        RECT  3.100 0.570 3.190 0.640 ;
        RECT  3.080 0.375 3.150 0.485 ;
        RECT  3.030 0.570 3.100 0.920 ;
        RECT  2.970 0.415 3.080 0.485 ;
        RECT  2.860 0.570 3.030 0.640 ;
        RECT  2.650 0.850 3.030 0.920 ;
        RECT  2.930 0.210 3.000 0.330 ;
        RECT  2.710 0.710 2.930 0.780 ;
        RECT  2.790 0.220 2.860 0.640 ;
        RECT  2.710 0.220 2.790 0.290 ;
        RECT  2.640 0.370 2.710 0.780 ;
        RECT  2.500 0.210 2.570 0.790 ;
        RECT  2.470 0.870 2.540 1.060 ;
        RECT  2.280 0.720 2.500 0.790 ;
        RECT  2.085 0.870 2.470 0.940 ;
        RECT  2.360 0.510 2.430 0.640 ;
        RECT  2.010 0.510 2.360 0.580 ;
        RECT  2.160 0.670 2.280 0.790 ;
        RECT  2.015 0.855 2.085 0.940 ;
        RECT  1.020 0.855 2.015 0.925 ;
        RECT  1.935 0.300 2.010 0.775 ;
        RECT  1.870 0.705 1.935 0.775 ;
        RECT  0.620 0.195 1.840 0.265 ;
        RECT  1.680 0.995 1.800 1.075 ;
        RECT  1.705 0.335 1.775 0.785 ;
        RECT  1.530 0.335 1.705 0.405 ;
        RECT  1.510 0.715 1.705 0.785 ;
        RECT  0.610 0.995 1.680 1.065 ;
        RECT  1.375 0.545 1.550 0.615 ;
        RECT  1.305 0.335 1.375 0.785 ;
        RECT  1.170 0.335 1.305 0.405 ;
        RECT  1.150 0.715 1.305 0.785 ;
        RECT  0.900 0.700 1.020 0.925 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFD1BWP

MACRO EDFD2BWP
    CLASS CORE ;
    FOREIGN EDFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.905 ;
        RECT  4.230 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.230 0.465 ;
        RECT  4.175 0.735 4.230 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.350 3.885 0.905 ;
        RECT  3.795 0.350 3.815 0.470 ;
        RECT  3.795 0.765 3.815 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.540 1.225 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 -0.115 4.480 0.115 ;
        RECT  4.355 -0.115 4.425 0.305 ;
        RECT  4.080 -0.115 4.355 0.115 ;
        RECT  3.960 -0.115 4.080 0.140 ;
        RECT  3.690 -0.115 3.960 0.115 ;
        RECT  3.570 -0.115 3.690 0.140 ;
        RECT  3.300 -0.115 3.570 0.115 ;
        RECT  3.180 -0.115 3.300 0.140 ;
        RECT  2.375 -0.115 3.180 0.115 ;
        RECT  2.305 -0.115 2.375 0.420 ;
        RECT  1.440 -0.115 2.305 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 1.145 4.480 1.375 ;
        RECT  4.355 0.960 4.425 1.375 ;
        RECT  4.080 1.145 4.355 1.375 ;
        RECT  3.960 1.120 4.080 1.375 ;
        RECT  3.690 1.145 3.960 1.375 ;
        RECT  3.570 1.120 3.690 1.375 ;
        RECT  3.300 1.145 3.570 1.375 ;
        RECT  3.180 1.135 3.300 1.375 ;
        RECT  2.400 1.145 3.180 1.375 ;
        RECT  2.275 1.020 2.400 1.375 ;
        RECT  1.420 1.145 2.275 1.375 ;
        RECT  1.300 1.135 1.420 1.375 ;
        RECT  1.120 1.145 1.300 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.085 0.520 4.130 0.640 ;
        RECT  4.015 0.210 4.085 1.050 ;
        RECT  3.070 0.210 4.015 0.280 ;
        RECT  3.265 0.980 4.015 1.050 ;
        RECT  3.640 0.520 3.745 0.640 ;
        RECT  3.570 0.365 3.640 0.910 ;
        RECT  3.240 0.365 3.570 0.435 ;
        RECT  3.380 0.840 3.570 0.910 ;
        RECT  3.345 0.520 3.415 0.770 ;
        RECT  3.070 0.700 3.345 0.770 ;
        RECT  3.195 0.980 3.265 1.065 ;
        RECT  3.140 0.365 3.240 0.630 ;
        RECT  2.540 0.995 3.195 1.065 ;
        RECT  2.970 0.210 3.070 0.310 ;
        RECT  3.000 0.540 3.070 0.925 ;
        RECT  2.860 0.540 3.000 0.610 ;
        RECT  2.670 0.855 3.000 0.925 ;
        RECT  2.710 0.715 2.920 0.785 ;
        RECT  2.790 0.220 2.860 0.610 ;
        RECT  2.710 0.220 2.790 0.290 ;
        RECT  2.640 0.370 2.710 0.785 ;
        RECT  2.500 0.210 2.570 0.790 ;
        RECT  2.470 0.870 2.540 1.065 ;
        RECT  2.280 0.720 2.500 0.790 ;
        RECT  2.085 0.870 2.470 0.940 ;
        RECT  2.360 0.510 2.430 0.640 ;
        RECT  2.010 0.510 2.360 0.580 ;
        RECT  2.160 0.670 2.280 0.790 ;
        RECT  2.015 0.855 2.085 0.940 ;
        RECT  1.020 0.855 2.015 0.925 ;
        RECT  1.935 0.300 2.010 0.775 ;
        RECT  1.870 0.705 1.935 0.775 ;
        RECT  0.620 0.195 1.840 0.265 ;
        RECT  1.680 0.995 1.800 1.075 ;
        RECT  1.705 0.335 1.775 0.785 ;
        RECT  1.530 0.335 1.705 0.405 ;
        RECT  1.510 0.715 1.705 0.785 ;
        RECT  0.610 0.995 1.680 1.065 ;
        RECT  1.375 0.545 1.550 0.615 ;
        RECT  1.305 0.335 1.375 0.785 ;
        RECT  1.170 0.335 1.305 0.405 ;
        RECT  1.150 0.715 1.305 0.785 ;
        RECT  0.900 0.700 1.020 0.925 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFD2BWP

MACRO EDFD4BWP
    CLASS CORE ;
    FOREIGN EDFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.765 4.945 1.065 ;
        RECT  4.795 0.355 4.875 0.465 ;
        RECT  4.795 0.765 4.875 0.905 ;
        RECT  4.585 0.355 4.795 0.905 ;
        RECT  4.565 0.355 4.585 0.465 ;
        RECT  4.495 0.765 4.585 1.075 ;
        RECT  4.495 0.185 4.565 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.710 4.230 0.800 ;
        RECT  4.095 0.355 4.210 0.450 ;
        RECT  3.885 0.355 4.095 0.800 ;
        RECT  3.710 0.355 3.885 0.450 ;
        RECT  3.750 0.710 3.885 0.800 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.210 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.055 -0.115 5.125 0.465 ;
        RECT  4.755 -0.115 5.055 0.115 ;
        RECT  4.685 -0.115 4.755 0.285 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.145 ;
        RECT  4.020 -0.115 4.280 0.115 ;
        RECT  3.900 -0.115 4.020 0.145 ;
        RECT  3.640 -0.115 3.900 0.115 ;
        RECT  3.520 -0.115 3.640 0.145 ;
        RECT  3.260 -0.115 3.520 0.115 ;
        RECT  3.140 -0.115 3.260 0.145 ;
        RECT  2.380 -0.115 3.140 0.115 ;
        RECT  2.260 -0.115 2.380 0.125 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.140 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.140 ;
        RECT  0.305 -0.115 1.000 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.055 0.680 5.125 1.375 ;
        RECT  4.755 1.145 5.055 1.375 ;
        RECT  4.685 0.975 4.755 1.375 ;
        RECT  4.410 1.145 4.685 1.375 ;
        RECT  4.290 1.010 4.410 1.375 ;
        RECT  4.050 1.145 4.290 1.375 ;
        RECT  3.930 1.010 4.050 1.375 ;
        RECT  3.680 1.145 3.930 1.375 ;
        RECT  3.560 1.010 3.680 1.375 ;
        RECT  3.300 1.145 3.560 1.375 ;
        RECT  3.180 1.130 3.300 1.375 ;
        RECT  2.395 1.145 3.180 1.375 ;
        RECT  2.325 1.010 2.395 1.375 ;
        RECT  1.460 1.145 2.325 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.100 1.145 1.340 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.765 4.945 1.065 ;
        RECT  4.865 0.355 4.875 0.465 ;
        RECT  4.865 0.765 4.875 0.905 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.765 4.515 1.075 ;
        RECT  4.165 0.710 4.230 0.800 ;
        RECT  4.165 0.355 4.210 0.450 ;
        RECT  3.710 0.355 3.815 0.450 ;
        RECT  3.750 0.710 3.815 0.800 ;
        RECT  4.370 0.545 4.490 0.615 ;
        RECT  4.300 0.215 4.370 0.940 ;
        RECT  3.030 0.215 4.300 0.285 ;
        RECT  3.475 0.870 4.300 0.940 ;
        RECT  3.600 0.545 3.780 0.615 ;
        RECT  3.530 0.370 3.600 0.800 ;
        RECT  3.170 0.370 3.530 0.440 ;
        RECT  3.380 0.700 3.530 0.800 ;
        RECT  3.405 0.870 3.475 1.060 ;
        RECT  3.310 0.545 3.450 0.615 ;
        RECT  2.590 0.990 3.405 1.060 ;
        RECT  3.240 0.545 3.310 0.920 ;
        RECT  2.750 0.850 3.240 0.920 ;
        RECT  3.100 0.370 3.170 0.630 ;
        RECT  3.070 0.530 3.100 0.630 ;
        RECT  2.960 0.215 3.030 0.385 ;
        RECT  2.890 0.675 2.990 0.745 ;
        RECT  2.820 0.195 2.890 0.745 ;
        RECT  2.720 0.195 2.820 0.265 ;
        RECT  2.680 0.345 2.750 0.920 ;
        RECT  2.570 0.185 2.720 0.265 ;
        RECT  2.540 0.345 2.610 0.780 ;
        RECT  2.520 0.850 2.590 1.060 ;
        RECT  2.040 0.195 2.570 0.265 ;
        RECT  2.270 0.345 2.540 0.415 ;
        RECT  2.490 0.710 2.540 0.780 ;
        RECT  1.020 0.850 2.520 0.920 ;
        RECT  2.410 0.520 2.460 0.640 ;
        RECT  2.340 0.520 2.410 0.780 ;
        RECT  2.015 0.710 2.340 0.780 ;
        RECT  2.200 0.345 2.270 0.630 ;
        RECT  1.945 0.350 2.015 0.780 ;
        RECT  1.910 0.710 1.945 0.780 ;
        RECT  0.920 0.210 1.850 0.280 ;
        RECT  0.920 0.990 1.830 1.060 ;
        RECT  1.740 0.350 1.810 0.780 ;
        RECT  1.550 0.350 1.740 0.420 ;
        RECT  1.530 0.710 1.740 0.780 ;
        RECT  1.450 0.545 1.570 0.615 ;
        RECT  1.380 0.350 1.450 0.780 ;
        RECT  1.170 0.350 1.380 0.420 ;
        RECT  1.150 0.710 1.380 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.850 0.195 0.920 0.280 ;
        RECT  0.850 0.990 0.920 1.065 ;
        RECT  0.620 0.195 0.850 0.265 ;
        RECT  0.610 0.995 0.850 1.065 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFD4BWP

MACRO EDFKCND1BWP
    CLASS CORE ;
    FOREIGN EDFKCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.185 4.445 1.045 ;
        RECT  4.355 0.185 4.375 0.465 ;
        RECT  4.355 0.735 4.375 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.350 4.045 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.645 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 -0.115 4.480 0.115 ;
        RECT  4.140 -0.115 4.260 0.140 ;
        RECT  3.620 -0.115 4.140 0.115 ;
        RECT  3.500 -0.115 3.620 0.140 ;
        RECT  2.775 -0.115 3.500 0.115 ;
        RECT  2.705 -0.115 2.775 0.420 ;
        RECT  1.800 -0.115 2.705 0.115 ;
        RECT  1.680 -0.115 1.800 0.125 ;
        RECT  1.440 -0.115 1.680 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  0.330 -0.115 1.320 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.145 4.480 1.375 ;
        RECT  4.140 1.130 4.260 1.375 ;
        RECT  3.620 1.145 4.140 1.375 ;
        RECT  3.500 1.130 3.620 1.375 ;
        RECT  2.780 1.145 3.500 1.375 ;
        RECT  2.655 1.020 2.780 1.375 ;
        RECT  1.800 1.145 2.655 1.375 ;
        RECT  1.680 1.135 1.800 1.375 ;
        RECT  1.220 1.145 1.680 1.375 ;
        RECT  1.100 1.120 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.230 0.520 4.295 0.640 ;
        RECT  4.160 0.210 4.230 1.060 ;
        RECT  3.400 0.210 4.160 0.280 ;
        RECT  2.940 0.990 4.160 1.060 ;
        RECT  3.815 0.375 3.885 0.870 ;
        RECT  3.540 0.375 3.815 0.445 ;
        RECT  3.680 0.800 3.815 0.870 ;
        RECT  3.580 0.545 3.700 0.640 ;
        RECT  3.500 0.570 3.580 0.640 ;
        RECT  3.470 0.375 3.540 0.485 ;
        RECT  3.430 0.570 3.500 0.920 ;
        RECT  3.370 0.415 3.470 0.485 ;
        RECT  3.260 0.570 3.430 0.640 ;
        RECT  3.050 0.850 3.430 0.920 ;
        RECT  3.330 0.210 3.400 0.330 ;
        RECT  3.110 0.710 3.330 0.780 ;
        RECT  3.190 0.220 3.260 0.640 ;
        RECT  3.110 0.220 3.190 0.290 ;
        RECT  3.040 0.370 3.110 0.780 ;
        RECT  2.900 0.210 2.970 0.790 ;
        RECT  2.870 0.870 2.940 1.060 ;
        RECT  2.680 0.720 2.900 0.790 ;
        RECT  2.465 0.870 2.870 0.940 ;
        RECT  2.760 0.510 2.830 0.640 ;
        RECT  2.390 0.510 2.760 0.580 ;
        RECT  2.560 0.670 2.680 0.790 ;
        RECT  2.395 0.855 2.465 0.940 ;
        RECT  1.710 0.855 2.395 0.925 ;
        RECT  2.315 0.300 2.390 0.775 ;
        RECT  2.250 0.705 2.315 0.775 ;
        RECT  0.750 0.200 2.220 0.270 ;
        RECT  2.060 0.995 2.180 1.075 ;
        RECT  2.085 0.355 2.155 0.775 ;
        RECT  1.890 0.355 2.085 0.425 ;
        RECT  1.890 0.705 2.085 0.775 ;
        RECT  1.540 0.995 2.060 1.065 ;
        RECT  1.785 0.545 1.910 0.615 ;
        RECT  1.715 0.355 1.785 0.770 ;
        RECT  1.470 0.355 1.715 0.425 ;
        RECT  1.470 0.700 1.715 0.770 ;
        RECT  1.640 0.840 1.710 0.925 ;
        RECT  1.115 0.840 1.640 0.910 ;
        RECT  1.470 0.980 1.540 1.065 ;
        RECT  0.810 0.980 1.470 1.050 ;
        RECT  0.485 0.340 1.230 0.410 ;
        RECT  1.045 0.520 1.115 0.910 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.790 0.810 1.050 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCND1BWP

MACRO EDFKCND2BWP
    CLASS CORE ;
    FOREIGN EDFKCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 0.355 4.585 0.905 ;
        RECT  4.515 0.185 4.525 1.035 ;
        RECT  4.455 0.185 4.515 0.465 ;
        RECT  4.455 0.735 4.515 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.350 4.165 0.905 ;
        RECT  4.080 0.350 4.095 0.470 ;
        RECT  4.075 0.775 4.095 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.645 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 -0.115 4.760 0.115 ;
        RECT  4.635 -0.115 4.705 0.300 ;
        RECT  4.360 -0.115 4.635 0.115 ;
        RECT  4.240 -0.115 4.360 0.140 ;
        RECT  3.970 -0.115 4.240 0.115 ;
        RECT  3.850 -0.115 3.970 0.140 ;
        RECT  3.600 -0.115 3.850 0.115 ;
        RECT  3.480 -0.115 3.600 0.140 ;
        RECT  2.735 -0.115 3.480 0.115 ;
        RECT  2.665 -0.115 2.735 0.420 ;
        RECT  1.780 -0.115 2.665 0.115 ;
        RECT  1.660 -0.115 1.780 0.125 ;
        RECT  1.440 -0.115 1.660 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  0.330 -0.115 1.320 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 1.145 4.760 1.375 ;
        RECT  4.635 0.960 4.705 1.375 ;
        RECT  4.360 1.145 4.635 1.375 ;
        RECT  4.240 1.130 4.360 1.375 ;
        RECT  3.970 1.145 4.240 1.375 ;
        RECT  3.850 1.130 3.970 1.375 ;
        RECT  3.600 1.145 3.850 1.375 ;
        RECT  3.480 1.130 3.600 1.375 ;
        RECT  2.760 1.145 3.480 1.375 ;
        RECT  2.635 1.020 2.760 1.375 ;
        RECT  1.780 1.145 2.635 1.375 ;
        RECT  1.660 1.135 1.780 1.375 ;
        RECT  1.220 1.145 1.660 1.375 ;
        RECT  1.100 1.120 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.545 4.440 0.615 ;
        RECT  4.280 0.210 4.350 1.060 ;
        RECT  3.375 0.210 4.280 0.280 ;
        RECT  2.900 0.990 4.280 1.060 ;
        RECT  3.970 0.520 4.025 0.640 ;
        RECT  3.900 0.365 3.970 0.920 ;
        RECT  3.540 0.365 3.900 0.435 ;
        RECT  3.670 0.850 3.900 0.920 ;
        RECT  3.625 0.520 3.695 0.780 ;
        RECT  3.380 0.710 3.625 0.780 ;
        RECT  3.450 0.365 3.540 0.640 ;
        RECT  3.310 0.520 3.380 0.920 ;
        RECT  3.285 0.185 3.375 0.445 ;
        RECT  3.210 0.520 3.310 0.590 ;
        RECT  3.030 0.850 3.310 0.920 ;
        RECT  3.070 0.660 3.240 0.780 ;
        RECT  3.140 0.190 3.210 0.590 ;
        RECT  3.030 0.190 3.140 0.260 ;
        RECT  3.000 0.340 3.070 0.780 ;
        RECT  2.860 0.190 2.930 0.790 ;
        RECT  2.830 0.870 2.900 1.060 ;
        RECT  2.640 0.720 2.860 0.790 ;
        RECT  2.445 0.870 2.830 0.940 ;
        RECT  2.720 0.510 2.790 0.640 ;
        RECT  2.370 0.510 2.720 0.580 ;
        RECT  2.520 0.670 2.640 0.790 ;
        RECT  2.375 0.855 2.445 0.940 ;
        RECT  1.710 0.855 2.375 0.925 ;
        RECT  2.295 0.300 2.370 0.775 ;
        RECT  2.230 0.705 2.295 0.775 ;
        RECT  0.750 0.200 2.200 0.270 ;
        RECT  2.040 0.995 2.160 1.075 ;
        RECT  2.065 0.355 2.135 0.775 ;
        RECT  1.870 0.355 2.065 0.425 ;
        RECT  1.870 0.705 2.065 0.775 ;
        RECT  1.540 0.995 2.040 1.065 ;
        RECT  1.785 0.545 1.890 0.615 ;
        RECT  1.715 0.355 1.785 0.770 ;
        RECT  1.490 0.355 1.715 0.425 ;
        RECT  1.490 0.700 1.715 0.770 ;
        RECT  1.640 0.840 1.710 0.925 ;
        RECT  1.115 0.840 1.640 0.910 ;
        RECT  1.470 0.980 1.540 1.065 ;
        RECT  0.810 0.980 1.470 1.050 ;
        RECT  0.485 0.340 1.230 0.410 ;
        RECT  1.045 0.520 1.115 0.910 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.790 0.810 1.050 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCND2BWP

MACRO EDFKCND4BWP
    CLASS CORE ;
    FOREIGN EDFKCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.155 0.185 5.225 0.465 ;
        RECT  5.155 0.775 5.225 1.075 ;
        RECT  5.075 0.355 5.155 0.465 ;
        RECT  5.075 0.775 5.155 0.905 ;
        RECT  4.885 0.355 5.075 0.905 ;
        RECT  4.865 0.355 4.885 1.075 ;
        RECT  4.795 0.185 4.865 0.465 ;
        RECT  4.795 0.775 4.865 1.075 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.710 4.530 0.800 ;
        RECT  4.375 0.355 4.510 0.460 ;
        RECT  4.165 0.355 4.375 0.800 ;
        RECT  4.010 0.355 4.165 0.460 ;
        RECT  4.050 0.710 4.165 0.800 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.650 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.405 -0.115 5.460 0.115 ;
        RECT  5.335 -0.115 5.405 0.465 ;
        RECT  5.045 -0.115 5.335 0.115 ;
        RECT  4.975 -0.115 5.045 0.285 ;
        RECT  4.700 -0.115 4.975 0.115 ;
        RECT  4.580 -0.115 4.700 0.145 ;
        RECT  4.320 -0.115 4.580 0.115 ;
        RECT  4.200 -0.115 4.320 0.145 ;
        RECT  3.940 -0.115 4.200 0.115 ;
        RECT  3.820 -0.115 3.940 0.145 ;
        RECT  3.560 -0.115 3.820 0.115 ;
        RECT  3.440 -0.115 3.560 0.145 ;
        RECT  2.680 -0.115 3.440 0.115 ;
        RECT  2.560 -0.115 2.680 0.125 ;
        RECT  1.780 -0.115 2.560 0.115 ;
        RECT  1.660 -0.115 1.780 0.140 ;
        RECT  1.420 -0.115 1.660 0.115 ;
        RECT  1.300 -0.115 1.420 0.140 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.405 1.145 5.460 1.375 ;
        RECT  5.335 0.680 5.405 1.375 ;
        RECT  5.045 1.145 5.335 1.375 ;
        RECT  4.975 0.975 5.045 1.375 ;
        RECT  4.710 1.145 4.975 1.375 ;
        RECT  4.590 1.010 4.710 1.375 ;
        RECT  4.350 1.145 4.590 1.375 ;
        RECT  4.230 1.010 4.350 1.375 ;
        RECT  3.980 1.145 4.230 1.375 ;
        RECT  3.860 1.130 3.980 1.375 ;
        RECT  3.580 1.145 3.860 1.375 ;
        RECT  3.460 1.130 3.580 1.375 ;
        RECT  2.740 1.145 3.460 1.375 ;
        RECT  2.620 1.015 2.740 1.375 ;
        RECT  1.780 1.145 2.620 1.375 ;
        RECT  1.660 1.130 1.780 1.375 ;
        RECT  1.220 1.145 1.660 1.375 ;
        RECT  1.100 1.130 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.155 0.185 5.225 0.465 ;
        RECT  5.155 0.775 5.225 1.075 ;
        RECT  5.145 0.355 5.155 0.465 ;
        RECT  5.145 0.775 5.155 0.905 ;
        RECT  4.445 0.710 4.530 0.800 ;
        RECT  4.445 0.355 4.510 0.460 ;
        RECT  4.010 0.355 4.095 0.460 ;
        RECT  4.050 0.710 4.095 0.800 ;
        RECT  4.670 0.545 4.780 0.615 ;
        RECT  4.600 0.215 4.670 0.940 ;
        RECT  3.330 0.215 4.600 0.285 ;
        RECT  4.110 0.870 4.600 0.940 ;
        RECT  4.040 0.870 4.110 1.060 ;
        RECT  3.900 0.545 4.080 0.615 ;
        RECT  2.910 0.990 4.040 1.060 ;
        RECT  3.830 0.370 3.900 0.815 ;
        RECT  3.470 0.370 3.830 0.440 ;
        RECT  3.680 0.695 3.830 0.815 ;
        RECT  3.610 0.545 3.750 0.615 ;
        RECT  3.540 0.545 3.610 0.920 ;
        RECT  3.050 0.850 3.540 0.920 ;
        RECT  3.400 0.370 3.470 0.630 ;
        RECT  3.370 0.530 3.400 0.630 ;
        RECT  3.260 0.215 3.330 0.430 ;
        RECT  3.190 0.685 3.290 0.755 ;
        RECT  3.120 0.195 3.190 0.755 ;
        RECT  3.000 0.195 3.120 0.265 ;
        RECT  2.980 0.345 3.050 0.920 ;
        RECT  2.880 0.185 3.000 0.265 ;
        RECT  2.840 0.345 2.910 0.790 ;
        RECT  2.840 0.870 2.910 1.060 ;
        RECT  2.460 0.195 2.880 0.265 ;
        RECT  2.600 0.345 2.840 0.415 ;
        RECT  2.740 0.870 2.840 0.940 ;
        RECT  2.700 0.520 2.770 0.795 ;
        RECT  2.670 0.865 2.740 0.940 ;
        RECT  2.230 0.725 2.700 0.795 ;
        RECT  2.110 0.865 2.670 0.935 ;
        RECT  2.530 0.345 2.600 0.640 ;
        RECT  2.390 0.195 2.460 0.615 ;
        RECT  2.310 0.545 2.390 0.615 ;
        RECT  2.250 0.260 2.320 0.440 ;
        RECT  2.230 0.370 2.250 0.440 ;
        RECT  2.160 0.370 2.230 0.795 ;
        RECT  1.205 0.210 2.170 0.280 ;
        RECT  1.970 1.005 2.150 1.075 ;
        RECT  2.040 0.850 2.110 0.935 ;
        RECT  1.995 0.350 2.065 0.780 ;
        RECT  1.115 0.850 2.040 0.920 ;
        RECT  1.870 0.350 1.995 0.420 ;
        RECT  1.860 0.680 1.995 0.780 ;
        RECT  1.900 0.990 1.970 1.075 ;
        RECT  0.810 0.990 1.900 1.060 ;
        RECT  1.790 0.540 1.840 0.610 ;
        RECT  1.720 0.355 1.790 0.780 ;
        RECT  1.470 0.355 1.720 0.425 ;
        RECT  1.470 0.710 1.720 0.780 ;
        RECT  1.065 0.350 1.230 0.420 ;
        RECT  1.135 0.200 1.205 0.280 ;
        RECT  0.750 0.200 1.135 0.270 ;
        RECT  1.045 0.520 1.115 0.920 ;
        RECT  0.995 0.340 1.065 0.420 ;
        RECT  0.485 0.340 0.995 0.410 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.800 0.810 1.060 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCND4BWP

MACRO EDFKCNQD1BWP
    CLASS CORE ;
    FOREIGN EDFKCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.185 4.165 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.645 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.970 -0.115 4.200 0.115 ;
        RECT  3.850 -0.115 3.970 0.140 ;
        RECT  3.600 -0.115 3.850 0.115 ;
        RECT  3.480 -0.115 3.600 0.140 ;
        RECT  2.755 -0.115 3.480 0.115 ;
        RECT  2.685 -0.115 2.755 0.420 ;
        RECT  1.800 -0.115 2.685 0.115 ;
        RECT  1.680 -0.115 1.800 0.125 ;
        RECT  1.440 -0.115 1.680 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  0.330 -0.115 1.320 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.970 1.145 4.200 1.375 ;
        RECT  3.850 1.130 3.970 1.375 ;
        RECT  3.600 1.145 3.850 1.375 ;
        RECT  3.480 1.130 3.600 1.375 ;
        RECT  2.760 1.145 3.480 1.375 ;
        RECT  2.635 1.020 2.760 1.375 ;
        RECT  1.800 1.145 2.635 1.375 ;
        RECT  1.680 1.135 1.800 1.375 ;
        RECT  1.220 1.145 1.680 1.375 ;
        RECT  1.100 1.120 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.935 0.210 4.005 1.060 ;
        RECT  3.380 0.210 3.935 0.280 ;
        RECT  2.920 0.990 3.935 1.060 ;
        RECT  3.795 0.375 3.865 0.870 ;
        RECT  3.520 0.375 3.795 0.445 ;
        RECT  3.660 0.800 3.795 0.870 ;
        RECT  3.560 0.545 3.680 0.640 ;
        RECT  3.480 0.570 3.560 0.640 ;
        RECT  3.450 0.375 3.520 0.485 ;
        RECT  3.410 0.570 3.480 0.920 ;
        RECT  3.350 0.415 3.450 0.485 ;
        RECT  3.240 0.570 3.410 0.640 ;
        RECT  3.030 0.850 3.410 0.920 ;
        RECT  3.310 0.210 3.380 0.330 ;
        RECT  3.090 0.710 3.310 0.780 ;
        RECT  3.170 0.220 3.240 0.640 ;
        RECT  3.090 0.220 3.170 0.290 ;
        RECT  3.020 0.370 3.090 0.780 ;
        RECT  2.880 0.210 2.950 0.790 ;
        RECT  2.850 0.870 2.920 1.060 ;
        RECT  2.660 0.720 2.880 0.790 ;
        RECT  2.465 0.870 2.850 0.940 ;
        RECT  2.740 0.510 2.810 0.640 ;
        RECT  2.390 0.510 2.740 0.580 ;
        RECT  2.540 0.670 2.660 0.790 ;
        RECT  2.395 0.855 2.465 0.940 ;
        RECT  1.710 0.855 2.395 0.925 ;
        RECT  2.315 0.300 2.390 0.775 ;
        RECT  2.250 0.705 2.315 0.775 ;
        RECT  0.750 0.200 2.220 0.270 ;
        RECT  2.060 0.995 2.180 1.075 ;
        RECT  2.085 0.355 2.155 0.775 ;
        RECT  1.890 0.355 2.085 0.425 ;
        RECT  1.890 0.705 2.085 0.775 ;
        RECT  1.540 0.995 2.060 1.065 ;
        RECT  1.785 0.545 1.910 0.615 ;
        RECT  1.715 0.355 1.785 0.770 ;
        RECT  1.470 0.355 1.715 0.425 ;
        RECT  1.470 0.700 1.715 0.770 ;
        RECT  1.640 0.840 1.710 0.925 ;
        RECT  1.115 0.840 1.640 0.910 ;
        RECT  1.470 0.980 1.540 1.065 ;
        RECT  0.810 0.980 1.470 1.050 ;
        RECT  0.485 0.340 1.230 0.410 ;
        RECT  1.045 0.520 1.115 0.910 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.790 0.810 1.050 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCNQD1BWP

MACRO EDFKCNQD2BWP
    CLASS CORE ;
    FOREIGN EDFKCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.905 ;
        RECT  4.235 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.235 0.465 ;
        RECT  4.175 0.735 4.235 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.645 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 -0.115 4.480 0.115 ;
        RECT  4.355 -0.115 4.425 0.300 ;
        RECT  4.090 -0.115 4.355 0.115 ;
        RECT  3.970 -0.115 4.090 0.275 ;
        RECT  3.640 -0.115 3.970 0.115 ;
        RECT  3.640 0.215 3.730 0.285 ;
        RECT  3.520 -0.115 3.640 0.285 ;
        RECT  2.735 -0.115 3.520 0.115 ;
        RECT  3.430 0.215 3.520 0.285 ;
        RECT  2.665 -0.115 2.735 0.420 ;
        RECT  1.780 -0.115 2.665 0.115 ;
        RECT  1.660 -0.115 1.780 0.125 ;
        RECT  1.440 -0.115 1.660 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  0.330 -0.115 1.320 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 1.145 4.480 1.375 ;
        RECT  4.355 0.960 4.425 1.375 ;
        RECT  3.720 1.145 4.355 1.375 ;
        RECT  3.600 1.005 3.720 1.375 ;
        RECT  2.740 1.145 3.600 1.375 ;
        RECT  2.615 1.020 2.740 1.375 ;
        RECT  1.780 1.145 2.615 1.375 ;
        RECT  1.660 1.135 1.780 1.375 ;
        RECT  1.220 1.145 1.660 1.375 ;
        RECT  1.100 1.120 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.520 4.130 0.640 ;
        RECT  4.000 0.365 4.070 0.940 ;
        RECT  3.900 0.365 4.000 0.435 ;
        RECT  3.790 0.870 4.000 0.940 ;
        RECT  3.800 0.190 3.900 0.435 ;
        RECT  3.745 0.520 3.815 0.800 ;
        RECT  3.630 0.365 3.800 0.435 ;
        RECT  3.670 0.730 3.745 0.800 ;
        RECT  3.600 0.730 3.670 0.925 ;
        RECT  3.560 0.365 3.630 0.620 ;
        RECT  3.350 0.855 3.600 0.925 ;
        RECT  2.900 0.995 3.510 1.065 ;
        RECT  3.420 0.365 3.490 0.770 ;
        RECT  3.350 0.365 3.420 0.435 ;
        RECT  3.280 0.200 3.350 0.435 ;
        RECT  3.280 0.520 3.350 0.925 ;
        RECT  3.210 0.520 3.280 0.590 ;
        RECT  3.010 0.855 3.280 0.925 ;
        RECT  3.140 0.190 3.210 0.590 ;
        RECT  3.070 0.660 3.210 0.780 ;
        RECT  3.030 0.190 3.140 0.260 ;
        RECT  3.000 0.340 3.070 0.780 ;
        RECT  2.860 0.190 2.930 0.790 ;
        RECT  2.830 0.870 2.900 1.065 ;
        RECT  2.640 0.720 2.860 0.790 ;
        RECT  2.445 0.870 2.830 0.940 ;
        RECT  2.720 0.510 2.790 0.640 ;
        RECT  2.370 0.510 2.720 0.580 ;
        RECT  2.520 0.670 2.640 0.790 ;
        RECT  2.375 0.855 2.445 0.940 ;
        RECT  1.710 0.855 2.375 0.925 ;
        RECT  2.295 0.300 2.370 0.775 ;
        RECT  2.230 0.705 2.295 0.775 ;
        RECT  0.750 0.200 2.200 0.270 ;
        RECT  2.040 0.995 2.160 1.075 ;
        RECT  2.065 0.355 2.135 0.775 ;
        RECT  1.870 0.355 2.065 0.425 ;
        RECT  1.870 0.705 2.065 0.775 ;
        RECT  1.540 0.995 2.040 1.065 ;
        RECT  1.785 0.545 1.890 0.615 ;
        RECT  1.715 0.355 1.785 0.770 ;
        RECT  1.490 0.355 1.715 0.425 ;
        RECT  1.490 0.700 1.715 0.770 ;
        RECT  1.640 0.840 1.710 0.925 ;
        RECT  1.115 0.840 1.640 0.910 ;
        RECT  1.470 0.980 1.540 1.065 ;
        RECT  0.810 0.980 1.470 1.050 ;
        RECT  0.485 0.340 1.230 0.410 ;
        RECT  1.045 0.520 1.115 0.910 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.790 0.810 1.050 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCNQD2BWP

MACRO EDFKCNQD4BWP
    CLASS CORE ;
    FOREIGN EDFKCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.595 0.185 4.665 0.465 ;
        RECT  4.595 0.775 4.665 1.075 ;
        RECT  4.515 0.355 4.595 0.465 ;
        RECT  4.515 0.775 4.595 0.905 ;
        RECT  4.305 0.355 4.515 0.905 ;
        RECT  4.235 0.185 4.305 0.465 ;
        RECT  4.235 0.775 4.305 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0428 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.620 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.650 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.245 0.495 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.465 ;
        RECT  4.510 -0.115 4.775 0.115 ;
        RECT  4.390 -0.115 4.510 0.280 ;
        RECT  4.140 -0.115 4.390 0.115 ;
        RECT  4.020 -0.115 4.140 0.275 ;
        RECT  3.680 -0.115 4.020 0.115 ;
        RECT  3.680 0.215 3.770 0.285 ;
        RECT  3.560 -0.115 3.680 0.285 ;
        RECT  2.775 -0.115 3.560 0.115 ;
        RECT  3.470 0.215 3.560 0.285 ;
        RECT  2.705 -0.115 2.775 0.420 ;
        RECT  1.800 -0.115 2.705 0.115 ;
        RECT  1.680 -0.115 1.800 0.140 ;
        RECT  1.430 -0.115 1.680 0.115 ;
        RECT  1.310 -0.115 1.430 0.140 ;
        RECT  0.330 -0.115 1.310 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.680 4.845 1.375 ;
        RECT  4.510 1.145 4.775 1.375 ;
        RECT  4.390 0.975 4.510 1.375 ;
        RECT  4.140 1.145 4.390 1.375 ;
        RECT  4.020 1.030 4.140 1.375 ;
        RECT  3.760 1.145 4.020 1.375 ;
        RECT  3.640 1.005 3.760 1.375 ;
        RECT  2.780 1.145 3.640 1.375 ;
        RECT  2.655 1.020 2.780 1.375 ;
        RECT  1.800 1.145 2.655 1.375 ;
        RECT  1.680 1.130 1.800 1.375 ;
        RECT  1.220 1.145 1.680 1.375 ;
        RECT  1.100 1.130 1.220 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.595 0.185 4.665 0.465 ;
        RECT  4.595 0.775 4.665 1.075 ;
        RECT  4.585 0.355 4.595 0.465 ;
        RECT  4.585 0.775 4.595 0.905 ;
        RECT  4.090 0.520 4.190 0.640 ;
        RECT  4.020 0.365 4.090 0.960 ;
        RECT  3.940 0.365 4.020 0.435 ;
        RECT  3.830 0.890 4.020 0.960 ;
        RECT  3.840 0.190 3.940 0.435 ;
        RECT  3.855 0.520 3.925 0.820 ;
        RECT  3.710 0.750 3.855 0.820 ;
        RECT  3.670 0.365 3.840 0.435 ;
        RECT  3.640 0.750 3.710 0.925 ;
        RECT  3.600 0.365 3.670 0.620 ;
        RECT  3.390 0.855 3.640 0.925 ;
        RECT  2.940 0.995 3.550 1.065 ;
        RECT  3.460 0.365 3.530 0.770 ;
        RECT  3.390 0.365 3.460 0.435 ;
        RECT  3.320 0.200 3.390 0.435 ;
        RECT  3.320 0.520 3.390 0.925 ;
        RECT  3.250 0.520 3.320 0.590 ;
        RECT  3.050 0.855 3.320 0.925 ;
        RECT  3.180 0.190 3.250 0.590 ;
        RECT  3.110 0.660 3.250 0.780 ;
        RECT  3.070 0.190 3.180 0.260 ;
        RECT  3.040 0.340 3.110 0.780 ;
        RECT  2.900 0.190 2.970 0.790 ;
        RECT  2.870 0.870 2.940 1.065 ;
        RECT  2.680 0.720 2.900 0.790 ;
        RECT  2.465 0.870 2.870 0.940 ;
        RECT  2.760 0.510 2.830 0.640 ;
        RECT  2.390 0.510 2.760 0.580 ;
        RECT  2.560 0.670 2.680 0.790 ;
        RECT  2.395 0.850 2.465 0.940 ;
        RECT  1.115 0.850 2.395 0.920 ;
        RECT  2.315 0.300 2.390 0.775 ;
        RECT  2.250 0.705 2.315 0.775 ;
        RECT  1.205 0.210 2.220 0.280 ;
        RECT  2.050 0.990 2.170 1.070 ;
        RECT  2.085 0.355 2.155 0.780 ;
        RECT  1.870 0.355 2.085 0.425 ;
        RECT  1.870 0.710 2.085 0.780 ;
        RECT  0.810 0.990 2.050 1.060 ;
        RECT  1.790 0.545 1.890 0.615 ;
        RECT  1.720 0.355 1.790 0.780 ;
        RECT  1.490 0.355 1.720 0.425 ;
        RECT  1.490 0.710 1.720 0.780 ;
        RECT  1.065 0.350 1.230 0.420 ;
        RECT  1.135 0.200 1.205 0.280 ;
        RECT  0.750 0.200 1.135 0.270 ;
        RECT  1.045 0.520 1.115 0.920 ;
        RECT  0.995 0.340 1.065 0.420 ;
        RECT  0.485 0.340 0.995 0.410 ;
        RECT  0.845 0.480 0.915 0.620 ;
        RECT  0.415 0.480 0.845 0.550 ;
        RECT  0.740 0.800 0.810 1.060 ;
        RECT  0.415 0.195 0.485 0.410 ;
        RECT  0.345 0.480 0.415 0.920 ;
        RECT  0.330 0.480 0.345 0.550 ;
        RECT  0.125 0.850 0.345 0.920 ;
        RECT  0.260 0.355 0.330 0.550 ;
        RECT  0.125 0.355 0.260 0.425 ;
        RECT  0.055 0.270 0.125 0.425 ;
        RECT  0.055 0.850 0.125 1.040 ;
    END
END EDFKCNQD4BWP

MACRO EDFQD1BWP
    CLASS CORE ;
    FOREIGN EDFQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.185 3.745 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.225 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 -0.115 3.780 0.115 ;
        RECT  3.440 -0.115 3.560 0.140 ;
        RECT  3.200 -0.115 3.440 0.115 ;
        RECT  3.080 -0.115 3.200 0.140 ;
        RECT  2.375 -0.115 3.080 0.115 ;
        RECT  2.305 -0.115 2.375 0.420 ;
        RECT  1.440 -0.115 2.305 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.145 3.780 1.375 ;
        RECT  3.440 1.130 3.560 1.375 ;
        RECT  3.200 1.145 3.440 1.375 ;
        RECT  3.080 1.130 3.200 1.375 ;
        RECT  2.400 1.145 3.080 1.375 ;
        RECT  2.275 1.020 2.400 1.375 ;
        RECT  1.420 1.145 2.275 1.375 ;
        RECT  1.300 1.135 1.420 1.375 ;
        RECT  1.120 1.145 1.300 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.515 0.210 3.585 1.060 ;
        RECT  2.990 0.210 3.515 0.280 ;
        RECT  2.540 0.990 3.515 1.060 ;
        RECT  3.375 0.375 3.445 0.870 ;
        RECT  3.120 0.375 3.375 0.445 ;
        RECT  3.260 0.800 3.375 0.870 ;
        RECT  3.160 0.545 3.280 0.640 ;
        RECT  3.080 0.570 3.160 0.640 ;
        RECT  3.050 0.375 3.120 0.485 ;
        RECT  3.010 0.570 3.080 0.920 ;
        RECT  2.950 0.415 3.050 0.485 ;
        RECT  2.850 0.570 3.010 0.640 ;
        RECT  2.670 0.850 3.010 0.920 ;
        RECT  2.920 0.210 2.990 0.330 ;
        RECT  2.710 0.710 2.930 0.780 ;
        RECT  2.780 0.220 2.850 0.640 ;
        RECT  2.690 0.220 2.780 0.290 ;
        RECT  2.640 0.370 2.710 0.780 ;
        RECT  2.500 0.210 2.570 0.790 ;
        RECT  2.470 0.870 2.540 1.060 ;
        RECT  2.280 0.720 2.500 0.790 ;
        RECT  2.085 0.870 2.470 0.940 ;
        RECT  2.360 0.510 2.430 0.640 ;
        RECT  2.010 0.510 2.360 0.580 ;
        RECT  2.160 0.670 2.280 0.790 ;
        RECT  2.015 0.855 2.085 0.940 ;
        RECT  1.020 0.855 2.015 0.925 ;
        RECT  1.935 0.300 2.010 0.775 ;
        RECT  1.870 0.705 1.935 0.775 ;
        RECT  0.620 0.195 1.840 0.265 ;
        RECT  1.680 0.995 1.800 1.075 ;
        RECT  1.705 0.335 1.775 0.785 ;
        RECT  1.530 0.335 1.705 0.405 ;
        RECT  1.510 0.715 1.705 0.785 ;
        RECT  0.610 0.995 1.680 1.065 ;
        RECT  1.375 0.545 1.550 0.615 ;
        RECT  1.305 0.335 1.375 0.785 ;
        RECT  1.170 0.335 1.305 0.405 ;
        RECT  1.150 0.715 1.305 0.785 ;
        RECT  0.900 0.695 1.020 0.925 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFQD1BWP

MACRO EDFQD2BWP
    CLASS CORE ;
    FOREIGN EDFQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 0.355 3.885 0.905 ;
        RECT  3.825 0.185 3.830 0.905 ;
        RECT  3.810 0.185 3.825 1.035 ;
        RECT  3.760 0.185 3.810 0.465 ;
        RECT  3.755 0.735 3.810 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.545 1.225 0.625 ;
        RECT  1.015 0.355 1.085 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.305 ;
        RECT  3.650 -0.115 3.935 0.115 ;
        RECT  3.530 -0.115 3.650 0.140 ;
        RECT  3.280 -0.115 3.530 0.115 ;
        RECT  3.160 -0.115 3.280 0.130 ;
        RECT  2.375 -0.115 3.160 0.115 ;
        RECT  2.305 -0.115 2.375 0.420 ;
        RECT  1.440 -0.115 2.305 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.305 -0.115 1.020 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.145 4.060 1.375 ;
        RECT  3.935 0.960 4.005 1.375 ;
        RECT  3.610 1.145 3.935 1.375 ;
        RECT  3.490 1.110 3.610 1.375 ;
        RECT  3.220 1.145 3.490 1.375 ;
        RECT  3.100 1.135 3.220 1.375 ;
        RECT  2.400 1.145 3.100 1.375 ;
        RECT  2.275 1.020 2.400 1.375 ;
        RECT  1.420 1.145 2.275 1.375 ;
        RECT  1.300 1.135 1.420 1.375 ;
        RECT  1.120 1.145 1.300 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.680 0.520 3.710 0.640 ;
        RECT  3.610 0.255 3.680 0.975 ;
        RECT  3.180 0.255 3.610 0.325 ;
        RECT  3.310 0.905 3.610 0.975 ;
        RECT  3.470 0.410 3.540 0.820 ;
        RECT  3.030 0.410 3.470 0.480 ;
        RECT  3.210 0.750 3.470 0.820 ;
        RECT  3.070 0.550 3.360 0.620 ;
        RECT  3.140 0.750 3.210 1.065 ;
        RECT  3.110 0.215 3.180 0.325 ;
        RECT  2.540 0.995 3.140 1.065 ;
        RECT  3.030 0.215 3.110 0.285 ;
        RECT  3.000 0.550 3.070 0.925 ;
        RECT  2.960 0.360 3.030 0.480 ;
        RECT  2.860 0.550 3.000 0.620 ;
        RECT  2.670 0.855 3.000 0.925 ;
        RECT  2.710 0.715 2.920 0.785 ;
        RECT  2.790 0.220 2.860 0.620 ;
        RECT  2.710 0.220 2.790 0.290 ;
        RECT  2.640 0.370 2.710 0.785 ;
        RECT  2.500 0.210 2.570 0.790 ;
        RECT  2.470 0.870 2.540 1.065 ;
        RECT  2.280 0.720 2.500 0.790 ;
        RECT  2.085 0.870 2.470 0.940 ;
        RECT  2.360 0.510 2.430 0.640 ;
        RECT  2.010 0.510 2.360 0.580 ;
        RECT  2.160 0.670 2.280 0.790 ;
        RECT  2.015 0.855 2.085 0.940 ;
        RECT  1.020 0.855 2.015 0.925 ;
        RECT  1.935 0.300 2.010 0.775 ;
        RECT  1.870 0.705 1.935 0.775 ;
        RECT  0.620 0.195 1.840 0.265 ;
        RECT  1.680 0.995 1.800 1.075 ;
        RECT  1.705 0.335 1.775 0.785 ;
        RECT  1.530 0.335 1.705 0.405 ;
        RECT  1.510 0.715 1.705 0.785 ;
        RECT  0.610 0.995 1.680 1.065 ;
        RECT  1.375 0.545 1.550 0.615 ;
        RECT  1.305 0.335 1.375 0.785 ;
        RECT  1.170 0.335 1.305 0.405 ;
        RECT  1.150 0.715 1.305 0.785 ;
        RECT  0.900 0.695 1.020 0.925 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFQD2BWP

MACRO EDFQD4BWP
    CLASS CORE ;
    FOREIGN EDFQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.185 4.245 0.465 ;
        RECT  4.235 0.775 4.245 1.075 ;
        RECT  4.175 0.185 4.235 1.075 ;
        RECT  4.025 0.355 4.175 0.905 ;
        RECT  3.885 0.355 4.025 0.465 ;
        RECT  3.885 0.775 4.025 0.905 ;
        RECT  3.815 0.185 3.885 0.465 ;
        RECT  3.815 0.775 3.885 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.530 1.225 0.630 ;
        RECT  1.015 0.355 1.085 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 -0.115 4.480 0.115 ;
        RECT  4.355 -0.115 4.425 0.465 ;
        RECT  4.090 -0.115 4.355 0.115 ;
        RECT  3.970 -0.115 4.090 0.275 ;
        RECT  3.720 -0.115 3.970 0.115 ;
        RECT  3.600 -0.115 3.720 0.140 ;
        RECT  3.340 -0.115 3.600 0.115 ;
        RECT  3.220 -0.115 3.340 0.130 ;
        RECT  2.435 -0.115 3.220 0.115 ;
        RECT  2.365 -0.115 2.435 0.420 ;
        RECT  1.480 -0.115 2.365 0.115 ;
        RECT  1.360 -0.115 1.480 0.140 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.140 ;
        RECT  0.305 -0.115 1.000 0.115 ;
        RECT  0.235 -0.115 0.305 0.330 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.425 1.145 4.480 1.375 ;
        RECT  4.355 0.680 4.425 1.375 ;
        RECT  4.065 1.145 4.355 1.375 ;
        RECT  3.995 0.975 4.065 1.375 ;
        RECT  3.700 1.145 3.995 1.375 ;
        RECT  3.580 1.110 3.700 1.375 ;
        RECT  3.280 1.145 3.580 1.375 ;
        RECT  3.160 1.135 3.280 1.375 ;
        RECT  2.460 1.145 3.160 1.375 ;
        RECT  2.335 1.020 2.460 1.375 ;
        RECT  1.480 1.145 2.335 1.375 ;
        RECT  1.360 1.130 1.480 1.375 ;
        RECT  1.110 1.145 1.360 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.355 3.955 0.465 ;
        RECT  3.885 0.775 3.955 0.905 ;
        RECT  3.815 0.185 3.885 0.465 ;
        RECT  3.815 0.775 3.885 1.075 ;
        RECT  3.740 0.545 3.850 0.615 ;
        RECT  3.670 0.255 3.740 0.975 ;
        RECT  3.240 0.255 3.670 0.325 ;
        RECT  3.370 0.905 3.670 0.975 ;
        RECT  3.530 0.410 3.600 0.820 ;
        RECT  3.090 0.410 3.530 0.480 ;
        RECT  3.270 0.750 3.530 0.820 ;
        RECT  3.130 0.550 3.440 0.620 ;
        RECT  3.200 0.750 3.270 1.065 ;
        RECT  3.170 0.215 3.240 0.325 ;
        RECT  2.600 0.995 3.200 1.065 ;
        RECT  3.090 0.215 3.170 0.285 ;
        RECT  3.060 0.550 3.130 0.925 ;
        RECT  3.020 0.360 3.090 0.480 ;
        RECT  2.920 0.550 3.060 0.620 ;
        RECT  2.730 0.855 3.060 0.925 ;
        RECT  2.770 0.715 2.980 0.785 ;
        RECT  2.850 0.220 2.920 0.620 ;
        RECT  2.770 0.220 2.850 0.290 ;
        RECT  2.700 0.370 2.770 0.785 ;
        RECT  2.560 0.210 2.630 0.790 ;
        RECT  2.530 0.870 2.600 1.065 ;
        RECT  2.340 0.720 2.560 0.790 ;
        RECT  2.145 0.870 2.530 0.940 ;
        RECT  2.420 0.510 2.490 0.640 ;
        RECT  2.070 0.510 2.420 0.580 ;
        RECT  2.220 0.670 2.340 0.790 ;
        RECT  2.075 0.850 2.145 0.940 ;
        RECT  1.020 0.850 2.075 0.920 ;
        RECT  1.995 0.300 2.070 0.770 ;
        RECT  1.930 0.700 1.995 0.770 ;
        RECT  0.920 0.210 1.900 0.280 ;
        RECT  0.920 0.990 1.850 1.060 ;
        RECT  1.725 0.350 1.795 0.780 ;
        RECT  1.550 0.350 1.725 0.420 ;
        RECT  1.550 0.710 1.725 0.780 ;
        RECT  1.460 0.545 1.570 0.615 ;
        RECT  1.390 0.350 1.460 0.780 ;
        RECT  1.170 0.350 1.390 0.420 ;
        RECT  1.170 0.710 1.390 0.780 ;
        RECT  0.900 0.700 1.020 0.920 ;
        RECT  0.850 0.195 0.920 0.280 ;
        RECT  0.850 0.990 0.920 1.065 ;
        RECT  0.620 0.195 0.850 0.265 ;
        RECT  0.610 0.995 0.850 1.065 ;
        RECT  0.735 0.490 0.810 0.920 ;
        RECT  0.125 0.850 0.735 0.920 ;
        RECT  0.595 0.355 0.665 0.780 ;
        RECT  0.410 0.355 0.595 0.425 ;
        RECT  0.410 0.710 0.595 0.780 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.105 0.850 0.125 1.050 ;
        RECT  0.035 0.210 0.105 1.050 ;
    END
END EDFQD4BWP

MACRO FA1D0BWP
    CLASS CORE ;
    FOREIGN FA1D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.045 0.325 3.100 0.395 ;
        RECT  2.970 0.325 3.045 0.780 ;
        RECT  2.940 0.680 2.970 0.780 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.290 3.465 0.905 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.545 2.830 0.625 ;
        RECT  2.695 0.355 2.765 0.625 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0472 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.110 0.495 1.155 0.640 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.115 3.500 0.115 ;
        RECT  3.180 -0.115 3.260 0.420 ;
        RECT  2.700 -0.115 3.180 0.115 ;
        RECT  2.580 -0.115 2.700 0.125 ;
        RECT  1.280 -0.115 2.580 0.115 ;
        RECT  1.160 -0.115 1.280 0.140 ;
        RECT  0.330 -0.115 1.160 0.115 ;
        RECT  0.210 -0.115 0.330 0.255 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.145 3.500 1.375 ;
        RECT  3.130 1.135 3.250 1.375 ;
        RECT  2.660 1.145 3.130 1.375 ;
        RECT  2.540 1.135 2.660 1.375 ;
        RECT  1.270 1.145 2.540 1.375 ;
        RECT  1.150 1.010 1.270 1.375 ;
        RECT  0.330 1.145 1.150 1.375 ;
        RECT  0.210 1.030 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.825 0.995 3.410 1.065 ;
        RECT  3.115 0.520 3.190 0.925 ;
        RECT  2.230 0.855 3.115 0.925 ;
        RECT  2.610 0.205 2.910 0.275 ;
        RECT  2.610 0.695 2.870 0.785 ;
        RECT  2.540 0.205 2.610 0.785 ;
        RECT  2.085 0.205 2.540 0.275 ;
        RECT  2.515 0.520 2.540 0.640 ;
        RECT  2.440 0.345 2.460 0.465 ;
        RECT  2.370 0.345 2.440 0.770 ;
        RECT  2.310 0.700 2.370 0.770 ;
        RECT  2.230 0.350 2.290 0.420 ;
        RECT  2.160 0.350 2.230 0.925 ;
        RECT  2.080 0.855 2.160 0.925 ;
        RECT  2.015 0.205 2.085 0.615 ;
        RECT  1.975 0.545 2.015 0.615 ;
        RECT  1.905 0.545 1.975 0.915 ;
        RECT  1.825 0.350 1.910 0.420 ;
        RECT  1.755 0.350 1.825 1.065 ;
        RECT  1.715 0.905 1.755 1.065 ;
        RECT  1.645 0.325 1.680 0.780 ;
        RECT  1.610 0.325 1.645 0.940 ;
        RECT  1.590 0.325 1.610 0.445 ;
        RECT  1.575 0.710 1.610 0.940 ;
        RECT  1.065 0.870 1.575 0.940 ;
        RECT  1.505 0.515 1.535 0.635 ;
        RECT  1.435 0.210 1.505 0.800 ;
        RECT  1.350 0.210 1.435 0.280 ;
        RECT  1.330 0.730 1.435 0.800 ;
        RECT  1.295 0.350 1.365 0.640 ;
        RECT  1.240 0.350 1.295 0.420 ;
        RECT  1.170 0.210 1.240 0.420 ;
        RECT  0.685 0.210 1.170 0.280 ;
        RECT  1.040 0.350 1.090 0.420 ;
        RECT  1.040 0.735 1.065 1.035 ;
        RECT  0.995 0.350 1.040 1.035 ;
        RECT  0.970 0.350 0.995 0.805 ;
        RECT  0.920 0.520 0.970 0.640 ;
        RECT  0.850 0.350 0.890 0.450 ;
        RECT  0.860 0.760 0.890 0.880 ;
        RECT  0.850 0.760 0.860 1.055 ;
        RECT  0.780 0.350 0.850 1.055 ;
        RECT  0.500 0.985 0.780 1.055 ;
        RECT  0.615 0.210 0.685 0.915 ;
        RECT  0.485 0.395 0.530 0.820 ;
        RECT  0.430 0.890 0.500 1.055 ;
        RECT  0.460 0.185 0.485 0.820 ;
        RECT  0.415 0.185 0.460 0.465 ;
        RECT  0.415 0.700 0.460 0.820 ;
        RECT  0.330 0.890 0.430 0.960 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.345 0.330 0.960 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.890 0.260 0.960 ;
        RECT  0.055 0.240 0.125 0.415 ;
        RECT  0.055 0.890 0.125 1.035 ;
    END
END FA1D0BWP

MACRO FA1D1BWP
    CLASS CORE ;
    FOREIGN FA1D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.215 3.885 0.485 ;
        RECT  3.800 0.215 3.870 0.800 ;
        RECT  3.670 0.215 3.800 0.285 ;
        RECT  3.680 0.700 3.800 0.800 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.045 ;
        RECT  4.075 0.185 4.095 0.465 ;
        RECT  4.080 0.730 4.095 1.045 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.355 3.465 0.625 ;
        RECT  3.340 0.540 3.395 0.625 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0480 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.000 0.625 ;
        RECT  0.875 0.355 0.945 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.270 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.985 -0.115 4.200 0.115 ;
        RECT  3.865 -0.115 3.985 0.140 ;
        RECT  3.610 -0.115 3.865 0.115 ;
        RECT  3.490 -0.115 3.610 0.140 ;
        RECT  3.220 -0.115 3.490 0.115 ;
        RECT  3.100 -0.115 3.220 0.135 ;
        RECT  1.845 -0.115 3.100 0.115 ;
        RECT  1.725 -0.115 1.845 0.130 ;
        RECT  0.890 -0.115 1.725 0.115 ;
        RECT  0.770 -0.115 0.890 0.135 ;
        RECT  0.485 -0.115 0.770 0.115 ;
        RECT  0.415 -0.115 0.485 0.305 ;
        RECT  0.140 -0.115 0.415 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.145 4.200 1.375 ;
        RECT  3.860 1.010 3.980 1.375 ;
        RECT  3.610 1.145 3.860 1.375 ;
        RECT  3.490 1.130 3.610 1.375 ;
        RECT  3.200 1.145 3.490 1.375 ;
        RECT  3.080 1.130 3.200 1.375 ;
        RECT  1.820 1.145 3.080 1.375 ;
        RECT  1.700 1.030 1.820 1.375 ;
        RECT  0.890 1.145 1.700 1.375 ;
        RECT  0.770 1.120 0.890 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.010 0.515 4.025 0.640 ;
        RECT  3.955 0.515 4.010 0.940 ;
        RECT  3.940 0.595 3.955 0.940 ;
        RECT  3.780 0.870 3.940 0.940 ;
        RECT  3.710 0.870 3.780 1.060 ;
        RECT  3.610 0.540 3.730 0.620 ;
        RECT  2.410 0.990 3.710 1.060 ;
        RECT  3.540 0.540 3.610 0.920 ;
        RECT  2.820 0.850 3.540 0.920 ;
        RECT  3.215 0.710 3.420 0.780 ;
        RECT  3.215 0.205 3.410 0.275 ;
        RECT  3.145 0.205 3.215 0.780 ;
        RECT  2.635 0.205 3.145 0.275 ;
        RECT  3.040 0.520 3.145 0.640 ;
        RECT  2.960 0.355 3.030 0.425 ;
        RECT  2.960 0.710 3.010 0.780 ;
        RECT  2.890 0.355 2.960 0.780 ;
        RECT  2.750 0.360 2.820 0.920 ;
        RECT  2.640 0.850 2.750 0.920 ;
        RECT  2.565 0.205 2.635 0.730 ;
        RECT  2.550 0.660 2.565 0.730 ;
        RECT  2.480 0.660 2.550 0.900 ;
        RECT  2.410 0.195 2.445 0.455 ;
        RECT  2.340 0.195 2.410 1.060 ;
        RECT  2.300 0.915 2.340 1.060 ;
        RECT  2.220 0.330 2.270 0.790 ;
        RECT  2.200 0.330 2.220 0.960 ;
        RECT  2.185 0.720 2.200 0.960 ;
        RECT  2.150 0.720 2.185 1.075 ;
        RECT  2.115 0.890 2.150 1.075 ;
        RECT  2.045 0.530 2.130 0.650 ;
        RECT  1.585 0.890 2.115 0.960 ;
        RECT  1.975 0.260 2.045 0.820 ;
        RECT  1.910 0.750 1.975 0.820 ;
        RECT  1.815 0.200 1.885 0.640 ;
        RECT  1.225 0.200 1.815 0.270 ;
        RECT  1.585 0.370 1.625 0.610 ;
        RECT  1.555 0.370 1.585 1.030 ;
        RECT  1.515 0.540 1.555 1.030 ;
        RECT  1.445 0.540 1.515 0.660 ;
        RECT  1.375 0.340 1.460 0.410 ;
        RECT  1.375 0.800 1.405 1.050 ;
        RECT  1.305 0.340 1.375 1.050 ;
        RECT  0.850 0.980 1.305 1.050 ;
        RECT  1.155 0.200 1.225 0.900 ;
        RECT  0.665 0.205 1.070 0.275 ;
        RECT  0.960 0.730 1.060 0.910 ;
        RECT  0.800 0.730 0.960 0.800 ;
        RECT  0.780 0.870 0.850 1.050 ;
        RECT  0.730 0.405 0.800 0.800 ;
        RECT  0.490 0.870 0.780 0.940 ;
        RECT  0.665 0.405 0.730 0.475 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.595 0.205 0.665 0.475 ;
        RECT  0.500 0.545 0.640 0.615 ;
        RECT  0.490 0.395 0.500 0.615 ;
        RECT  0.420 0.395 0.490 0.940 ;
        RECT  0.305 0.395 0.420 0.465 ;
        RECT  0.305 0.870 0.420 0.940 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FA1D1BWP

MACRO FA1D2BWP
    CLASS CORE ;
    FOREIGN FA1D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.185 3.745 0.820 ;
        RECT  3.655 0.185 3.675 0.465 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.105 0.355 4.165 0.805 ;
        RECT  4.095 0.185 4.105 1.035 ;
        RECT  4.035 0.185 4.095 0.465 ;
        RECT  4.035 0.735 4.095 1.035 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.545 3.375 0.630 ;
        RECT  3.255 0.355 3.325 0.630 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0480 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.000 0.625 ;
        RECT  0.875 0.355 0.945 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.270 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.115 4.340 0.115 ;
        RECT  4.215 -0.115 4.285 0.300 ;
        RECT  3.925 -0.115 4.215 0.115 ;
        RECT  3.855 -0.115 3.925 0.465 ;
        RECT  3.530 -0.115 3.855 0.115 ;
        RECT  3.460 -0.115 3.530 0.430 ;
        RECT  3.180 -0.115 3.460 0.115 ;
        RECT  3.060 -0.115 3.180 0.135 ;
        RECT  1.840 -0.115 3.060 0.115 ;
        RECT  1.720 -0.115 1.840 0.130 ;
        RECT  0.890 -0.115 1.720 0.115 ;
        RECT  0.770 -0.115 0.890 0.135 ;
        RECT  0.485 -0.115 0.770 0.115 ;
        RECT  0.415 -0.115 0.485 0.305 ;
        RECT  0.140 -0.115 0.415 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 1.145 4.340 1.375 ;
        RECT  4.215 0.905 4.285 1.375 ;
        RECT  3.950 1.145 4.215 1.375 ;
        RECT  3.830 1.030 3.950 1.375 ;
        RECT  3.560 1.145 3.830 1.375 ;
        RECT  3.440 1.130 3.560 1.375 ;
        RECT  3.160 1.145 3.440 1.375 ;
        RECT  3.040 1.130 3.160 1.375 ;
        RECT  1.790 1.145 3.040 1.375 ;
        RECT  1.670 1.030 1.790 1.375 ;
        RECT  0.890 1.145 1.670 1.375 ;
        RECT  0.770 1.120 0.890 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.930 0.545 4.020 0.615 ;
        RECT  3.860 0.545 3.930 0.960 ;
        RECT  3.750 0.890 3.860 0.960 ;
        RECT  3.680 0.890 3.750 1.060 ;
        RECT  2.370 0.990 3.680 1.060 ;
        RECT  3.585 0.520 3.605 0.640 ;
        RECT  3.515 0.520 3.585 0.920 ;
        RECT  2.780 0.850 3.515 0.920 ;
        RECT  3.155 0.205 3.370 0.275 ;
        RECT  3.155 0.710 3.360 0.780 ;
        RECT  3.085 0.205 3.155 0.780 ;
        RECT  2.610 0.205 3.085 0.275 ;
        RECT  3.000 0.520 3.085 0.640 ;
        RECT  2.930 0.355 2.990 0.425 ;
        RECT  2.860 0.355 2.930 0.780 ;
        RECT  2.710 0.360 2.780 0.920 ;
        RECT  2.600 0.850 2.710 0.920 ;
        RECT  2.540 0.205 2.610 0.730 ;
        RECT  2.510 0.660 2.540 0.730 ;
        RECT  2.440 0.660 2.510 0.900 ;
        RECT  2.370 0.195 2.405 0.455 ;
        RECT  2.300 0.195 2.370 1.060 ;
        RECT  2.240 0.915 2.300 1.060 ;
        RECT  2.170 0.330 2.230 0.790 ;
        RECT  2.160 0.330 2.170 0.960 ;
        RECT  2.125 0.720 2.160 0.960 ;
        RECT  2.100 0.720 2.125 1.075 ;
        RECT  2.055 0.890 2.100 1.075 ;
        RECT  2.020 0.530 2.080 0.650 ;
        RECT  1.585 0.890 2.055 0.960 ;
        RECT  1.950 0.195 2.020 0.820 ;
        RECT  1.850 0.750 1.950 0.820 ;
        RECT  1.810 0.200 1.880 0.640 ;
        RECT  1.225 0.200 1.810 0.270 ;
        RECT  1.585 0.370 1.625 0.610 ;
        RECT  1.555 0.370 1.585 1.030 ;
        RECT  1.515 0.540 1.555 1.030 ;
        RECT  1.445 0.540 1.515 0.660 ;
        RECT  1.375 0.340 1.460 0.410 ;
        RECT  1.375 0.800 1.405 1.050 ;
        RECT  1.305 0.340 1.375 1.050 ;
        RECT  0.850 0.980 1.305 1.050 ;
        RECT  1.155 0.200 1.225 0.900 ;
        RECT  0.665 0.205 1.070 0.275 ;
        RECT  0.960 0.730 1.060 0.910 ;
        RECT  0.800 0.730 0.960 0.800 ;
        RECT  0.780 0.870 0.850 1.050 ;
        RECT  0.730 0.405 0.800 0.800 ;
        RECT  0.490 0.870 0.780 0.940 ;
        RECT  0.665 0.405 0.730 0.475 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.595 0.205 0.665 0.475 ;
        RECT  0.500 0.545 0.640 0.615 ;
        RECT  0.490 0.395 0.500 0.615 ;
        RECT  0.420 0.395 0.490 0.940 ;
        RECT  0.305 0.395 0.420 0.465 ;
        RECT  0.305 0.870 0.420 0.940 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FA1D2BWP

MACRO FA1D4BWP
    CLASS CORE ;
    FOREIGN FA1D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.720 4.950 0.800 ;
        RECT  4.855 0.185 4.925 0.465 ;
        RECT  4.795 0.355 4.855 0.465 ;
        RECT  4.585 0.355 4.795 0.800 ;
        RECT  4.545 0.355 4.585 0.465 ;
        RECT  4.450 0.720 4.585 0.800 ;
        RECT  4.475 0.185 4.545 0.465 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.185 5.645 0.465 ;
        RECT  5.635 0.745 5.645 1.075 ;
        RECT  5.575 0.185 5.635 1.075 ;
        RECT  5.425 0.345 5.575 0.905 ;
        RECT  5.285 0.345 5.425 0.465 ;
        RECT  5.285 0.745 5.425 0.905 ;
        RECT  5.215 0.185 5.285 0.465 ;
        RECT  5.215 0.745 5.285 1.075 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 0.355 4.175 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.205 0.765 ;
        RECT  2.030 0.495 2.135 0.640 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.825 -0.115 5.880 0.115 ;
        RECT  5.755 -0.115 5.825 0.465 ;
        RECT  5.490 -0.115 5.755 0.115 ;
        RECT  5.370 -0.115 5.490 0.270 ;
        RECT  5.105 -0.115 5.370 0.115 ;
        RECT  5.035 -0.115 5.105 0.465 ;
        RECT  4.760 -0.115 5.035 0.115 ;
        RECT  4.640 -0.115 4.760 0.280 ;
        RECT  4.355 -0.115 4.640 0.115 ;
        RECT  4.285 -0.115 4.355 0.465 ;
        RECT  4.000 -0.115 4.285 0.115 ;
        RECT  3.880 -0.115 4.000 0.140 ;
        RECT  3.610 -0.115 3.880 0.115 ;
        RECT  3.490 -0.115 3.610 0.140 ;
        RECT  2.200 -0.115 3.490 0.115 ;
        RECT  2.080 -0.115 2.200 0.140 ;
        RECT  1.060 -0.115 2.080 0.115 ;
        RECT  0.940 -0.115 1.060 0.140 ;
        RECT  0.665 -0.115 0.940 0.115 ;
        RECT  0.595 -0.115 0.665 0.465 ;
        RECT  0.330 -0.115 0.595 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.825 1.145 5.880 1.375 ;
        RECT  5.755 0.680 5.825 1.375 ;
        RECT  5.490 1.145 5.755 1.375 ;
        RECT  5.370 0.975 5.490 1.375 ;
        RECT  5.130 1.145 5.370 1.375 ;
        RECT  5.010 1.010 5.130 1.375 ;
        RECT  4.760 1.145 5.010 1.375 ;
        RECT  4.640 1.010 4.760 1.375 ;
        RECT  4.380 1.145 4.640 1.375 ;
        RECT  4.260 1.130 4.380 1.375 ;
        RECT  3.980 1.145 4.260 1.375 ;
        RECT  3.860 1.130 3.980 1.375 ;
        RECT  3.530 1.145 3.860 1.375 ;
        RECT  3.410 1.130 3.530 1.375 ;
        RECT  2.200 1.145 3.410 1.375 ;
        RECT  2.080 1.030 2.200 1.375 ;
        RECT  1.060 1.145 2.080 1.375 ;
        RECT  0.940 1.120 1.060 1.375 ;
        RECT  0.690 1.145 0.940 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.025 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.345 5.355 0.465 ;
        RECT  5.285 0.745 5.355 0.905 ;
        RECT  5.215 0.185 5.285 0.465 ;
        RECT  5.215 0.745 5.285 1.075 ;
        RECT  4.865 0.720 4.950 0.800 ;
        RECT  4.865 0.185 4.925 0.465 ;
        RECT  4.475 0.185 4.515 0.465 ;
        RECT  4.450 0.720 4.515 0.800 ;
        RECT  5.105 0.545 5.260 0.615 ;
        RECT  5.035 0.545 5.105 0.940 ;
        RECT  4.550 0.870 5.035 0.940 ;
        RECT  4.480 0.870 4.550 1.060 ;
        RECT  4.370 0.545 4.500 0.615 ;
        RECT  2.780 0.990 4.480 1.060 ;
        RECT  4.300 0.545 4.370 0.920 ;
        RECT  3.085 0.850 4.300 0.920 ;
        RECT  3.980 0.210 4.190 0.280 ;
        RECT  3.980 0.710 4.190 0.780 ;
        RECT  3.910 0.210 3.980 0.780 ;
        RECT  3.025 0.210 3.910 0.280 ;
        RECT  3.590 0.545 3.910 0.615 ;
        RECT  3.365 0.350 3.810 0.420 ;
        RECT  3.365 0.710 3.780 0.780 ;
        RECT  3.295 0.350 3.365 0.780 ;
        RECT  3.230 0.710 3.295 0.780 ;
        RECT  3.145 0.350 3.215 0.570 ;
        RECT  3.085 0.500 3.145 0.570 ;
        RECT  3.015 0.500 3.085 0.920 ;
        RECT  2.955 0.210 3.025 0.420 ;
        RECT  2.930 0.350 2.955 0.420 ;
        RECT  2.860 0.350 2.930 0.910 ;
        RECT  2.710 0.320 2.780 1.060 ;
        RECT  2.680 0.870 2.710 1.060 ;
        RECT  2.600 0.370 2.630 0.780 ;
        RECT  2.560 0.370 2.600 0.960 ;
        RECT  2.510 0.370 2.560 0.440 ;
        RECT  2.530 0.710 2.560 0.960 ;
        RECT  1.960 0.890 2.530 0.960 ;
        RECT  2.400 0.185 2.520 0.280 ;
        RECT  2.405 0.520 2.480 0.640 ;
        RECT  2.385 0.350 2.405 0.640 ;
        RECT  1.585 0.210 2.400 0.280 ;
        RECT  2.335 0.350 2.385 0.820 ;
        RECT  2.315 0.520 2.335 0.820 ;
        RECT  1.960 0.350 2.010 0.420 ;
        RECT  1.890 0.350 1.960 1.035 ;
        RECT  1.875 0.520 1.890 1.035 ;
        RECT  1.815 0.520 1.875 0.640 ;
        RECT  1.735 0.360 1.820 0.430 ;
        RECT  1.735 0.745 1.760 0.865 ;
        RECT  1.665 0.360 1.735 1.050 ;
        RECT  0.850 0.980 1.665 1.050 ;
        RECT  1.515 0.210 1.585 0.910 ;
        RECT  1.375 0.375 1.445 0.770 ;
        RECT  1.050 0.210 1.430 0.280 ;
        RECT  1.050 0.840 1.430 0.910 ;
        RECT  1.130 0.375 1.375 0.445 ;
        RECT  1.130 0.700 1.375 0.770 ;
        RECT  0.980 0.210 1.050 0.910 ;
        RECT  0.845 0.395 0.980 0.465 ;
        RECT  0.750 0.725 0.980 0.795 ;
        RECT  0.485 0.545 0.870 0.615 ;
        RECT  0.780 0.865 0.850 1.050 ;
        RECT  0.775 0.185 0.845 0.465 ;
        RECT  0.485 0.865 0.780 0.935 ;
        RECT  0.415 0.185 0.485 1.015 ;
        RECT  0.125 0.345 0.415 0.415 ;
        RECT  0.125 0.865 0.415 0.935 ;
        RECT  0.055 0.230 0.125 0.415 ;
        RECT  0.055 0.865 0.125 1.015 ;
    END
END FA1D4BWP

MACRO FCICIND1BWP
    CLASS CORE ;
    FOREIGN FCICIND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.395 1.505 0.795 ;
        RECT  1.385 0.395 1.435 0.465 ;
        RECT  1.290 0.725 1.435 0.795 ;
        RECT  1.295 0.185 1.385 0.465 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.645 0.675 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.475 0.885 0.640 ;
        RECT  0.525 0.475 0.815 0.545 ;
        RECT  0.455 0.475 0.525 0.765 ;
        RECT  0.400 0.550 0.455 0.650 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 -0.115 1.820 0.115 ;
        RECT  1.500 -0.115 1.580 0.275 ;
        RECT  0.560 -0.115 1.500 0.115 ;
        RECT  0.440 -0.115 0.560 0.260 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.145 1.820 1.375 ;
        RECT  1.480 1.010 1.600 1.375 ;
        RECT  0.525 1.145 1.480 1.375 ;
        RECT  0.455 0.870 0.525 1.375 ;
        RECT  0.000 1.145 0.455 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.205 1.785 1.020 ;
        RECT  1.670 0.205 1.715 0.275 ;
        RECT  1.695 0.870 1.715 1.020 ;
        RECT  1.360 0.870 1.695 0.940 ;
        RECT  1.290 0.870 1.360 1.065 ;
        RECT  1.035 0.545 1.340 0.615 ;
        RECT  0.665 0.995 1.290 1.065 ;
        RECT  0.805 0.855 1.210 0.925 ;
        RECT  1.115 0.195 1.185 0.455 ;
        RECT  0.680 0.195 1.115 0.265 ;
        RECT  0.965 0.335 1.035 0.785 ;
        RECT  0.330 0.335 0.965 0.405 ;
        RECT  0.890 0.715 0.965 0.785 ;
        RECT  0.735 0.785 0.805 0.925 ;
        RECT  0.665 0.615 0.715 0.685 ;
        RECT  0.595 0.615 0.665 1.065 ;
        RECT  0.260 0.335 0.330 0.960 ;
        RECT  0.125 0.335 0.260 0.405 ;
        RECT  0.125 0.890 0.260 0.960 ;
        RECT  0.055 0.260 0.125 0.405 ;
        RECT  0.055 0.890 0.125 1.040 ;
    END
END FCICIND1BWP

MACRO FCICIND2BWP
    CLASS CORE ;
    FOREIGN FCICIND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.510 0.725 1.560 0.795 ;
        RECT  1.510 0.185 1.525 0.465 ;
        RECT  1.430 0.185 1.510 0.795 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.775 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.475 0.875 0.640 ;
        RECT  0.525 0.475 0.805 0.545 ;
        RECT  0.455 0.475 0.525 0.765 ;
        RECT  0.400 0.550 0.455 0.650 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.115 1.960 0.115 ;
        RECT  1.640 -0.115 1.720 0.415 ;
        RECT  1.345 -0.115 1.640 0.115 ;
        RECT  1.275 -0.115 1.345 0.465 ;
        RECT  0.560 -0.115 1.275 0.115 ;
        RECT  0.440 -0.115 0.560 0.260 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.145 1.960 1.375 ;
        RECT  1.620 1.010 1.740 1.375 ;
        RECT  0.525 1.145 1.620 1.375 ;
        RECT  0.455 0.870 0.525 1.375 ;
        RECT  0.000 1.145 0.455 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.855 0.240 1.925 1.020 ;
        RECT  1.835 0.240 1.855 0.380 ;
        RECT  1.835 0.870 1.855 1.020 ;
        RECT  1.520 0.870 1.835 0.940 ;
        RECT  1.450 0.870 1.520 1.065 ;
        RECT  0.665 0.995 1.450 1.065 ;
        RECT  1.025 0.545 1.320 0.615 ;
        RECT  0.805 0.855 1.190 0.925 ;
        RECT  1.095 0.195 1.165 0.455 ;
        RECT  0.680 0.195 1.095 0.265 ;
        RECT  0.955 0.335 1.025 0.785 ;
        RECT  0.330 0.335 0.955 0.405 ;
        RECT  0.890 0.715 0.955 0.785 ;
        RECT  0.735 0.785 0.805 0.925 ;
        RECT  0.665 0.615 0.715 0.685 ;
        RECT  0.595 0.615 0.665 1.065 ;
        RECT  0.260 0.335 0.330 0.960 ;
        RECT  0.125 0.335 0.260 0.405 ;
        RECT  0.125 0.890 0.260 0.960 ;
        RECT  0.055 0.260 0.125 0.405 ;
        RECT  0.055 0.890 0.125 1.040 ;
    END
END FCICIND2BWP

MACRO FCICOND1BWP
    CLASS CORE ;
    FOREIGN FCICOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CON
        ANTENNADIFFAREA 0.1585 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.070 0.490 1.085 0.800 ;
        RECT  1.025 0.335 1.070 0.800 ;
        RECT  1.000 0.335 1.025 0.895 ;
        RECT  0.330 0.335 1.000 0.405 ;
        RECT  0.955 0.730 1.000 0.895 ;
        RECT  0.260 0.335 0.330 0.905 ;
        RECT  0.125 0.335 0.260 0.410 ;
        RECT  0.125 0.835 0.260 0.905 ;
        RECT  0.035 0.215 0.125 0.410 ;
        RECT  0.055 0.835 0.125 1.045 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.615 0.750 0.685 ;
        RECT  0.595 0.615 0.665 0.905 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0424 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.475 0.920 0.660 ;
        RECT  0.525 0.475 0.845 0.545 ;
        RECT  0.455 0.475 0.525 0.765 ;
        RECT  0.415 0.560 0.455 0.680 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0528 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 -0.115 1.260 0.115 ;
        RECT  0.490 -0.115 0.610 0.265 ;
        RECT  0.000 -0.115 0.490 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 1.260 1.375 ;
        RECT  0.500 0.980 0.580 1.375 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.140 0.195 1.210 0.325 ;
        RECT  1.135 0.900 1.205 1.055 ;
        RECT  0.720 0.195 1.140 0.265 ;
        RECT  0.835 0.985 1.135 1.055 ;
        RECT  0.765 0.765 0.835 1.055 ;
    END
END FCICOND1BWP

MACRO FCICOND2BWP
    CLASS CORE ;
    FOREIGN FCICOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN CON
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.725 0.355 1.785 0.805 ;
        RECT  1.715 0.185 1.725 1.035 ;
        RECT  1.655 0.185 1.715 0.465 ;
        RECT  1.655 0.735 1.715 1.035 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.615 0.715 0.685 ;
        RECT  0.595 0.615 0.665 0.905 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.475 0.885 0.660 ;
        RECT  0.525 0.475 0.815 0.545 ;
        RECT  0.455 0.475 0.525 0.765 ;
        RECT  0.405 0.560 0.455 0.680 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0544 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.830 -0.115 1.910 0.300 ;
        RECT  1.550 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.550 0.305 ;
        RECT  0.550 -0.115 1.470 0.115 ;
        RECT  0.430 -0.115 0.550 0.260 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.905 1.145 1.960 1.375 ;
        RECT  1.835 0.905 1.905 1.375 ;
        RECT  1.550 1.145 1.835 1.375 ;
        RECT  1.470 0.860 1.550 1.375 ;
        RECT  0.580 1.145 1.470 1.375 ;
        RECT  0.500 0.985 0.580 1.375 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.585 0.520 1.610 0.640 ;
        RECT  1.515 0.385 1.585 0.790 ;
        RECT  1.365 0.385 1.515 0.455 ;
        RECT  1.365 0.720 1.515 0.790 ;
        RECT  1.345 0.530 1.445 0.630 ;
        RECT  1.295 0.195 1.365 0.455 ;
        RECT  1.295 0.720 1.365 1.035 ;
        RECT  1.035 0.530 1.345 0.600 ;
        RECT  1.115 0.195 1.185 0.455 ;
        RECT  1.115 0.765 1.185 1.055 ;
        RECT  0.680 0.195 1.115 0.265 ;
        RECT  0.805 0.985 1.115 1.055 ;
        RECT  0.965 0.335 1.035 0.895 ;
        RECT  0.330 0.335 0.965 0.405 ;
        RECT  0.925 0.755 0.965 0.895 ;
        RECT  0.735 0.765 0.805 1.055 ;
        RECT  0.260 0.335 0.330 0.960 ;
        RECT  0.125 0.335 0.260 0.405 ;
        RECT  0.125 0.890 0.260 0.960 ;
        RECT  0.055 0.260 0.125 0.405 ;
        RECT  0.055 0.890 0.125 1.040 ;
    END
END FCICOND2BWP

MACRO FCSICIND1BWP
    CLASS CORE ;
    FOREIGN FCSICIND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.175 0.185 7.245 1.045 ;
        RECT  7.155 0.185 7.175 0.465 ;
        RECT  7.160 0.745 7.175 1.045 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.940 0.215 6.970 0.485 ;
        RECT  6.895 0.215 6.940 0.640 ;
        RECT  6.860 0.415 6.895 0.640 ;
        END
    END CS
    PIN CO1
        ANTENNADIFFAREA 0.0871 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.090 0.775 4.165 0.915 ;
        RECT  4.090 0.475 4.140 0.545 ;
        RECT  4.020 0.475 4.090 0.915 ;
        END
    END CO1
    PIN CO0
        ANTENNADIFFAREA 0.0769 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.905 0.475 3.950 0.565 ;
        RECT  3.815 0.475 3.905 0.915 ;
        END
    END CO0
    PIN CIN1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.495 5.730 0.640 ;
        END
    END CIN1
    PIN CIN0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.530 2.250 0.635 ;
        RECT  2.135 0.355 2.205 0.635 ;
        RECT  2.115 0.355 2.135 0.460 ;
        END
    END CIN0
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.040 -0.115 7.280 0.115 ;
        RECT  6.920 -0.115 7.040 0.145 ;
        RECT  5.840 -0.115 6.920 0.115 ;
        RECT  5.720 -0.115 5.840 0.130 ;
        RECT  4.400 -0.115 5.720 0.115 ;
        RECT  4.280 -0.115 4.400 0.125 ;
        RECT  3.720 -0.115 4.280 0.115 ;
        RECT  3.600 -0.115 3.720 0.125 ;
        RECT  2.200 -0.115 3.600 0.115 ;
        RECT  2.075 -0.115 2.200 0.140 ;
        RECT  1.830 -0.115 2.075 0.115 ;
        RECT  1.705 -0.115 1.830 0.140 ;
        RECT  0.870 -0.115 1.705 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.270 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.060 1.145 7.280 1.375 ;
        RECT  6.940 1.010 7.060 1.375 ;
        RECT  5.880 1.145 6.940 1.375 ;
        RECT  5.760 1.130 5.880 1.375 ;
        RECT  4.320 1.145 5.760 1.375 ;
        RECT  4.200 1.135 4.320 1.375 ;
        RECT  3.720 1.145 4.200 1.375 ;
        RECT  3.600 1.135 3.720 1.375 ;
        RECT  2.180 1.145 3.600 1.375 ;
        RECT  2.060 1.130 2.180 1.375 ;
        RECT  1.810 1.145 2.060 1.375 ;
        RECT  1.690 1.130 1.810 1.375 ;
        RECT  0.890 1.145 1.690 1.375 ;
        RECT  0.765 1.125 0.890 1.375 ;
        RECT  0.510 1.145 0.765 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.090 0.540 7.105 0.660 ;
        RECT  7.020 0.540 7.090 0.940 ;
        RECT  6.840 0.870 7.020 0.940 ;
        RECT  6.790 0.720 6.870 0.790 ;
        RECT  6.770 0.870 6.840 1.065 ;
        RECT  6.790 0.230 6.815 0.350 ;
        RECT  6.720 0.230 6.790 0.790 ;
        RECT  6.445 0.995 6.770 1.065 ;
        RECT  6.670 0.520 6.720 0.640 ;
        RECT  6.600 0.845 6.650 0.915 ;
        RECT  6.600 0.325 6.620 0.445 ;
        RECT  6.530 0.195 6.600 0.915 ;
        RECT  6.030 0.195 6.530 0.265 ;
        RECT  6.375 0.355 6.445 1.065 ;
        RECT  6.355 0.805 6.375 1.065 ;
        RECT  6.175 0.335 6.245 1.060 ;
        RECT  6.150 0.335 6.175 0.460 ;
        RECT  5.210 0.990 6.175 1.060 ;
        RECT  6.010 0.340 6.080 0.920 ;
        RECT  5.960 0.195 6.030 0.270 ;
        RECT  5.940 0.340 6.010 0.460 ;
        RECT  5.105 0.850 6.010 0.920 ;
        RECT  5.680 0.200 5.960 0.270 ;
        RECT  5.870 0.530 5.940 0.630 ;
        RECT  5.800 0.345 5.870 0.780 ;
        RECT  5.530 0.345 5.800 0.415 ;
        RECT  5.390 0.710 5.800 0.780 ;
        RECT  5.610 0.195 5.680 0.270 ;
        RECT  2.640 0.195 5.610 0.265 ;
        RECT  5.355 0.335 5.425 0.565 ;
        RECT  5.310 0.495 5.355 0.565 ;
        RECT  5.240 0.495 5.310 0.780 ;
        RECT  5.170 0.345 5.260 0.415 ;
        RECT  5.200 0.680 5.240 0.780 ;
        RECT  5.105 0.345 5.170 0.605 ;
        RECT  5.100 0.345 5.105 0.960 ;
        RECT  5.035 0.535 5.100 0.960 ;
        RECT  4.960 0.345 5.025 0.465 ;
        RECT  4.890 0.345 4.960 0.920 ;
        RECT  4.340 0.850 4.890 0.920 ;
        RECT  4.750 0.345 4.820 0.780 ;
        RECT  4.620 0.690 4.750 0.780 ;
        RECT  1.585 0.990 4.750 1.060 ;
        RECT  4.605 0.540 4.680 0.610 ;
        RECT  4.550 0.345 4.605 0.610 ;
        RECT  4.535 0.345 4.550 0.780 ;
        RECT  4.480 0.540 4.535 0.780 ;
        RECT  4.420 0.690 4.480 0.780 ;
        RECT  4.320 0.335 4.410 0.550 ;
        RECT  4.270 0.625 4.340 0.920 ;
        RECT  3.625 0.335 4.320 0.405 ;
        RECT  4.160 0.625 4.270 0.695 ;
        RECT  3.675 0.615 3.745 0.920 ;
        RECT  3.045 0.850 3.675 0.920 ;
        RECT  3.555 0.335 3.625 0.550 ;
        RECT  3.455 0.710 3.500 0.780 ;
        RECT  3.380 0.345 3.455 0.780 ;
        RECT  3.300 0.545 3.380 0.615 ;
        RECT  3.225 0.710 3.300 0.780 ;
        RECT  3.155 0.345 3.225 0.780 ;
        RECT  2.975 0.345 3.045 0.920 ;
        RECT  2.835 0.370 2.905 0.920 ;
        RECT  2.710 0.370 2.835 0.440 ;
        RECT  1.825 0.850 2.835 0.920 ;
        RECT  2.655 0.545 2.725 0.770 ;
        RECT  2.640 0.545 2.655 0.615 ;
        RECT  2.570 0.195 2.640 0.615 ;
        RECT  2.470 0.370 2.570 0.440 ;
        RECT  2.400 0.710 2.570 0.780 ;
        RECT  2.380 0.185 2.500 0.280 ;
        RECT  2.330 0.355 2.400 0.780 ;
        RECT  1.225 0.210 2.380 0.280 ;
        RECT  2.280 0.355 2.330 0.455 ;
        RECT  2.065 0.710 2.330 0.780 ;
        RECT  1.965 0.530 2.065 0.780 ;
        RECT  1.825 0.375 2.010 0.445 ;
        RECT  1.755 0.375 1.825 0.920 ;
        RECT  1.585 0.350 1.605 0.590 ;
        RECT  1.535 0.350 1.585 1.060 ;
        RECT  1.515 0.520 1.535 1.060 ;
        RECT  1.435 0.520 1.515 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.210 1.225 0.905 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FCSICIND1BWP

MACRO FCSICIND2BWP
    CLASS CORE ;
    FOREIGN FCSICIND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0994 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.595 0.355 7.665 0.815 ;
        RECT  7.450 0.355 7.595 0.435 ;
        RECT  7.470 0.735 7.595 0.815 ;
        RECT  7.400 0.735 7.470 1.035 ;
        RECT  7.370 0.185 7.450 0.465 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0484 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.180 0.215 7.250 0.485 ;
        RECT  7.175 0.215 7.180 0.640 ;
        RECT  7.100 0.415 7.175 0.640 ;
        END
    END CS
    PIN CO1
        ANTENNADIFFAREA 0.0992 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.475 4.400 0.545 ;
        RECT  4.305 0.825 4.370 0.905 ;
        RECT  4.235 0.475 4.305 0.905 ;
        END
    END CO1
    PIN CO0
        ANTENNADIFFAREA 0.1118 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.475 4.025 0.905 ;
        RECT  3.810 0.475 3.955 0.545 ;
        RECT  3.830 0.825 3.955 0.905 ;
        END
    END CO0
    PIN CIN1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.495 5.990 0.640 ;
        END
    END CIN1
    PIN CIN0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.530 2.250 0.635 ;
        RECT  2.135 0.355 2.205 0.635 ;
        RECT  2.115 0.355 2.135 0.430 ;
        END
    END CIN0
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.640 -0.115 7.700 0.115 ;
        RECT  7.540 -0.115 7.640 0.270 ;
        RECT  7.280 -0.115 7.540 0.115 ;
        RECT  7.160 -0.115 7.280 0.135 ;
        RECT  6.100 -0.115 7.160 0.115 ;
        RECT  5.980 -0.115 6.100 0.130 ;
        RECT  4.620 -0.115 5.980 0.115 ;
        RECT  4.500 -0.115 4.620 0.125 ;
        RECT  4.180 -0.115 4.500 0.115 ;
        RECT  4.060 -0.115 4.180 0.125 ;
        RECT  3.700 -0.115 4.060 0.115 ;
        RECT  3.580 -0.115 3.700 0.125 ;
        RECT  2.200 -0.115 3.580 0.115 ;
        RECT  2.075 -0.115 2.200 0.140 ;
        RECT  1.830 -0.115 2.075 0.115 ;
        RECT  1.705 -0.115 1.830 0.140 ;
        RECT  0.870 -0.115 1.705 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.270 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.035 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.645 1.145 7.700 1.375 ;
        RECT  7.575 0.905 7.645 1.375 ;
        RECT  7.280 1.145 7.575 1.375 ;
        RECT  7.200 1.010 7.280 1.375 ;
        RECT  6.160 1.145 7.200 1.375 ;
        RECT  6.040 1.135 6.160 1.375 ;
        RECT  4.580 1.145 6.040 1.375 ;
        RECT  4.460 1.135 4.580 1.375 ;
        RECT  4.160 1.145 4.460 1.375 ;
        RECT  4.040 1.135 4.160 1.375 ;
        RECT  3.740 1.145 4.040 1.375 ;
        RECT  3.620 1.135 3.740 1.375 ;
        RECT  2.180 1.145 3.620 1.375 ;
        RECT  2.060 1.130 2.180 1.375 ;
        RECT  1.810 1.145 2.060 1.375 ;
        RECT  1.690 1.130 1.810 1.375 ;
        RECT  0.890 1.145 1.690 1.375 ;
        RECT  0.765 1.125 0.890 1.375 ;
        RECT  0.510 1.145 0.765 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.330 0.555 7.495 0.625 ;
        RECT  7.260 0.555 7.330 0.940 ;
        RECT  7.105 0.870 7.260 0.940 ;
        RECT  7.020 0.710 7.110 0.780 ;
        RECT  7.035 0.870 7.105 1.065 ;
        RECT  7.020 0.230 7.060 0.350 ;
        RECT  6.700 0.995 7.035 1.065 ;
        RECT  6.950 0.230 7.020 0.780 ;
        RECT  6.920 0.520 6.950 0.640 ;
        RECT  6.840 0.855 6.930 0.925 ;
        RECT  6.840 0.325 6.880 0.445 ;
        RECT  6.770 0.200 6.840 0.925 ;
        RECT  5.940 0.200 6.770 0.270 ;
        RECT  6.630 0.360 6.700 1.065 ;
        RECT  6.475 0.345 6.545 1.065 ;
        RECT  6.410 0.345 6.475 0.470 ;
        RECT  5.470 0.995 6.475 1.065 ;
        RECT  6.270 0.340 6.340 0.925 ;
        RECT  6.200 0.340 6.270 0.460 ;
        RECT  5.350 0.855 6.270 0.925 ;
        RECT  6.130 0.530 6.200 0.630 ;
        RECT  6.060 0.345 6.130 0.785 ;
        RECT  5.790 0.345 6.060 0.415 ;
        RECT  5.650 0.715 6.060 0.785 ;
        RECT  5.870 0.195 5.940 0.270 ;
        RECT  2.640 0.195 5.870 0.265 ;
        RECT  5.615 0.345 5.685 0.625 ;
        RECT  5.570 0.555 5.615 0.625 ;
        RECT  5.500 0.555 5.570 0.785 ;
        RECT  5.430 0.345 5.510 0.415 ;
        RECT  5.450 0.715 5.500 0.785 ;
        RECT  5.360 0.345 5.430 0.545 ;
        RECT  5.350 0.475 5.360 0.545 ;
        RECT  5.280 0.475 5.350 0.965 ;
        RECT  5.190 0.335 5.280 0.405 ;
        RECT  5.120 0.335 5.190 0.925 ;
        RECT  4.510 0.855 5.120 0.925 ;
        RECT  4.980 0.345 5.050 0.785 ;
        RECT  2.925 0.995 5.010 1.065 ;
        RECT  4.880 0.695 4.980 0.785 ;
        RECT  4.845 0.545 4.910 0.615 ;
        RECT  4.810 0.345 4.845 0.615 ;
        RECT  4.775 0.345 4.810 0.785 ;
        RECT  4.740 0.545 4.775 0.785 ;
        RECT  4.680 0.715 4.740 0.785 ;
        RECT  4.595 0.335 4.670 0.635 ;
        RECT  3.620 0.335 4.595 0.405 ;
        RECT  4.440 0.645 4.510 0.925 ;
        RECT  4.375 0.645 4.440 0.715 ;
        RECT  3.760 0.645 3.880 0.715 ;
        RECT  3.690 0.645 3.760 0.925 ;
        RECT  3.070 0.855 3.690 0.925 ;
        RECT  3.550 0.335 3.620 0.640 ;
        RECT  3.470 0.715 3.520 0.785 ;
        RECT  3.400 0.345 3.470 0.785 ;
        RECT  3.390 0.345 3.400 0.615 ;
        RECT  3.285 0.545 3.390 0.615 ;
        RECT  3.215 0.695 3.320 0.785 ;
        RECT  3.215 0.345 3.280 0.425 ;
        RECT  3.145 0.345 3.215 0.785 ;
        RECT  3.000 0.355 3.070 0.925 ;
        RECT  2.855 0.370 2.925 0.920 ;
        RECT  2.855 0.990 2.925 1.065 ;
        RECT  2.730 0.370 2.855 0.440 ;
        RECT  1.825 0.850 2.855 0.920 ;
        RECT  1.585 0.990 2.855 1.060 ;
        RECT  2.665 0.545 2.735 0.770 ;
        RECT  2.640 0.545 2.665 0.615 ;
        RECT  2.570 0.195 2.640 0.615 ;
        RECT  2.490 0.355 2.570 0.425 ;
        RECT  2.400 0.710 2.570 0.780 ;
        RECT  2.380 0.185 2.500 0.280 ;
        RECT  2.330 0.355 2.400 0.780 ;
        RECT  1.225 0.210 2.380 0.280 ;
        RECT  2.280 0.355 2.330 0.455 ;
        RECT  2.065 0.710 2.330 0.780 ;
        RECT  1.995 0.530 2.065 0.780 ;
        RECT  1.825 0.375 2.010 0.445 ;
        RECT  1.965 0.530 1.995 0.630 ;
        RECT  1.755 0.375 1.825 0.920 ;
        RECT  1.585 0.350 1.605 0.590 ;
        RECT  1.535 0.350 1.585 1.060 ;
        RECT  1.515 0.520 1.535 1.060 ;
        RECT  1.435 0.520 1.515 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.210 1.225 0.905 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FCSICIND2BWP

MACRO FCSICOND1BWP
    CLASS CORE ;
    FOREIGN FCSICOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.875 0.185 7.945 1.045 ;
        RECT  7.855 0.185 7.875 0.465 ;
        RECT  7.855 0.745 7.875 1.045 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.615 0.215 7.670 0.485 ;
        RECT  7.595 0.215 7.615 0.640 ;
        RECT  7.545 0.415 7.595 0.640 ;
        END
    END CS
    PIN CON1
        ANTENNADIFFAREA 0.0900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.485 4.540 0.555 ;
        RECT  4.445 0.840 4.530 0.910 ;
        RECT  4.375 0.485 4.445 0.910 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.0900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.485 4.165 0.910 ;
        RECT  4.020 0.485 4.095 0.555 ;
        RECT  4.030 0.840 4.095 0.910 ;
        END
    END CON0
    PIN CI1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.585 0.495 6.685 0.765 ;
        END
    END CI1
    PIN CI0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.495 1.935 0.765 ;
        END
    END CI0
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.740 -0.115 7.980 0.115 ;
        RECT  7.620 -0.115 7.740 0.135 ;
        RECT  6.480 -0.115 7.620 0.115 ;
        RECT  6.360 -0.115 6.480 0.135 ;
        RECT  4.960 -0.115 6.360 0.115 ;
        RECT  4.840 -0.115 4.960 0.135 ;
        RECT  4.340 -0.115 4.840 0.115 ;
        RECT  4.220 -0.115 4.340 0.135 ;
        RECT  3.720 -0.115 4.220 0.115 ;
        RECT  3.600 -0.115 3.720 0.135 ;
        RECT  2.200 -0.115 3.600 0.115 ;
        RECT  2.075 -0.115 2.200 0.140 ;
        RECT  1.830 -0.115 2.075 0.115 ;
        RECT  1.705 -0.115 1.830 0.140 ;
        RECT  0.870 -0.115 1.705 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.270 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.145 7.980 1.375 ;
        RECT  7.620 1.020 7.740 1.375 ;
        RECT  6.540 1.145 7.620 1.375 ;
        RECT  6.420 1.130 6.540 1.375 ;
        RECT  4.960 1.145 6.420 1.375 ;
        RECT  4.840 1.130 4.960 1.375 ;
        RECT  4.340 1.145 4.840 1.375 ;
        RECT  4.220 1.130 4.340 1.375 ;
        RECT  3.720 1.145 4.220 1.375 ;
        RECT  3.600 1.130 3.720 1.375 ;
        RECT  2.180 1.145 3.600 1.375 ;
        RECT  2.060 1.130 2.180 1.375 ;
        RECT  1.810 1.145 2.060 1.375 ;
        RECT  1.690 1.130 1.810 1.375 ;
        RECT  0.895 1.145 1.690 1.375 ;
        RECT  0.770 1.125 0.895 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.765 0.520 7.805 0.665 ;
        RECT  7.735 0.520 7.765 0.950 ;
        RECT  7.695 0.595 7.735 0.950 ;
        RECT  7.520 0.880 7.695 0.950 ;
        RECT  7.460 0.730 7.530 0.800 ;
        RECT  7.450 0.880 7.520 1.050 ;
        RECT  7.460 0.230 7.505 0.350 ;
        RECT  7.390 0.230 7.460 0.800 ;
        RECT  7.085 0.980 7.450 1.050 ;
        RECT  7.305 0.520 7.390 0.640 ;
        RECT  7.235 0.840 7.310 0.910 ;
        RECT  7.235 0.350 7.290 0.420 ;
        RECT  7.165 0.205 7.235 0.910 ;
        RECT  2.640 0.205 7.165 0.275 ;
        RECT  7.015 0.355 7.085 1.050 ;
        RECT  6.835 0.345 6.905 1.060 ;
        RECT  6.760 0.345 6.835 0.415 ;
        RECT  5.850 0.990 6.835 1.060 ;
        RECT  6.515 0.850 6.740 0.920 ;
        RECT  6.515 0.350 6.680 0.420 ;
        RECT  6.445 0.350 6.515 0.920 ;
        RECT  6.290 0.545 6.445 0.615 ;
        RECT  5.735 0.850 6.445 0.920 ;
        RECT  6.030 0.690 6.350 0.780 ;
        RECT  6.005 0.345 6.075 0.610 ;
        RECT  5.950 0.540 6.005 0.610 ;
        RECT  5.850 0.540 5.950 0.780 ;
        RECT  5.735 0.370 5.890 0.440 ;
        RECT  5.665 0.370 5.735 0.970 ;
        RECT  5.515 0.355 5.585 0.920 ;
        RECT  4.890 0.850 5.515 0.920 ;
        RECT  5.335 0.345 5.405 0.780 ;
        RECT  1.585 0.990 5.390 1.060 ;
        RECT  5.260 0.710 5.335 0.780 ;
        RECT  5.180 0.545 5.260 0.615 ;
        RECT  5.105 0.360 5.180 0.780 ;
        RECT  5.060 0.710 5.105 0.780 ;
        RECT  4.965 0.345 5.035 0.640 ;
        RECT  3.595 0.345 4.965 0.415 ;
        RECT  4.860 0.690 4.890 0.920 ;
        RECT  4.820 0.610 4.860 0.920 ;
        RECT  4.790 0.610 4.820 0.760 ;
        RECT  4.690 0.840 4.750 0.910 ;
        RECT  4.690 0.485 4.745 0.555 ;
        RECT  4.620 0.485 4.690 0.910 ;
        RECT  4.550 0.635 4.620 0.705 ;
        RECT  3.940 0.635 4.010 0.705 ;
        RECT  3.870 0.485 3.940 0.910 ;
        RECT  3.820 0.485 3.870 0.555 ;
        RECT  3.810 0.840 3.870 0.910 ;
        RECT  3.740 0.610 3.770 0.760 ;
        RECT  3.700 0.610 3.740 0.920 ;
        RECT  3.670 0.690 3.700 0.920 ;
        RECT  3.045 0.850 3.670 0.920 ;
        RECT  3.525 0.345 3.595 0.640 ;
        RECT  3.455 0.710 3.500 0.780 ;
        RECT  3.380 0.370 3.455 0.780 ;
        RECT  3.300 0.545 3.380 0.615 ;
        RECT  3.225 0.710 3.300 0.780 ;
        RECT  3.155 0.345 3.225 0.780 ;
        RECT  2.975 0.355 3.045 0.920 ;
        RECT  2.835 0.370 2.905 0.920 ;
        RECT  2.710 0.370 2.835 0.440 ;
        RECT  2.170 0.850 2.835 0.920 ;
        RECT  2.640 0.540 2.705 0.770 ;
        RECT  2.635 0.205 2.640 0.770 ;
        RECT  2.570 0.205 2.635 0.610 ;
        RECT  2.490 0.350 2.570 0.470 ;
        RECT  2.410 0.710 2.550 0.780 ;
        RECT  2.380 0.185 2.500 0.280 ;
        RECT  2.340 0.380 2.410 0.780 ;
        RECT  1.225 0.210 2.380 0.280 ;
        RECT  2.270 0.380 2.340 0.450 ;
        RECT  2.250 0.710 2.340 0.780 ;
        RECT  2.170 0.545 2.270 0.615 ;
        RECT  2.100 0.350 2.170 0.920 ;
        RECT  1.880 0.350 2.100 0.420 ;
        RECT  1.860 0.850 2.100 0.920 ;
        RECT  1.585 0.350 1.605 0.590 ;
        RECT  1.535 0.350 1.585 1.060 ;
        RECT  1.515 0.520 1.535 1.060 ;
        RECT  1.435 0.520 1.515 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.210 1.225 0.895 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FCSICOND1BWP

MACRO FCSICOND2BWP
    CLASS CORE ;
    FOREIGN FCSICOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.435 0.355 8.505 0.815 ;
        RECT  8.305 0.355 8.435 0.425 ;
        RECT  8.305 0.745 8.435 0.815 ;
        RECT  8.235 0.185 8.305 0.485 ;
        RECT  8.235 0.745 8.305 1.045 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.020 0.215 8.090 0.485 ;
        RECT  8.015 0.215 8.020 0.640 ;
        RECT  7.940 0.415 8.015 0.640 ;
        END
    END CS
    PIN CON1
        ANTENNADIFFAREA 0.1016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.585 0.485 4.740 0.555 ;
        RECT  4.585 0.775 4.725 0.905 ;
        RECT  4.515 0.485 4.585 0.905 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.1080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.485 4.445 0.905 ;
        RECT  4.210 0.485 4.375 0.555 ;
        RECT  4.235 0.775 4.375 0.905 ;
        END
    END CON0
    PIN CI1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.035 0.495 7.105 0.765 ;
        RECT  6.965 0.495 7.035 0.640 ;
        END
    END CI1
    PIN CI0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.495 1.935 0.765 ;
        END
    END CI0
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.500 -0.115 8.540 0.115 ;
        RECT  8.400 -0.115 8.500 0.270 ;
        RECT  8.120 -0.115 8.400 0.115 ;
        RECT  8.000 -0.115 8.120 0.135 ;
        RECT  6.865 -0.115 8.000 0.115 ;
        RECT  6.740 -0.115 6.865 0.135 ;
        RECT  5.340 -0.115 6.740 0.115 ;
        RECT  5.220 -0.115 5.340 0.135 ;
        RECT  4.940 -0.115 5.220 0.115 ;
        RECT  4.815 -0.115 4.940 0.135 ;
        RECT  4.540 -0.115 4.815 0.115 ;
        RECT  4.415 -0.115 4.540 0.135 ;
        RECT  4.130 -0.115 4.415 0.115 ;
        RECT  4.005 -0.115 4.130 0.135 ;
        RECT  3.720 -0.115 4.005 0.115 ;
        RECT  3.600 -0.115 3.720 0.135 ;
        RECT  2.200 -0.115 3.600 0.115 ;
        RECT  2.075 -0.115 2.200 0.140 ;
        RECT  1.830 -0.115 2.075 0.115 ;
        RECT  1.705 -0.115 1.830 0.140 ;
        RECT  0.870 -0.115 1.705 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.270 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.490 1.145 8.540 1.375 ;
        RECT  8.410 0.915 8.490 1.375 ;
        RECT  8.120 1.145 8.410 1.375 ;
        RECT  8.000 1.020 8.120 1.375 ;
        RECT  6.920 1.145 8.000 1.375 ;
        RECT  6.800 1.130 6.920 1.375 ;
        RECT  5.340 1.145 6.800 1.375 ;
        RECT  5.220 1.130 5.340 1.375 ;
        RECT  4.930 1.145 5.220 1.375 ;
        RECT  4.810 1.130 4.930 1.375 ;
        RECT  4.540 1.145 4.810 1.375 ;
        RECT  4.420 1.130 4.540 1.375 ;
        RECT  4.130 1.145 4.420 1.375 ;
        RECT  4.005 1.130 4.130 1.375 ;
        RECT  3.720 1.145 4.005 1.375 ;
        RECT  3.600 1.130 3.720 1.375 ;
        RECT  2.180 1.145 3.600 1.375 ;
        RECT  2.060 1.130 2.180 1.375 ;
        RECT  1.810 1.145 2.060 1.375 ;
        RECT  1.690 1.130 1.810 1.375 ;
        RECT  0.895 1.145 1.690 1.375 ;
        RECT  0.770 1.125 0.895 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.165 0.555 8.325 0.625 ;
        RECT  8.095 0.555 8.165 0.950 ;
        RECT  7.900 0.880 8.095 0.950 ;
        RECT  7.860 0.255 7.910 0.325 ;
        RECT  7.860 0.730 7.910 0.800 ;
        RECT  7.830 0.880 7.900 1.050 ;
        RECT  7.790 0.255 7.860 0.800 ;
        RECT  7.465 0.980 7.830 1.050 ;
        RECT  7.685 0.520 7.790 0.640 ;
        RECT  7.615 0.840 7.690 0.910 ;
        RECT  7.615 0.350 7.670 0.420 ;
        RECT  7.545 0.205 7.615 0.910 ;
        RECT  2.640 0.205 7.545 0.275 ;
        RECT  7.395 0.355 7.465 1.050 ;
        RECT  7.215 0.345 7.285 1.060 ;
        RECT  7.140 0.345 7.215 0.415 ;
        RECT  6.230 0.990 7.215 1.060 ;
        RECT  6.895 0.850 7.120 0.920 ;
        RECT  6.895 0.350 7.060 0.420 ;
        RECT  6.825 0.350 6.895 0.920 ;
        RECT  6.670 0.545 6.825 0.615 ;
        RECT  6.115 0.850 6.825 0.920 ;
        RECT  6.410 0.690 6.730 0.780 ;
        RECT  6.385 0.345 6.455 0.610 ;
        RECT  6.330 0.540 6.385 0.610 ;
        RECT  6.230 0.540 6.330 0.780 ;
        RECT  6.115 0.370 6.270 0.440 ;
        RECT  6.045 0.370 6.115 0.960 ;
        RECT  5.895 0.355 5.965 0.920 ;
        RECT  5.270 0.850 5.895 0.920 ;
        RECT  5.715 0.345 5.785 0.780 ;
        RECT  1.585 0.990 5.770 1.060 ;
        RECT  5.640 0.710 5.715 0.780 ;
        RECT  5.560 0.545 5.640 0.615 ;
        RECT  5.485 0.360 5.560 0.780 ;
        RECT  5.440 0.710 5.485 0.780 ;
        RECT  5.345 0.345 5.415 0.640 ;
        RECT  3.595 0.345 5.345 0.415 ;
        RECT  5.200 0.635 5.270 0.920 ;
        RECT  5.120 0.635 5.200 0.705 ;
        RECT  4.890 0.840 5.130 0.910 ;
        RECT  4.890 0.485 5.115 0.555 ;
        RECT  4.820 0.485 4.890 0.910 ;
        RECT  4.055 0.485 4.125 0.910 ;
        RECT  3.825 0.485 4.055 0.555 ;
        RECT  3.810 0.840 4.055 0.910 ;
        RECT  3.740 0.635 3.820 0.705 ;
        RECT  3.670 0.635 3.740 0.920 ;
        RECT  3.045 0.850 3.670 0.920 ;
        RECT  3.525 0.345 3.595 0.640 ;
        RECT  3.455 0.710 3.500 0.780 ;
        RECT  3.380 0.370 3.455 0.780 ;
        RECT  3.300 0.545 3.380 0.615 ;
        RECT  3.225 0.710 3.300 0.780 ;
        RECT  3.155 0.345 3.225 0.780 ;
        RECT  2.975 0.355 3.045 0.920 ;
        RECT  2.835 0.370 2.905 0.920 ;
        RECT  2.710 0.370 2.835 0.440 ;
        RECT  2.170 0.850 2.835 0.920 ;
        RECT  2.640 0.540 2.705 0.770 ;
        RECT  2.635 0.205 2.640 0.770 ;
        RECT  2.570 0.205 2.635 0.610 ;
        RECT  2.490 0.350 2.570 0.470 ;
        RECT  2.410 0.710 2.550 0.780 ;
        RECT  2.380 0.185 2.500 0.280 ;
        RECT  2.340 0.380 2.410 0.780 ;
        RECT  1.225 0.210 2.380 0.280 ;
        RECT  2.270 0.380 2.340 0.450 ;
        RECT  2.250 0.710 2.340 0.780 ;
        RECT  2.170 0.545 2.270 0.615 ;
        RECT  2.100 0.350 2.170 0.920 ;
        RECT  1.880 0.350 2.100 0.420 ;
        RECT  1.860 0.850 2.100 0.920 ;
        RECT  1.585 0.350 1.605 0.590 ;
        RECT  1.535 0.350 1.585 1.060 ;
        RECT  1.515 0.520 1.535 1.060 ;
        RECT  1.435 0.520 1.515 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.210 1.225 0.895 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FCSICOND2BWP

MACRO FICIND1BWP
    CLASS CORE ;
    FOREIGN FICIND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0868 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.700 3.650 0.770 ;
        RECT  3.530 0.185 3.625 0.770 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 3.075 0.640 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.740 -0.115 3.820 0.450 ;
        RECT  3.240 -0.115 3.740 0.115 ;
        RECT  3.120 -0.115 3.240 0.140 ;
        RECT  1.820 -0.115 3.120 0.115 ;
        RECT  1.700 -0.115 1.820 0.135 ;
        RECT  0.870 -0.115 1.700 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.270 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.145 4.060 1.375 ;
        RECT  3.720 1.005 3.840 1.375 ;
        RECT  3.200 1.145 3.720 1.375 ;
        RECT  3.080 1.130 3.200 1.375 ;
        RECT  1.810 1.145 3.080 1.375 ;
        RECT  1.690 1.010 1.810 1.375 ;
        RECT  0.895 1.145 1.690 1.375 ;
        RECT  0.770 1.125 0.895 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.855 0.520 3.880 0.640 ;
        RECT  3.785 0.520 3.855 0.920 ;
        RECT  2.765 0.850 3.785 0.920 ;
        RECT  2.345 0.990 3.540 1.060 ;
        RECT  3.360 0.210 3.430 0.780 ;
        RECT  2.625 0.210 3.360 0.280 ;
        RECT  3.290 0.690 3.360 0.780 ;
        RECT  3.220 0.540 3.290 0.610 ;
        RECT  3.150 0.350 3.220 0.780 ;
        RECT  2.910 0.350 3.150 0.420 ;
        RECT  2.860 0.710 3.150 0.780 ;
        RECT  2.765 0.350 2.830 0.420 ;
        RECT  2.695 0.350 2.765 0.920 ;
        RECT  2.620 0.850 2.695 0.920 ;
        RECT  2.555 0.210 2.625 0.575 ;
        RECT  2.525 0.505 2.555 0.575 ;
        RECT  2.455 0.505 2.525 0.910 ;
        RECT  2.345 0.355 2.450 0.425 ;
        RECT  2.275 0.355 2.345 1.060 ;
        RECT  2.160 0.335 2.205 0.920 ;
        RECT  2.135 0.335 2.160 1.075 ;
        RECT  2.060 0.850 2.135 1.075 ;
        RECT  1.995 0.385 2.065 0.780 ;
        RECT  1.605 0.850 2.060 0.920 ;
        RECT  1.985 0.385 1.995 0.455 ;
        RECT  1.870 0.710 1.995 0.780 ;
        RECT  1.915 0.195 1.985 0.455 ;
        RECT  1.805 0.545 1.900 0.615 ;
        RECT  1.735 0.205 1.805 0.615 ;
        RECT  1.225 0.205 1.735 0.275 ;
        RECT  1.535 0.345 1.605 1.035 ;
        RECT  1.530 0.345 1.535 0.640 ;
        RECT  1.465 0.520 1.530 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.205 1.225 0.905 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FICIND1BWP

MACRO FICIND2BWP
    CLASS CORE ;
    FOREIGN FICIND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 0.185 4.310 0.790 ;
        RECT  4.235 0.185 4.240 0.485 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.670 0.355 4.725 0.805 ;
        RECT  4.665 0.355 4.670 1.035 ;
        RECT  4.655 0.185 4.665 1.035 ;
        RECT  4.595 0.185 4.655 0.465 ;
        RECT  4.600 0.735 4.655 1.035 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.625 0.765 ;
        END
    END CIN
    PIN B
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.495 1.925 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.330 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.300 ;
        RECT  4.485 -0.115 4.775 0.115 ;
        RECT  4.415 -0.115 4.485 0.420 ;
        RECT  4.115 -0.115 4.415 0.115 ;
        RECT  4.045 -0.115 4.115 0.305 ;
        RECT  3.760 -0.115 4.045 0.115 ;
        RECT  3.640 -0.115 3.760 0.135 ;
        RECT  3.370 -0.115 3.640 0.115 ;
        RECT  3.250 -0.115 3.370 0.135 ;
        RECT  2.040 -0.115 3.250 0.115 ;
        RECT  1.920 -0.115 2.040 0.140 ;
        RECT  0.880 -0.115 1.920 0.115 ;
        RECT  0.760 -0.115 0.880 0.140 ;
        RECT  0.490 -0.115 0.760 0.115 ;
        RECT  0.410 -0.115 0.490 0.275 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.895 4.845 1.375 ;
        RECT  4.510 1.145 4.775 1.375 ;
        RECT  4.390 1.010 4.510 1.375 ;
        RECT  4.120 1.145 4.390 1.375 ;
        RECT  4.000 1.135 4.120 1.375 ;
        RECT  3.700 1.145 4.000 1.375 ;
        RECT  3.580 1.135 3.700 1.375 ;
        RECT  1.990 1.145 3.580 1.375 ;
        RECT  1.870 1.025 1.990 1.375 ;
        RECT  0.880 1.145 1.870 1.375 ;
        RECT  0.760 1.120 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.530 0.520 4.550 0.640 ;
        RECT  4.460 0.520 4.530 0.940 ;
        RECT  4.310 0.870 4.460 0.940 ;
        RECT  4.240 0.870 4.310 1.065 ;
        RECT  2.570 0.995 4.240 1.065 ;
        RECT  4.095 0.515 4.170 0.925 ;
        RECT  2.920 0.855 4.095 0.925 ;
        RECT  3.955 0.390 4.025 0.785 ;
        RECT  3.925 0.390 3.955 0.470 ;
        RECT  3.790 0.715 3.955 0.785 ;
        RECT  3.855 0.205 3.925 0.470 ;
        RECT  3.775 0.545 3.860 0.615 ;
        RECT  2.780 0.205 3.855 0.275 ;
        RECT  3.705 0.355 3.775 0.615 ;
        RECT  3.140 0.355 3.705 0.425 ;
        RECT  3.395 0.655 3.465 0.785 ;
        RECT  3.140 0.715 3.395 0.785 ;
        RECT  3.070 0.355 3.140 0.785 ;
        RECT  3.010 0.715 3.070 0.785 ;
        RECT  2.920 0.360 3.000 0.460 ;
        RECT  2.850 0.360 2.920 0.925 ;
        RECT  2.790 0.855 2.850 0.925 ;
        RECT  2.710 0.205 2.780 0.630 ;
        RECT  2.640 0.560 2.710 0.910 ;
        RECT  2.570 0.345 2.620 0.415 ;
        RECT  2.500 0.345 2.570 1.065 ;
        RECT  2.430 0.995 2.500 1.065 ;
        RECT  2.365 0.320 2.430 0.810 ;
        RECT  2.360 0.320 2.365 0.955 ;
        RECT  2.335 0.320 2.360 0.440 ;
        RECT  2.295 0.740 2.360 0.955 ;
        RECT  1.760 0.885 2.295 0.955 ;
        RECT  2.225 0.520 2.290 0.640 ;
        RECT  2.155 0.195 2.225 0.815 ;
        RECT  2.050 0.745 2.155 0.815 ;
        RECT  2.015 0.210 2.085 0.640 ;
        RECT  1.405 0.210 2.015 0.280 ;
        RECT  1.760 0.350 1.830 0.420 ;
        RECT  1.690 0.350 1.760 1.055 ;
        RECT  1.630 0.540 1.690 0.640 ;
        RECT  1.555 0.350 1.620 0.470 ;
        RECT  1.565 0.790 1.585 0.910 ;
        RECT  1.555 0.790 1.565 1.050 ;
        RECT  1.485 0.350 1.555 1.050 ;
        RECT  0.665 0.980 1.485 1.050 ;
        RECT  1.335 0.210 1.405 0.910 ;
        RECT  0.860 0.840 1.250 0.910 ;
        RECT  1.155 0.210 1.225 0.370 ;
        RECT  1.070 0.545 1.180 0.615 ;
        RECT  0.860 0.210 1.155 0.280 ;
        RECT  0.995 0.355 1.070 0.760 ;
        RECT  0.950 0.355 0.995 0.425 ;
        RECT  0.950 0.690 0.995 0.760 ;
        RECT  0.790 0.210 0.860 0.910 ;
        RECT  0.570 0.345 0.790 0.415 ;
        RECT  0.570 0.730 0.790 0.800 ;
        RECT  0.595 0.870 0.665 1.050 ;
        RECT  0.485 0.545 0.650 0.615 ;
        RECT  0.485 0.870 0.595 0.940 ;
        RECT  0.415 0.345 0.485 0.940 ;
        RECT  0.330 0.345 0.415 0.415 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.205 0.330 0.415 ;
        RECT  0.235 0.750 0.305 1.045 ;
    END
END FICIND2BWP

MACRO FICOND1BWP
    CLASS CORE ;
    FOREIGN FICOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.185 4.305 1.070 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.925 0.405 3.995 0.780 ;
        RECT  3.920 0.405 3.925 0.485 ;
        RECT  3.830 0.710 3.925 0.780 ;
        RECT  3.815 0.205 3.920 0.485 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.355 3.340 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.960 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.105 -0.115 4.340 0.115 ;
        RECT  4.035 -0.115 4.105 0.315 ;
        RECT  3.745 -0.115 4.035 0.115 ;
        RECT  3.675 -0.115 3.745 0.465 ;
        RECT  3.220 -0.115 3.675 0.115 ;
        RECT  3.100 -0.115 3.220 0.140 ;
        RECT  1.840 -0.115 3.100 0.115 ;
        RECT  1.720 -0.115 1.840 0.125 ;
        RECT  0.870 -0.115 1.720 0.115 ;
        RECT  0.750 -0.115 0.870 0.260 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.260 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.145 4.340 1.375 ;
        RECT  4.010 1.010 4.130 1.375 ;
        RECT  3.770 1.145 4.010 1.375 ;
        RECT  3.650 1.005 3.770 1.375 ;
        RECT  3.180 1.145 3.650 1.375 ;
        RECT  3.060 1.130 3.180 1.375 ;
        RECT  1.800 1.145 3.060 1.375 ;
        RECT  1.680 1.010 1.800 1.375 ;
        RECT  0.890 1.145 1.680 1.375 ;
        RECT  0.765 1.125 0.890 1.375 ;
        RECT  0.510 1.145 0.765 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.075 0.510 4.145 0.920 ;
        RECT  2.760 0.850 4.075 0.920 ;
        RECT  3.590 0.555 3.840 0.625 ;
        RECT  3.565 0.555 3.590 0.780 ;
        RECT  3.495 0.185 3.565 0.780 ;
        RECT  3.470 0.710 3.495 0.780 ;
        RECT  2.350 0.990 3.480 1.060 ;
        RECT  3.170 0.210 3.410 0.280 ;
        RECT  3.170 0.710 3.370 0.780 ;
        RECT  3.100 0.210 3.170 0.780 ;
        RECT  2.620 0.210 3.100 0.280 ;
        RECT  3.030 0.520 3.100 0.640 ;
        RECT  2.960 0.360 3.030 0.430 ;
        RECT  2.960 0.700 2.990 0.770 ;
        RECT  2.890 0.360 2.960 0.770 ;
        RECT  2.870 0.700 2.890 0.770 ;
        RECT  2.760 0.350 2.820 0.450 ;
        RECT  2.690 0.350 2.760 0.920 ;
        RECT  2.620 0.850 2.690 0.920 ;
        RECT  2.550 0.210 2.620 0.725 ;
        RECT  2.525 0.655 2.550 0.725 ;
        RECT  2.455 0.655 2.525 0.900 ;
        RECT  2.350 0.350 2.415 0.550 ;
        RECT  2.040 0.195 2.350 0.275 ;
        RECT  2.345 0.350 2.350 1.060 ;
        RECT  2.280 0.480 2.345 1.060 ;
        RECT  2.130 0.355 2.200 0.940 ;
        RECT  1.600 0.870 2.130 0.940 ;
        RECT  1.960 0.195 2.040 0.800 ;
        RECT  1.870 0.730 1.960 0.800 ;
        RECT  1.850 0.520 1.890 0.640 ;
        RECT  1.780 0.205 1.850 0.640 ;
        RECT  1.225 0.205 1.780 0.275 ;
        RECT  1.530 0.345 1.600 1.035 ;
        RECT  1.515 0.520 1.530 1.035 ;
        RECT  1.435 0.520 1.515 0.640 ;
        RECT  1.365 0.355 1.450 0.425 ;
        RECT  1.365 0.775 1.405 0.895 ;
        RECT  1.295 0.355 1.365 1.055 ;
        RECT  0.650 0.985 1.295 1.055 ;
        RECT  1.150 0.205 1.225 0.905 ;
        RECT  1.135 0.205 1.150 0.325 ;
        RECT  0.800 0.845 1.070 0.915 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.800 0.340 0.940 0.425 ;
        RECT  0.730 0.340 0.800 0.915 ;
        RECT  0.680 0.340 0.730 0.425 ;
        RECT  0.570 0.730 0.730 0.800 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.580 0.870 0.650 1.055 ;
        RECT  0.485 0.545 0.640 0.615 ;
        RECT  0.485 0.870 0.580 0.940 ;
        RECT  0.415 0.340 0.485 0.940 ;
        RECT  0.330 0.340 0.415 0.410 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.210 0.200 0.330 0.410 ;
        RECT  0.235 0.735 0.305 1.035 ;
    END
END FICOND1BWP

MACRO FICOND2BWP
    CLASS CORE ;
    FOREIGN FICOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.670 0.355 4.725 0.805 ;
        RECT  4.665 0.355 4.670 1.035 ;
        RECT  4.655 0.185 4.665 1.035 ;
        RECT  4.595 0.185 4.655 0.465 ;
        RECT  4.595 0.735 4.655 1.035 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.370 0.215 4.445 0.345 ;
        RECT  4.300 0.215 4.370 0.785 ;
        RECT  4.215 0.215 4.300 0.475 ;
        RECT  4.190 0.715 4.300 0.785 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.625 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.0776 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.495 1.925 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.270 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.300 ;
        RECT  4.500 -0.115 4.775 0.115 ;
        RECT  4.380 -0.115 4.500 0.130 ;
        RECT  4.105 -0.115 4.380 0.115 ;
        RECT  4.035 -0.115 4.105 0.460 ;
        RECT  3.745 -0.115 4.035 0.115 ;
        RECT  3.675 -0.115 3.745 0.280 ;
        RECT  3.400 -0.115 3.675 0.115 ;
        RECT  3.280 -0.115 3.400 0.140 ;
        RECT  2.020 -0.115 3.280 0.115 ;
        RECT  1.900 -0.115 2.020 0.140 ;
        RECT  0.880 -0.115 1.900 0.115 ;
        RECT  0.760 -0.115 0.880 0.140 ;
        RECT  0.490 -0.115 0.760 0.115 ;
        RECT  0.410 -0.115 0.490 0.275 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.895 4.845 1.375 ;
        RECT  4.500 1.145 4.775 1.375 ;
        RECT  4.380 1.005 4.500 1.375 ;
        RECT  4.100 1.145 4.380 1.375 ;
        RECT  3.980 1.135 4.100 1.375 ;
        RECT  3.800 1.145 3.980 1.375 ;
        RECT  3.680 1.135 3.800 1.375 ;
        RECT  3.380 1.145 3.680 1.375 ;
        RECT  3.260 1.135 3.380 1.375 ;
        RECT  1.990 1.145 3.260 1.375 ;
        RECT  1.870 1.025 1.990 1.375 ;
        RECT  0.880 1.145 1.870 1.375 ;
        RECT  0.760 1.120 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.010 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.525 0.545 4.585 0.615 ;
        RECT  4.455 0.545 4.525 0.925 ;
        RECT  2.920 0.855 4.455 0.925 ;
        RECT  3.950 0.545 4.215 0.615 ;
        RECT  3.925 0.545 3.950 0.775 ;
        RECT  3.830 0.995 3.950 1.070 ;
        RECT  3.855 0.185 3.925 0.775 ;
        RECT  3.830 0.705 3.855 0.775 ;
        RECT  2.530 0.995 3.830 1.065 ;
        RECT  3.360 0.210 3.590 0.280 ;
        RECT  3.360 0.715 3.590 0.785 ;
        RECT  3.290 0.210 3.360 0.785 ;
        RECT  2.780 0.210 3.290 0.280 ;
        RECT  3.220 0.520 3.290 0.640 ;
        RECT  3.150 0.360 3.210 0.430 ;
        RECT  3.080 0.360 3.150 0.785 ;
        RECT  3.030 0.715 3.080 0.785 ;
        RECT  2.920 0.360 3.010 0.430 ;
        RECT  2.850 0.360 2.920 0.925 ;
        RECT  2.790 0.855 2.850 0.925 ;
        RECT  2.710 0.210 2.780 0.630 ;
        RECT  2.705 0.560 2.710 0.630 ;
        RECT  2.635 0.560 2.705 0.910 ;
        RECT  2.530 0.345 2.600 0.415 ;
        RECT  2.460 0.345 2.530 1.065 ;
        RECT  2.320 0.320 2.390 0.955 ;
        RECT  2.295 0.320 2.320 0.440 ;
        RECT  1.760 0.885 2.320 0.955 ;
        RECT  2.215 0.520 2.250 0.640 ;
        RECT  2.145 0.210 2.215 0.815 ;
        RECT  2.090 0.210 2.145 0.280 ;
        RECT  2.050 0.745 2.145 0.815 ;
        RECT  2.005 0.350 2.075 0.640 ;
        RECT  1.990 0.350 2.005 0.420 ;
        RECT  1.920 0.210 1.990 0.420 ;
        RECT  1.405 0.210 1.920 0.280 ;
        RECT  1.760 0.350 1.830 0.420 ;
        RECT  1.690 0.350 1.760 1.055 ;
        RECT  1.625 0.540 1.690 0.640 ;
        RECT  1.555 0.350 1.620 0.470 ;
        RECT  1.565 0.790 1.585 0.910 ;
        RECT  1.555 0.790 1.565 1.050 ;
        RECT  1.485 0.350 1.555 1.050 ;
        RECT  0.665 0.980 1.485 1.050 ;
        RECT  1.335 0.210 1.405 0.910 ;
        RECT  0.860 0.840 1.250 0.910 ;
        RECT  1.155 0.210 1.225 0.370 ;
        RECT  1.070 0.545 1.180 0.615 ;
        RECT  0.860 0.210 1.155 0.280 ;
        RECT  0.995 0.355 1.070 0.760 ;
        RECT  0.950 0.355 0.995 0.425 ;
        RECT  0.950 0.690 0.995 0.760 ;
        RECT  0.790 0.210 0.860 0.910 ;
        RECT  0.570 0.345 0.790 0.415 ;
        RECT  0.570 0.730 0.790 0.800 ;
        RECT  0.595 0.870 0.665 1.050 ;
        RECT  0.485 0.545 0.650 0.615 ;
        RECT  0.485 0.870 0.595 0.940 ;
        RECT  0.415 0.395 0.485 0.940 ;
        RECT  0.305 0.395 0.415 0.465 ;
        RECT  0.305 0.870 0.415 0.940 ;
        RECT  0.235 0.205 0.305 0.465 ;
        RECT  0.235 0.750 0.305 1.045 ;
    END
END FICOND2BWP

MACRO FIICOND1BWP
    CLASS CORE ;
    FOREIGN FIICOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.045 ;
        RECT  4.075 0.185 4.095 0.465 ;
        RECT  4.075 0.735 4.095 1.045 ;
        END
    END S
    PIN CON1
        ANTENNADIFFAREA 0.0947 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.730 0.945 0.800 ;
        RECT  0.670 0.355 0.750 0.425 ;
        RECT  0.595 0.355 0.670 0.800 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.0997 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.735 0.315 1.035 ;
        RECT  0.105 0.735 0.245 0.805 ;
        RECT  0.105 0.215 0.125 0.355 ;
        RECT  0.035 0.215 0.105 0.805 ;
        END
    END CON0
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.490 3.755 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1044 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.990 2.400 1.070 ;
        RECT  1.645 0.990 2.280 1.060 ;
        RECT  1.575 0.870 1.645 1.060 ;
        RECT  0.525 0.870 1.575 0.940 ;
        RECT  0.455 0.495 0.525 0.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1128 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.210 0.945 0.640 ;
        RECT  0.385 0.210 0.875 0.280 ;
        RECT  0.315 0.210 0.385 0.640 ;
        RECT  0.175 0.520 0.315 0.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 -0.115 4.200 0.115 ;
        RECT  3.860 -0.115 3.980 0.140 ;
        RECT  3.600 -0.115 3.860 0.115 ;
        RECT  3.480 -0.115 3.600 0.140 ;
        RECT  2.625 -0.115 3.480 0.115 ;
        RECT  2.555 -0.115 2.625 0.455 ;
        RECT  1.740 -0.115 2.555 0.115 ;
        RECT  1.620 -0.115 1.740 0.140 ;
        RECT  1.340 -0.115 1.620 0.115 ;
        RECT  1.220 -0.115 1.340 0.140 ;
        RECT  0.940 -0.115 1.220 0.115 ;
        RECT  0.820 -0.115 0.940 0.140 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.140 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.955 1.145 4.200 1.375 ;
        RECT  3.885 0.735 3.955 1.375 ;
        RECT  3.610 1.145 3.885 1.375 ;
        RECT  3.490 1.030 3.610 1.375 ;
        RECT  2.690 1.145 3.490 1.375 ;
        RECT  2.570 0.995 2.690 1.375 ;
        RECT  1.800 1.145 2.570 1.375 ;
        RECT  1.680 1.130 1.800 1.375 ;
        RECT  1.430 1.145 1.680 1.375 ;
        RECT  1.310 1.010 1.430 1.375 ;
        RECT  1.070 1.145 1.310 1.375 ;
        RECT  0.950 1.010 1.070 1.375 ;
        RECT  0.530 1.145 0.950 1.375 ;
        RECT  0.410 1.030 0.530 1.375 ;
        RECT  0.125 1.145 0.410 1.375 ;
        RECT  0.055 0.895 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.985 0.520 4.020 0.640 ;
        RECT  3.915 0.210 3.985 0.640 ;
        RECT  3.230 0.210 3.915 0.280 ;
        RECT  3.595 0.350 3.790 0.420 ;
        RECT  3.595 0.890 3.790 0.960 ;
        RECT  3.525 0.350 3.595 0.960 ;
        RECT  3.450 0.520 3.525 0.640 ;
        RECT  3.405 0.890 3.525 0.960 ;
        RECT  3.380 0.720 3.430 0.790 ;
        RECT  3.335 0.890 3.405 1.065 ;
        RECT  3.310 0.360 3.380 0.790 ;
        RECT  3.090 0.995 3.335 1.065 ;
        RECT  3.160 0.185 3.230 0.915 ;
        RECT  3.090 0.185 3.160 0.255 ;
        RECT  3.020 0.330 3.090 1.065 ;
        RECT  2.890 0.330 3.020 0.400 ;
        RECT  2.930 0.995 3.020 1.065 ;
        RECT  2.880 0.470 2.950 0.855 ;
        RECT  2.805 0.470 2.880 0.540 ;
        RECT  2.845 0.785 2.880 0.855 ;
        RECT  2.775 0.785 2.845 1.045 ;
        RECT  2.735 0.185 2.805 0.540 ;
        RECT  2.670 0.610 2.800 0.680 ;
        RECT  2.600 0.610 2.670 0.920 ;
        RECT  2.090 0.850 2.600 0.920 ;
        RECT  2.470 0.680 2.500 0.780 ;
        RECT  2.400 0.185 2.470 0.780 ;
        RECT  2.375 0.185 2.400 0.610 ;
        RECT  2.310 0.490 2.375 0.610 ;
        RECT  2.240 0.680 2.320 0.780 ;
        RECT  2.240 0.210 2.290 0.280 ;
        RECT  2.170 0.210 2.240 0.780 ;
        RECT  1.105 0.210 2.170 0.280 ;
        RECT  2.020 0.360 2.090 0.920 ;
        RECT  1.970 0.360 2.020 0.430 ;
        RECT  1.885 0.730 1.945 0.900 ;
        RECT  1.875 0.350 1.885 0.900 ;
        RECT  1.815 0.350 1.875 0.800 ;
        RECT  1.420 0.350 1.815 0.420 ;
        RECT  1.490 0.730 1.815 0.800 ;
        RECT  1.110 0.545 1.580 0.615 ;
        RECT  1.110 0.730 1.260 0.800 ;
        RECT  1.105 0.545 1.110 0.800 ;
        RECT  1.035 0.210 1.105 0.800 ;
    END
END FIICOND1BWP

MACRO FIICOND2BWP
    CLASS CORE ;
    FOREIGN FIICOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.805 0.350 4.865 0.805 ;
        RECT  4.795 0.185 4.805 1.035 ;
        RECT  4.735 0.185 4.795 0.465 ;
        RECT  4.735 0.735 4.795 1.035 ;
        END
    END S
    PIN CON1
        ANTENNADIFFAREA 0.1442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.340 1.515 0.410 ;
        RECT  1.295 0.340 1.365 0.790 ;
        RECT  1.085 0.720 1.295 0.790 ;
        RECT  1.010 0.350 1.085 0.790 ;
        RECT  0.950 0.350 1.010 0.420 ;
        END
    END CON1
    PIN CON0
        ANTENNADIFFAREA 0.1582 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.710 0.690 0.780 ;
        RECT  0.415 0.185 0.485 0.465 ;
        RECT  0.385 0.355 0.415 0.465 ;
        RECT  0.315 0.355 0.385 0.780 ;
        RECT  0.175 0.690 0.315 0.780 ;
        END
    END CON0
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.365 0.495 4.455 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1640 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.980 3.010 1.075 ;
        RECT  2.205 0.980 2.880 1.050 ;
        RECT  2.135 0.850 2.205 1.050 ;
        RECT  1.510 0.850 2.135 0.920 ;
        RECT  1.505 0.495 1.510 0.920 ;
        RECT  1.435 0.495 1.505 0.930 ;
        RECT  0.875 0.860 1.435 0.930 ;
        RECT  0.805 0.520 0.875 0.930 ;
        RECT  0.105 0.850 0.805 0.920 ;
        RECT  0.105 0.495 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.920 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.665 0.550 1.840 0.620 ;
        RECT  1.595 0.200 1.665 0.620 ;
        RECT  1.225 0.200 1.595 0.270 ;
        RECT  1.155 0.200 1.225 0.640 ;
        RECT  0.665 0.200 1.155 0.270 ;
        RECT  0.590 0.200 0.665 0.615 ;
        RECT  0.470 0.545 0.590 0.615 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.000 -0.115 5.040 0.115 ;
        RECT  4.900 -0.115 5.000 0.270 ;
        RECT  4.640 -0.115 4.900 0.115 ;
        RECT  4.520 -0.115 4.640 0.140 ;
        RECT  4.260 -0.115 4.520 0.115 ;
        RECT  4.140 -0.115 4.260 0.140 ;
        RECT  3.285 -0.115 4.140 0.115 ;
        RECT  3.215 -0.115 3.285 0.450 ;
        RECT  2.400 -0.115 3.215 0.115 ;
        RECT  2.280 -0.115 2.400 0.140 ;
        RECT  2.020 -0.115 2.280 0.115 ;
        RECT  1.900 -0.115 2.020 0.140 ;
        RECT  1.640 -0.115 1.900 0.115 ;
        RECT  1.520 -0.115 1.640 0.130 ;
        RECT  1.260 -0.115 1.520 0.115 ;
        RECT  1.140 -0.115 1.260 0.130 ;
        RECT  0.880 -0.115 1.140 0.115 ;
        RECT  0.760 -0.115 0.880 0.130 ;
        RECT  0.140 -0.115 0.760 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 1.145 5.040 1.375 ;
        RECT  4.915 0.895 4.985 1.375 ;
        RECT  4.615 1.145 4.915 1.375 ;
        RECT  4.545 0.700 4.615 1.375 ;
        RECT  4.260 1.145 4.545 1.375 ;
        RECT  4.140 1.025 4.260 1.375 ;
        RECT  3.310 1.145 4.140 1.375 ;
        RECT  3.190 0.995 3.310 1.375 ;
        RECT  2.390 1.145 3.190 1.375 ;
        RECT  2.270 1.120 2.390 1.375 ;
        RECT  2.000 1.145 2.270 1.375 ;
        RECT  1.880 1.005 2.000 1.375 ;
        RECT  1.620 1.145 1.880 1.375 ;
        RECT  1.500 1.005 1.620 1.375 ;
        RECT  0.880 1.145 1.500 1.375 ;
        RECT  0.760 1.005 0.880 1.375 ;
        RECT  0.510 1.145 0.760 1.375 ;
        RECT  0.390 1.005 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.990 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.640 0.545 4.720 0.615 ;
        RECT  4.570 0.210 4.640 0.615 ;
        RECT  3.845 0.210 4.570 0.280 ;
        RECT  4.285 0.350 4.450 0.420 ;
        RECT  4.285 0.885 4.450 0.955 ;
        RECT  4.215 0.350 4.285 0.955 ;
        RECT  4.085 0.520 4.215 0.640 ;
        RECT  4.035 0.885 4.215 0.955 ;
        RECT  4.010 0.355 4.070 0.425 ;
        RECT  4.010 0.735 4.060 0.805 ;
        RECT  3.965 0.885 4.035 1.040 ;
        RECT  3.940 0.355 4.010 0.805 ;
        RECT  3.700 0.970 3.965 1.040 ;
        RECT  3.775 0.210 3.845 0.890 ;
        RECT  3.630 0.325 3.700 1.040 ;
        RECT  3.580 0.325 3.630 0.445 ;
        RECT  3.550 0.970 3.630 1.040 ;
        RECT  3.500 0.520 3.560 0.640 ;
        RECT  3.465 0.185 3.500 0.835 ;
        RECT  3.430 0.185 3.465 1.045 ;
        RECT  3.395 0.185 3.430 0.445 ;
        RECT  3.395 0.755 3.430 1.045 ;
        RECT  3.300 0.520 3.360 0.640 ;
        RECT  3.230 0.520 3.300 0.910 ;
        RECT  2.725 0.840 3.230 0.910 ;
        RECT  3.105 0.695 3.130 0.765 ;
        RECT  3.035 0.185 3.105 0.765 ;
        RECT  3.010 0.510 3.035 0.765 ;
        RECT  2.950 0.510 3.010 0.630 ;
        RECT  2.880 0.210 2.950 0.280 ;
        RECT  2.880 0.700 2.930 0.770 ;
        RECT  2.810 0.210 2.880 0.770 ;
        RECT  1.990 0.210 2.810 0.280 ;
        RECT  2.655 0.350 2.725 0.910 ;
        RECT  2.500 0.365 2.570 0.910 ;
        RECT  2.090 0.365 2.500 0.435 ;
        RECT  2.450 0.710 2.500 0.910 ;
        RECT  2.070 0.710 2.450 0.780 ;
        RECT  1.990 0.540 2.215 0.620 ;
        RECT  1.920 0.210 1.990 0.780 ;
        RECT  1.805 0.210 1.920 0.280 ;
        RECT  1.680 0.710 1.920 0.780 ;
        RECT  1.735 0.210 1.805 0.470 ;
    END
END FIICOND2BWP

MACRO FILL16BWP
    CLASS CORE ;
    FOREIGN FILL16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.240 1.375 ;
        END
    END VDD
END FILL16BWP

MACRO FILL1BWP
    CLASS CORE ;
    FOREIGN FILL1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.140 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.140 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.140 1.375 ;
        END
    END VDD
END FILL1BWP

MACRO FILL2BWP
    CLASS CORE ;
    FOREIGN FILL2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.280 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.280 1.375 ;
        END
    END VDD
END FILL2BWP

MACRO FILL32BWP
    CLASS CORE ;
    FOREIGN FILL32BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.480 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 4.480 1.375 ;
        END
    END VDD
END FILL32BWP

MACRO FILL3BWP
    CLASS CORE ;
    FOREIGN FILL3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
END FILL3BWP

MACRO FILL4BWP
    CLASS CORE ;
    FOREIGN FILL4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.560 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.560 1.375 ;
        END
    END VDD
END FILL4BWP

MACRO FILL64BWP
    CLASS CORE ;
    FOREIGN FILL64BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 8.960 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 8.960 1.375 ;
        END
    END VDD
END FILL64BWP

MACRO FILL8BWP
    CLASS CORE ;
    FOREIGN FILL8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 1.120 1.375 ;
        END
    END VDD
END FILL8BWP

MACRO GAN2D1BWP
    CLASS CORE ;
    FOREIGN GAN2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.200 1.365 1.060 ;
        RECT  1.160 0.200 1.295 0.280 ;
        RECT  1.180 0.980 1.295 1.060 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.320 ;
        RECT  0.900 -0.115 1.010 0.115 ;
        RECT  0.820 -0.115 0.900 0.320 ;
        RECT  0.220 -0.115 0.820 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.900 1.145 0.990 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.600 1.145 0.820 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.200 1.145 0.480 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.500 1.225 0.785 ;
        RECT  0.945 0.715 1.155 0.785 ;
        RECT  0.875 0.500 0.945 0.785 ;
        RECT  0.665 0.715 0.875 0.785 ;
        RECT  0.595 0.200 0.665 0.915 ;
        RECT  0.480 0.200 0.595 0.280 ;
        RECT  0.270 0.845 0.595 0.915 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAN2D1BWP

MACRO GAN2D2BWP
    CLASS CORE ;
    FOREIGN GAN2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.370 1.365 0.880 ;
        RECT  1.100 0.370 1.295 0.440 ;
        RECT  1.085 0.810 1.295 0.880 ;
        RECT  1.015 0.190 1.100 0.440 ;
        RECT  1.015 0.810 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.300 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.220 -0.115 0.800 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.950 1.280 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.200 1.145 0.480 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.515 1.225 0.640 ;
        RECT  0.870 0.355 0.945 0.915 ;
        RECT  0.590 0.355 0.870 0.425 ;
        RECT  0.270 0.845 0.870 0.915 ;
        RECT  0.490 0.190 0.590 0.425 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAN2D2BWP

MACRO GAOI21D1BWP
    CLASS CORE ;
    FOREIGN GAOI21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2237 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.190 1.290 0.290 ;
        RECT  1.190 0.190 1.260 0.415 ;
        RECT  0.920 0.345 1.190 0.415 ;
        RECT  0.850 0.205 0.920 0.415 ;
        RECT  0.665 0.205 0.850 0.275 ;
        RECT  0.595 0.205 0.665 0.915 ;
        RECT  0.480 0.205 0.595 0.275 ;
        RECT  0.270 0.845 0.595 0.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 1.250 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.245 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 1.400 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.220 -0.115 0.990 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  0.990 0.850 1.110 1.375 ;
        RECT  0.000 1.145 0.990 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.970 1.300 1.070 ;
        RECT  1.190 0.710 1.260 1.070 ;
        RECT  0.920 0.710 1.190 0.780 ;
        RECT  0.850 0.710 0.920 1.055 ;
        RECT  0.080 0.985 0.850 1.055 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAOI21D1BWP

MACRO GAOI21D2BWP
    CLASS CORE ;
    FOREIGN GAOI21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3420 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.190 2.065 0.915 ;
        RECT  1.890 0.190 1.995 0.290 ;
        RECT  0.805 0.845 1.995 0.915 ;
        RECT  0.810 0.190 0.910 0.410 ;
        RECT  0.805 0.340 0.810 0.410 ;
        RECT  0.735 0.340 0.805 0.915 ;
        RECT  0.590 0.340 0.735 0.410 ;
        RECT  0.490 0.190 0.590 0.410 ;
        RECT  0.220 0.340 0.490 0.410 ;
        RECT  0.150 0.200 0.220 0.410 ;
        RECT  0.035 0.200 0.150 0.280 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.245 0.695 0.455 0.765 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.670 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.775 ;
        RECT  0.945 0.705 1.855 0.775 ;
        RECT  0.875 0.495 0.945 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.620 -0.115 2.100 0.115 ;
        RECT  1.500 -0.115 1.620 0.280 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.280 ;
        RECT  0.410 -0.115 1.180 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.145 2.100 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.600 0.985 2.020 1.055 ;
        RECT  1.700 0.185 1.800 0.405 ;
        RECT  1.000 0.185 1.100 0.405 ;
        RECT  0.480 0.850 0.600 1.055 ;
        RECT  0.100 0.850 0.210 1.070 ;
        LAYER VIA1 ;
        RECT  0.505 0.945 0.575 1.015 ;
        RECT  0.125 0.945 0.195 1.015 ;
        LAYER M2 ;
        RECT  0.075 0.945 0.625 1.015 ;
    END
END GAOI21D2BWP

MACRO GAOI22D1BWP
    CLASS CORE ;
    FOREIGN GAOI22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2448 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.990 1.365 1.060 ;
        RECT  0.805 0.200 0.920 0.275 ;
        RECT  0.735 0.200 0.805 1.060 ;
        RECT  0.480 0.200 0.735 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.640 ;
        RECT  1.155 0.495 1.295 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.220 -0.115 1.180 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 1.400 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.845 1.200 0.920 ;
        RECT  1.085 0.185 1.100 0.290 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.755 1.085 0.920 ;
        RECT  1.000 0.185 1.015 0.290 ;
        RECT  0.905 0.845 1.015 0.920 ;
        RECT  0.300 0.185 0.400 0.405 ;
        RECT  0.315 0.745 0.385 1.065 ;
        LAYER VIA1 ;
        RECT  1.015 0.805 1.085 0.875 ;
        RECT  0.315 0.805 0.385 0.875 ;
        LAYER M2 ;
        RECT  0.265 0.805 1.135 0.875 ;
    END
END GAOI22D1BWP

MACRO GBUFFD1BWP
    CLASS CORE ;
    FOREIGN GBUFFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.200 0.665 1.060 ;
        RECT  0.480 0.200 0.595 0.280 ;
        RECT  0.480 0.980 0.595 1.060 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.355 0.265 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.400 -0.115 0.700 0.115 ;
        RECT  0.300 -0.115 0.400 0.290 ;
        RECT  0.000 -0.115 0.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.145 0.700 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.500 0.525 0.780 ;
        RECT  0.105 0.710 0.450 0.780 ;
        RECT  0.105 0.200 0.220 0.280 ;
        RECT  0.105 0.980 0.220 1.060 ;
        RECT  0.035 0.200 0.105 1.060 ;
    END
END GBUFFD1BWP

MACRO GBUFFD2BWP
    CLASS CORE ;
    FOREIGN GBUFFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.365 1.365 0.845 ;
        RECT  1.100 0.365 1.295 0.435 ;
        RECT  1.085 0.775 1.295 0.845 ;
        RECT  1.015 0.190 1.100 0.435 ;
        RECT  1.015 0.775 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.545 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.290 0.290 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.210 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.210 0.290 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.515 1.225 0.640 ;
        RECT  0.870 0.350 0.945 0.780 ;
        RECT  0.400 0.350 0.870 0.420 ;
        RECT  0.385 0.710 0.870 0.780 ;
        RECT  0.300 0.190 0.400 0.420 ;
        RECT  0.315 0.710 0.385 0.965 ;
    END
END GBUFFD2BWP

MACRO GBUFFD3BWP
    CLASS CORE ;
    FOREIGN GBUFFD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.2376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.360 1.365 0.920 ;
        RECT  1.100 0.360 1.295 0.430 ;
        RECT  0.590 0.850 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.430 ;
        RECT  0.590 0.360 1.000 0.430 ;
        RECT  0.490 0.190 0.590 0.430 ;
        RECT  0.490 0.850 0.590 1.070 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.355 0.265 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.290 0.290 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.390 -0.115 0.800 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.400 1.375 ;
        RECT  1.180 0.990 1.300 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.410 1.145 0.800 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.510 1.225 0.780 ;
        RECT  0.950 0.710 1.155 0.780 ;
        RECT  0.870 0.510 0.950 0.780 ;
        RECT  0.530 0.710 0.870 0.780 ;
        RECT  0.450 0.510 0.530 0.780 ;
        RECT  0.105 0.710 0.450 0.780 ;
        RECT  0.105 0.200 0.220 0.280 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.200 0.105 1.070 ;
    END
END GBUFFD3BWP

MACRO GBUFFD4BWP
    CLASS CORE ;
    FOREIGN GBUFFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.2304 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.370 2.065 0.875 ;
        RECT  1.800 0.370 1.995 0.440 ;
        RECT  1.785 0.805 1.995 0.875 ;
        RECT  1.700 0.190 1.800 0.440 ;
        RECT  1.715 0.805 1.785 0.965 ;
        RECT  1.085 0.805 1.715 0.875 ;
        RECT  1.100 0.370 1.700 0.440 ;
        RECT  1.015 0.190 1.100 0.440 ;
        RECT  1.015 0.805 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.665 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 -0.115 2.100 0.115 ;
        RECT  1.900 -0.115 1.980 0.300 ;
        RECT  1.620 -0.115 1.900 0.115 ;
        RECT  1.500 -0.115 1.620 0.280 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.280 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.200 -0.115 0.480 0.115 ;
        RECT  0.120 -0.115 0.200 0.320 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.145 2.100 1.375 ;
        RECT  1.900 0.960 1.980 1.375 ;
        RECT  1.600 1.145 1.900 1.375 ;
        RECT  1.520 0.960 1.600 1.375 ;
        RECT  1.280 1.145 1.520 1.375 ;
        RECT  1.200 0.960 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.960 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.960 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.935 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.515 1.925 0.640 ;
        RECT  0.870 0.355 0.945 0.875 ;
        RECT  0.400 0.355 0.870 0.425 ;
        RECT  0.385 0.805 0.870 0.875 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.315 0.805 0.385 0.965 ;
    END
END GBUFFD4BWP

MACRO GBUFFD8BWP
    CLASS CORE ;
    FOREIGN GBUFFD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.4608 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.370 4.165 0.875 ;
        RECT  3.900 0.370 4.095 0.440 ;
        RECT  3.885 0.805 4.095 0.875 ;
        RECT  3.800 0.190 3.900 0.440 ;
        RECT  3.815 0.805 3.885 0.965 ;
        RECT  3.185 0.805 3.815 0.875 ;
        RECT  3.200 0.370 3.800 0.440 ;
        RECT  3.100 0.190 3.200 0.440 ;
        RECT  3.115 0.805 3.185 0.965 ;
        RECT  2.485 0.805 3.115 0.875 ;
        RECT  2.500 0.370 3.100 0.440 ;
        RECT  2.400 0.190 2.500 0.440 ;
        RECT  2.415 0.805 2.485 0.965 ;
        RECT  1.785 0.805 2.415 0.875 ;
        RECT  1.800 0.370 2.400 0.440 ;
        RECT  1.715 0.190 1.800 0.440 ;
        RECT  1.715 0.805 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 1.295 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.080 -0.115 4.200 0.115 ;
        RECT  4.000 -0.115 4.080 0.300 ;
        RECT  3.720 -0.115 4.000 0.115 ;
        RECT  3.600 -0.115 3.720 0.280 ;
        RECT  3.410 -0.115 3.600 0.115 ;
        RECT  3.280 -0.115 3.410 0.280 ;
        RECT  3.020 -0.115 3.280 0.115 ;
        RECT  2.900 -0.115 3.020 0.280 ;
        RECT  2.700 -0.115 2.900 0.115 ;
        RECT  2.580 -0.115 2.700 0.280 ;
        RECT  2.320 -0.115 2.580 0.115 ;
        RECT  2.200 -0.115 2.320 0.280 ;
        RECT  2.000 -0.115 2.200 0.115 ;
        RECT  1.880 -0.115 2.000 0.280 ;
        RECT  1.620 -0.115 1.880 0.115 ;
        RECT  1.500 -0.115 1.620 0.280 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.280 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.200 -0.115 0.480 0.115 ;
        RECT  0.120 -0.115 0.200 0.320 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.080 1.145 4.200 1.375 ;
        RECT  4.000 0.960 4.080 1.375 ;
        RECT  3.700 1.145 4.000 1.375 ;
        RECT  3.620 0.960 3.700 1.375 ;
        RECT  3.380 1.145 3.620 1.375 ;
        RECT  3.300 0.960 3.380 1.375 ;
        RECT  3.000 1.145 3.300 1.375 ;
        RECT  2.920 0.960 3.000 1.375 ;
        RECT  2.680 1.145 2.920 1.375 ;
        RECT  2.600 0.960 2.680 1.375 ;
        RECT  2.300 1.145 2.600 1.375 ;
        RECT  2.220 0.960 2.300 1.375 ;
        RECT  1.980 1.145 2.220 1.375 ;
        RECT  1.900 0.960 1.980 1.375 ;
        RECT  1.600 1.145 1.900 1.375 ;
        RECT  1.520 0.960 1.600 1.375 ;
        RECT  1.280 1.145 1.520 1.375 ;
        RECT  1.200 0.960 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.960 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.960 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.935 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.515 4.025 0.640 ;
        RECT  1.570 0.355 1.645 0.875 ;
        RECT  1.100 0.355 1.570 0.425 ;
        RECT  1.085 0.805 1.570 0.875 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  1.015 0.805 1.085 0.965 ;
        RECT  0.385 0.805 1.015 0.875 ;
        RECT  0.400 0.355 1.000 0.425 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.315 0.805 0.385 0.965 ;
    END
END GBUFFD8BWP

MACRO GDCAP10BWP
    CLASS CORE ;
    FOREIGN GDCAP10BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.690 -0.115 7.000 0.115 ;
        RECT  6.610 -0.115 6.690 0.300 ;
        RECT  6.500 -0.115 6.610 0.115 ;
        RECT  6.420 -0.115 6.500 0.300 ;
        RECT  5.990 -0.115 6.420 0.115 ;
        RECT  5.910 -0.115 5.990 0.300 ;
        RECT  5.800 -0.115 5.910 0.115 ;
        RECT  5.720 -0.115 5.800 0.300 ;
        RECT  5.290 -0.115 5.720 0.115 ;
        RECT  5.210 -0.115 5.290 0.300 ;
        RECT  5.100 -0.115 5.210 0.115 ;
        RECT  5.020 -0.115 5.100 0.300 ;
        RECT  4.590 -0.115 5.020 0.115 ;
        RECT  4.510 -0.115 4.590 0.300 ;
        RECT  4.400 -0.115 4.510 0.115 ;
        RECT  4.320 -0.115 4.400 0.300 ;
        RECT  3.890 -0.115 4.320 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.700 -0.115 3.810 0.115 ;
        RECT  3.620 -0.115 3.700 0.300 ;
        RECT  3.190 -0.115 3.620 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  3.000 -0.115 3.110 0.115 ;
        RECT  2.920 -0.115 3.000 0.300 ;
        RECT  2.490 -0.115 2.920 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.300 -0.115 2.410 0.115 ;
        RECT  2.220 -0.115 2.300 0.300 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.600 -0.115 1.710 0.115 ;
        RECT  1.520 -0.115 1.600 0.300 ;
        RECT  1.090 -0.115 1.520 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.900 -0.115 1.010 0.115 ;
        RECT  0.820 -0.115 0.900 0.300 ;
        RECT  0.390 -0.115 0.820 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.200 -0.115 0.310 0.115 ;
        RECT  0.120 -0.115 0.200 0.300 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.880 1.145 7.000 1.375 ;
        RECT  6.800 0.850 6.880 1.375 ;
        RECT  6.590 0.850 6.800 0.920 ;
        RECT  6.180 1.145 6.800 1.375 ;
        RECT  6.100 0.850 6.180 1.375 ;
        RECT  5.890 0.850 6.100 0.920 ;
        RECT  5.480 1.145 6.100 1.375 ;
        RECT  5.400 0.850 5.480 1.375 ;
        RECT  5.190 0.850 5.400 0.920 ;
        RECT  4.780 1.145 5.400 1.375 ;
        RECT  4.700 0.850 4.780 1.375 ;
        RECT  4.490 0.850 4.700 0.920 ;
        RECT  4.080 1.145 4.700 1.375 ;
        RECT  4.000 0.850 4.080 1.375 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.380 1.145 4.000 1.375 ;
        RECT  3.300 0.850 3.380 1.375 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  2.680 1.145 3.300 1.375 ;
        RECT  2.600 0.850 2.680 1.375 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  1.980 1.145 2.600 1.375 ;
        RECT  1.900 0.850 1.980 1.375 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.280 1.145 1.900 1.375 ;
        RECT  1.200 0.850 1.280 1.375 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.580 1.145 1.200 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.790 0.190 6.900 0.450 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.550 0.380 6.790 0.450 ;
        RECT  6.510 0.710 6.745 0.780 ;
        RECT  6.470 0.380 6.550 0.640 ;
        RECT  6.410 0.710 6.510 1.070 ;
        RECT  6.190 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.410 0.780 ;
        RECT  6.090 0.190 6.190 0.450 ;
        RECT  6.050 0.520 6.130 0.780 ;
        RECT  5.850 0.380 6.090 0.450 ;
        RECT  5.810 0.710 6.050 0.780 ;
        RECT  5.770 0.380 5.850 0.640 ;
        RECT  5.710 0.710 5.810 1.070 ;
        RECT  5.490 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.710 0.780 ;
        RECT  5.390 0.190 5.490 0.450 ;
        RECT  5.350 0.520 5.430 0.780 ;
        RECT  5.150 0.380 5.390 0.450 ;
        RECT  5.110 0.710 5.350 0.780 ;
        RECT  5.070 0.380 5.150 0.640 ;
        RECT  5.010 0.710 5.110 1.070 ;
        RECT  4.790 0.380 5.070 0.450 ;
        RECT  4.735 0.710 5.010 0.780 ;
        RECT  4.690 0.190 4.790 0.450 ;
        RECT  4.650 0.520 4.735 0.780 ;
        RECT  4.450 0.380 4.690 0.450 ;
        RECT  4.410 0.710 4.650 0.780 ;
        RECT  4.370 0.380 4.450 0.640 ;
        RECT  4.310 0.710 4.410 1.070 ;
        RECT  4.090 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.310 0.780 ;
        RECT  3.990 0.190 4.090 0.450 ;
        RECT  3.950 0.520 4.030 0.780 ;
        RECT  3.750 0.380 3.990 0.450 ;
        RECT  3.710 0.710 3.950 0.780 ;
        RECT  3.670 0.380 3.750 0.640 ;
        RECT  3.610 0.710 3.710 1.070 ;
        RECT  3.390 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.610 0.780 ;
        RECT  3.290 0.190 3.390 0.450 ;
        RECT  3.250 0.520 3.330 0.780 ;
        RECT  3.050 0.380 3.290 0.450 ;
        RECT  3.010 0.710 3.250 0.780 ;
        RECT  2.970 0.380 3.050 0.640 ;
        RECT  2.910 0.710 3.010 1.070 ;
        RECT  2.690 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.910 0.780 ;
        RECT  2.590 0.190 2.690 0.450 ;
        RECT  2.550 0.520 2.630 0.780 ;
        RECT  2.350 0.380 2.590 0.450 ;
        RECT  2.310 0.710 2.550 0.780 ;
        RECT  2.270 0.380 2.350 0.640 ;
        RECT  2.210 0.710 2.310 1.070 ;
        RECT  1.990 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.210 0.780 ;
        RECT  1.890 0.190 1.990 0.450 ;
        RECT  1.850 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.610 0.710 1.850 0.780 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GDCAP10BWP

MACRO GDCAP2BWP
    CLASS CORE ;
    FOREIGN GDCAP2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.900 -0.115 1.010 0.115 ;
        RECT  0.820 -0.115 0.900 0.300 ;
        RECT  0.390 -0.115 0.820 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.200 -0.115 0.310 0.115 ;
        RECT  0.120 -0.115 0.200 0.300 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.850 1.280 1.375 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.580 1.145 1.200 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.190 1.300 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.910 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GDCAP2BWP

MACRO GDCAP3BWP
    CLASS CORE ;
    FOREIGN GDCAP3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 -0.115 2.100 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.600 -0.115 1.710 0.115 ;
        RECT  1.520 -0.115 1.600 0.300 ;
        RECT  1.090 -0.115 1.520 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.900 -0.115 1.010 0.115 ;
        RECT  0.820 -0.115 0.900 0.300 ;
        RECT  0.390 -0.115 0.820 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.200 -0.115 0.310 0.115 ;
        RECT  0.120 -0.115 0.200 0.300 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.145 2.100 1.375 ;
        RECT  1.900 0.850 1.980 1.375 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.280 1.145 1.900 1.375 ;
        RECT  1.200 0.850 1.280 1.375 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.580 1.145 1.200 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.890 0.190 2.000 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.610 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GDCAP3BWP

MACRO GDCAP4BWP
    CLASS CORE ;
    FOREIGN GDCAP4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.490 -0.115 2.800 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.300 -0.115 2.410 0.115 ;
        RECT  2.220 -0.115 2.300 0.300 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.600 -0.115 1.710 0.115 ;
        RECT  1.520 -0.115 1.600 0.300 ;
        RECT  1.090 -0.115 1.520 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.900 -0.115 1.010 0.115 ;
        RECT  0.820 -0.115 0.900 0.300 ;
        RECT  0.390 -0.115 0.820 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.200 -0.115 0.310 0.115 ;
        RECT  0.120 -0.115 0.200 0.300 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 1.145 2.800 1.375 ;
        RECT  2.600 0.850 2.680 1.375 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  1.980 1.145 2.600 1.375 ;
        RECT  1.900 0.850 1.980 1.375 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.280 1.145 1.900 1.375 ;
        RECT  1.200 0.850 1.280 1.375 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.580 1.145 1.200 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.590 0.190 2.700 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.350 0.380 2.590 0.450 ;
        RECT  2.310 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.350 0.640 ;
        RECT  2.210 0.710 2.310 1.070 ;
        RECT  1.990 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.210 0.780 ;
        RECT  1.890 0.190 1.990 0.450 ;
        RECT  1.850 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.610 0.710 1.850 0.780 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GDCAP4BWP

MACRO GDCAPBWP
    CLASS CORE ;
    FOREIGN GDCAPBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.390 -0.115 0.700 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.200 -0.115 0.310 0.115 ;
        RECT  0.120 -0.115 0.200 0.300 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.700 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.490 0.190 0.600 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.210 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GDCAPBWP

MACRO GDFCNQD1BWP
    CLASS CORE ;
    FOREIGN GDFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.205 4.865 1.055 ;
        RECT  4.680 0.205 4.795 0.275 ;
        RECT  4.680 0.985 4.795 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.610 0.665 1.275 0.735 ;
        LAYER M1 ;
        RECT  0.675 0.665 0.760 0.735 ;
        RECT  0.605 0.665 0.675 0.785 ;
        RECT  0.245 0.715 0.605 0.785 ;
        RECT  0.175 0.495 0.245 0.785 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.395 0.665 4.075 0.735 ;
        RECT  2.325 0.525 2.395 0.735 ;
        RECT  1.940 0.525 2.325 0.595 ;
        LAYER M1 ;
        RECT  3.955 0.355 4.025 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.610 -0.115 4.900 0.115 ;
        RECT  4.490 -0.115 4.610 0.270 ;
        RECT  3.700 -0.115 4.490 0.115 ;
        RECT  3.615 -0.115 3.700 0.315 ;
        RECT  2.495 -0.115 3.615 0.115 ;
        RECT  2.420 -0.115 2.495 0.315 ;
        RECT  2.000 -0.115 2.420 0.115 ;
        RECT  1.910 -0.115 2.000 0.310 ;
        RECT  0.410 -0.115 1.910 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.610 1.145 4.900 1.375 ;
        RECT  4.520 0.805 4.610 1.375 ;
        RECT  3.890 1.145 4.520 1.375 ;
        RECT  3.815 0.820 3.890 1.375 ;
        RECT  2.510 1.145 3.815 1.375 ;
        RECT  2.390 0.850 2.510 1.375 ;
        RECT  1.810 1.145 2.390 1.375 ;
        RECT  1.690 0.850 1.810 1.375 ;
        RECT  0.410 1.145 1.690 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.520 4.725 0.640 ;
        RECT  4.375 0.520 4.445 0.905 ;
        RECT  4.305 0.205 4.420 0.275 ;
        RECT  4.305 0.985 4.420 1.055 ;
        RECT  4.235 0.205 4.305 1.055 ;
        RECT  4.095 0.205 4.165 1.055 ;
        RECT  3.980 0.205 4.095 0.275 ;
        RECT  3.980 0.985 4.095 1.055 ;
        RECT  3.885 0.195 3.910 0.290 ;
        RECT  3.780 0.195 3.885 0.475 ;
        RECT  3.535 0.545 3.820 0.615 ;
        RECT  3.610 0.770 3.710 1.070 ;
        RECT  3.515 0.385 3.655 0.455 ;
        RECT  3.465 0.545 3.535 0.780 ;
        RECT  3.445 0.200 3.515 0.455 ;
        RECT  3.185 0.710 3.465 0.780 ;
        RECT  3.275 0.200 3.445 0.280 ;
        RECT  3.290 0.850 3.390 1.070 ;
        RECT  3.255 0.385 3.345 0.640 ;
        RECT  3.185 0.185 3.205 0.315 ;
        RECT  3.115 0.185 3.185 0.965 ;
        RECT  2.975 0.185 3.045 0.370 ;
        RECT  2.975 0.520 3.045 0.905 ;
        RECT  2.905 0.985 3.015 1.055 ;
        RECT  2.835 0.185 2.975 0.275 ;
        RECT  2.835 0.355 2.905 1.055 ;
        RECT  2.695 0.205 2.765 1.055 ;
        RECT  2.580 0.205 2.695 0.275 ;
        RECT  2.580 0.985 2.695 1.055 ;
        RECT  2.555 0.485 2.625 0.765 ;
        RECT  1.225 0.695 2.555 0.765 ;
        RECT  2.345 0.545 2.395 0.615 ;
        RECT  2.275 0.345 2.345 0.615 ;
        RECT  2.160 0.190 2.325 0.270 ;
        RECT  2.210 0.850 2.310 1.070 ;
        RECT  2.250 0.545 2.275 0.615 ;
        RECT  1.800 0.515 2.170 0.615 ;
        RECT  2.090 0.190 2.160 0.365 ;
        RECT  1.890 0.850 1.990 1.070 ;
        RECT  1.690 0.185 1.810 0.395 ;
        RECT  1.365 0.515 1.695 0.615 ;
        RECT  1.180 0.205 1.620 0.275 ;
        RECT  1.510 0.850 1.610 1.070 ;
        RECT  1.295 0.355 1.365 0.615 ;
        RECT  1.190 0.850 1.290 1.070 ;
        RECT  1.155 0.520 1.225 0.765 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.870 0.355 0.945 0.645 ;
        RECT  0.480 0.205 0.920 0.275 ;
        RECT  0.790 0.805 0.920 1.075 ;
        RECT  0.420 0.355 0.870 0.425 ;
        RECT  0.570 0.865 0.665 1.075 ;
        RECT  0.480 0.960 0.570 1.075 ;
        RECT  0.350 0.345 0.420 0.425 ;
        RECT  0.210 0.345 0.350 0.415 ;
        RECT  0.105 0.985 0.220 1.055 ;
        RECT  0.110 0.190 0.210 0.415 ;
        RECT  0.105 0.345 0.110 0.415 ;
        RECT  0.035 0.345 0.105 1.055 ;
        LAYER VIA1 ;
        RECT  4.375 0.805 4.445 0.875 ;
        RECT  4.235 0.245 4.305 0.315 ;
        RECT  4.235 0.945 4.305 1.015 ;
        RECT  4.095 0.805 4.165 0.875 ;
        RECT  3.955 0.665 4.025 0.735 ;
        RECT  3.625 0.805 3.695 0.875 ;
        RECT  3.535 0.385 3.605 0.455 ;
        RECT  3.305 0.945 3.375 1.015 ;
        RECT  3.255 0.525 3.325 0.595 ;
        RECT  2.975 0.245 3.045 0.315 ;
        RECT  2.975 0.805 3.045 0.875 ;
        RECT  2.835 0.385 2.905 0.455 ;
        RECT  2.835 0.945 2.905 1.015 ;
        RECT  2.695 0.805 2.765 0.875 ;
        RECT  2.555 0.525 2.625 0.595 ;
        RECT  2.275 0.385 2.345 0.455 ;
        RECT  2.225 0.945 2.295 1.015 ;
        RECT  2.090 0.245 2.160 0.315 ;
        RECT  1.995 0.525 2.065 0.595 ;
        RECT  1.905 0.945 1.975 1.015 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.295 0.385 1.365 0.455 ;
        RECT  1.205 0.945 1.275 1.015 ;
        RECT  1.155 0.665 1.225 0.735 ;
        RECT  1.015 0.525 1.085 0.595 ;
        RECT  0.820 0.805 0.890 0.875 ;
        RECT  0.660 0.665 0.730 0.735 ;
        RECT  0.595 0.895 0.665 0.965 ;
        LAYER M2 ;
        RECT  3.575 0.805 4.495 0.875 ;
        RECT  2.925 0.245 4.355 0.315 ;
        RECT  3.255 0.945 4.355 1.015 ;
        RECT  2.625 0.385 3.655 0.455 ;
        RECT  2.505 0.525 3.375 0.595 ;
        RECT  2.645 0.805 3.095 0.875 ;
        RECT  2.175 0.945 2.955 1.015 ;
        RECT  2.555 0.245 2.625 0.455 ;
        RECT  1.645 0.245 2.555 0.315 ;
        RECT  1.785 0.385 2.395 0.455 ;
        RECT  1.505 0.945 2.025 1.015 ;
        RECT  1.715 0.385 1.785 0.595 ;
        RECT  0.965 0.525 1.715 0.595 ;
        RECT  1.575 0.245 1.645 0.455 ;
        RECT  1.245 0.385 1.575 0.455 ;
        RECT  1.435 0.805 1.505 1.015 ;
        RECT  0.770 0.805 1.435 0.875 ;
        RECT  0.665 0.945 1.325 1.015 ;
        RECT  0.595 0.840 0.665 1.015 ;
    END
END GDFCNQD1BWP

MACRO GDFQD1BWP
    CLASS CORE ;
    FOREIGN GDFQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.205 4.165 1.055 ;
        RECT  3.980 0.205 4.095 0.275 ;
        RECT  3.980 0.985 4.095 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.125 0.385 2.880 0.455 ;
        LAYER M1 ;
        RECT  0.175 0.355 0.245 0.685 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 -0.115 4.200 0.115 ;
        RECT  3.790 -0.115 3.910 0.275 ;
        RECT  3.190 -0.115 3.790 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  1.810 -0.115 3.110 0.115 ;
        RECT  1.690 -0.115 1.810 0.275 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 1.145 4.200 1.375 ;
        RECT  3.790 0.850 3.910 1.375 ;
        RECT  3.210 1.145 3.790 1.375 ;
        RECT  3.090 0.850 3.210 1.375 ;
        RECT  1.810 1.145 3.090 1.375 ;
        RECT  1.690 0.850 1.810 1.375 ;
        RECT  0.400 1.145 1.690 1.375 ;
        RECT  0.300 0.835 0.400 1.375 ;
        RECT  0.000 1.145 0.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.955 0.355 4.025 0.780 ;
        RECT  3.710 0.355 3.955 0.425 ;
        RECT  3.710 0.710 3.955 0.780 ;
        RECT  3.535 0.510 3.755 0.640 ;
        RECT  3.610 0.190 3.710 0.425 ;
        RECT  3.640 0.710 3.710 1.070 ;
        RECT  3.610 0.970 3.640 1.070 ;
        RECT  3.395 0.200 3.465 1.055 ;
        RECT  3.280 0.200 3.395 0.275 ;
        RECT  3.280 0.985 3.395 1.055 ;
        RECT  3.255 0.450 3.325 0.780 ;
        RECT  3.115 0.380 3.185 0.780 ;
        RECT  3.010 0.380 3.115 0.450 ;
        RECT  3.010 0.710 3.115 0.780 ;
        RECT  2.860 0.520 3.045 0.640 ;
        RECT  2.940 0.190 3.010 0.450 ;
        RECT  2.910 0.710 3.010 1.070 ;
        RECT  2.910 0.190 2.940 0.290 ;
        RECT  2.625 0.710 2.910 0.780 ;
        RECT  2.790 0.385 2.860 0.640 ;
        RECT  2.580 0.195 2.800 0.315 ;
        RECT  2.730 0.385 2.790 0.455 ;
        RECT  2.590 0.850 2.690 1.070 ;
        RECT  2.555 0.520 2.625 0.780 ;
        RECT  2.485 0.190 2.500 0.290 ;
        RECT  2.415 0.190 2.485 0.965 ;
        RECT  2.400 0.190 2.415 0.290 ;
        RECT  2.255 0.355 2.345 0.640 ;
        RECT  2.065 0.205 2.320 0.275 ;
        RECT  2.210 0.775 2.310 1.070 ;
        RECT  1.995 0.205 2.065 0.930 ;
        RECT  1.880 0.205 1.995 0.275 ;
        RECT  1.650 0.360 1.995 0.430 ;
        RECT  1.990 0.860 1.995 0.930 ;
        RECT  1.890 0.860 1.990 1.070 ;
        RECT  1.835 0.510 1.925 0.780 ;
        RECT  1.570 0.360 1.650 0.640 ;
        RECT  1.180 0.205 1.620 0.275 ;
        RECT  1.510 0.775 1.610 1.070 ;
        RECT  1.190 0.775 1.290 1.070 ;
        RECT  1.160 0.355 1.250 0.640 ;
        RECT  1.090 0.190 1.100 0.290 ;
        RECT  1.020 0.190 1.090 0.965 ;
        RECT  1.000 0.190 1.020 0.290 ;
        RECT  0.810 0.775 0.950 1.070 ;
        RECT  0.705 0.520 0.945 0.640 ;
        RECT  0.480 0.205 0.920 0.275 ;
        RECT  0.610 0.520 0.705 0.905 ;
        RECT  0.540 0.980 0.620 1.070 ;
        RECT  0.470 0.845 0.540 1.070 ;
        RECT  0.105 0.205 0.220 0.275 ;
        RECT  0.110 0.800 0.210 1.070 ;
        RECT  0.105 0.800 0.110 0.880 ;
        RECT  0.035 0.205 0.105 0.880 ;
        LAYER VIA1 ;
        RECT  3.955 0.665 4.025 0.735 ;
        RECT  3.605 0.525 3.675 0.595 ;
        RECT  3.395 0.245 3.465 0.315 ;
        RECT  3.395 0.805 3.465 0.875 ;
        RECT  3.255 0.665 3.325 0.735 ;
        RECT  2.760 0.385 2.830 0.455 ;
        RECT  2.620 0.245 2.690 0.315 ;
        RECT  2.605 0.945 2.675 1.015 ;
        RECT  2.415 0.525 2.485 0.595 ;
        RECT  2.265 0.385 2.335 0.455 ;
        RECT  2.225 0.805 2.295 0.875 ;
        RECT  1.910 0.945 1.980 1.015 ;
        RECT  1.855 0.665 1.925 0.735 ;
        RECT  1.525 0.805 1.595 0.875 ;
        RECT  1.205 0.945 1.275 1.015 ;
        RECT  1.160 0.385 1.230 0.455 ;
        RECT  1.020 0.665 1.090 0.735 ;
        RECT  0.880 0.805 0.950 0.875 ;
        RECT  0.610 0.805 0.680 0.875 ;
        RECT  0.470 0.945 0.540 1.015 ;
        RECT  0.175 0.385 0.245 0.455 ;
        RECT  0.100 0.805 0.170 0.875 ;
        LAYER M2 ;
        RECT  3.205 0.665 4.075 0.735 ;
        RECT  2.365 0.525 3.725 0.595 ;
        RECT  2.570 0.245 3.515 0.315 ;
        RECT  2.175 0.805 3.515 0.875 ;
        RECT  1.860 0.945 2.725 1.015 ;
        RECT  0.970 0.665 1.975 0.735 ;
        RECT  0.830 0.805 1.645 0.875 ;
        RECT  0.420 0.945 1.325 1.015 ;
        RECT  0.050 0.805 0.730 0.875 ;
    END
END GDFQD1BWP

MACRO GFILL10BWP
    CLASS CORE ;
    FOREIGN GFILL10BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 7.000 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 7.000 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.790 0.190 6.900 0.450 ;
        RECT  6.790 0.850 6.900 1.070 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.550 0.380 6.790 0.450 ;
        RECT  6.590 0.850 6.790 0.920 ;
        RECT  6.510 0.710 6.745 0.780 ;
        RECT  6.380 0.200 6.710 0.280 ;
        RECT  6.470 0.380 6.550 0.640 ;
        RECT  6.410 0.710 6.510 1.070 ;
        RECT  6.190 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.410 0.780 ;
        RECT  6.090 0.190 6.190 0.450 ;
        RECT  6.090 0.850 6.190 1.070 ;
        RECT  6.050 0.520 6.130 0.780 ;
        RECT  5.850 0.380 6.090 0.450 ;
        RECT  5.890 0.850 6.090 0.920 ;
        RECT  5.810 0.710 6.050 0.780 ;
        RECT  5.680 0.200 6.010 0.280 ;
        RECT  5.770 0.380 5.850 0.640 ;
        RECT  5.710 0.710 5.810 1.070 ;
        RECT  5.490 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.710 0.780 ;
        RECT  5.390 0.190 5.490 0.450 ;
        RECT  5.390 0.850 5.490 1.070 ;
        RECT  5.350 0.520 5.430 0.780 ;
        RECT  5.150 0.380 5.390 0.450 ;
        RECT  5.190 0.850 5.390 0.920 ;
        RECT  5.110 0.710 5.350 0.780 ;
        RECT  4.980 0.200 5.310 0.280 ;
        RECT  5.070 0.380 5.150 0.640 ;
        RECT  5.010 0.710 5.110 1.070 ;
        RECT  4.790 0.380 5.070 0.450 ;
        RECT  4.730 0.710 5.010 0.780 ;
        RECT  4.690 0.190 4.790 0.450 ;
        RECT  4.690 0.850 4.790 1.070 ;
        RECT  4.650 0.520 4.730 0.780 ;
        RECT  4.450 0.380 4.690 0.450 ;
        RECT  4.490 0.850 4.690 0.920 ;
        RECT  4.410 0.710 4.650 0.780 ;
        RECT  4.280 0.200 4.610 0.280 ;
        RECT  4.370 0.380 4.450 0.640 ;
        RECT  4.310 0.710 4.410 1.070 ;
        RECT  4.090 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.310 0.780 ;
        RECT  3.990 0.190 4.090 0.450 ;
        RECT  3.990 0.850 4.090 1.070 ;
        RECT  3.950 0.520 4.030 0.780 ;
        RECT  3.750 0.380 3.990 0.450 ;
        RECT  3.790 0.850 3.990 0.920 ;
        RECT  3.710 0.710 3.950 0.780 ;
        RECT  3.580 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.750 0.640 ;
        RECT  3.610 0.710 3.710 1.070 ;
        RECT  3.390 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.610 0.780 ;
        RECT  3.290 0.190 3.390 0.450 ;
        RECT  3.290 0.850 3.390 1.070 ;
        RECT  3.250 0.520 3.330 0.780 ;
        RECT  3.050 0.380 3.290 0.450 ;
        RECT  3.090 0.850 3.290 0.920 ;
        RECT  3.010 0.710 3.250 0.780 ;
        RECT  2.880 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.050 0.640 ;
        RECT  2.910 0.710 3.010 1.070 ;
        RECT  2.690 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.910 0.780 ;
        RECT  2.590 0.190 2.690 0.450 ;
        RECT  2.590 0.850 2.690 1.070 ;
        RECT  2.550 0.520 2.630 0.780 ;
        RECT  2.350 0.380 2.590 0.450 ;
        RECT  2.390 0.850 2.590 0.920 ;
        RECT  2.310 0.710 2.550 0.780 ;
        RECT  2.180 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.350 0.640 ;
        RECT  2.210 0.710 2.310 1.070 ;
        RECT  1.990 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.210 0.780 ;
        RECT  1.890 0.190 1.990 0.450 ;
        RECT  1.890 0.850 1.990 1.070 ;
        RECT  1.850 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.690 0.850 1.890 0.920 ;
        RECT  1.610 0.710 1.850 0.780 ;
        RECT  1.480 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.190 0.850 1.290 1.070 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.990 0.850 1.190 0.920 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.780 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.490 0.850 0.590 1.070 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.290 0.850 0.490 0.920 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.080 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GFILL10BWP

MACRO GFILL2BWP
    CLASS CORE ;
    FOREIGN GFILL2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 1.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.190 1.300 0.450 ;
        RECT  1.190 0.850 1.300 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.990 0.850 1.190 0.920 ;
        RECT  0.910 0.710 1.145 0.780 ;
        RECT  0.780 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.490 0.850 0.590 1.070 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.290 0.850 0.490 0.920 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.080 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GFILL2BWP

MACRO GFILL3BWP
    CLASS CORE ;
    FOREIGN GFILL3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.890 0.190 2.000 0.450 ;
        RECT  1.890 0.850 2.000 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.690 0.850 1.890 0.920 ;
        RECT  1.610 0.710 1.845 0.780 ;
        RECT  1.480 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.190 0.850 1.290 1.070 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.990 0.850 1.190 0.920 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.780 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.490 0.850 0.590 1.070 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.290 0.850 0.490 0.920 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.080 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GFILL3BWP

MACRO GFILL4BWP
    CLASS CORE ;
    FOREIGN GFILL4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.800 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.590 0.190 2.700 0.450 ;
        RECT  2.590 0.850 2.700 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.350 0.380 2.590 0.450 ;
        RECT  2.390 0.850 2.590 0.920 ;
        RECT  2.310 0.710 2.545 0.780 ;
        RECT  2.180 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.350 0.640 ;
        RECT  2.210 0.710 2.310 1.070 ;
        RECT  1.990 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.210 0.780 ;
        RECT  1.890 0.190 1.990 0.450 ;
        RECT  1.890 0.850 1.990 1.070 ;
        RECT  1.850 0.520 1.930 0.780 ;
        RECT  1.650 0.380 1.890 0.450 ;
        RECT  1.690 0.850 1.890 0.920 ;
        RECT  1.610 0.710 1.850 0.780 ;
        RECT  1.480 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.650 0.640 ;
        RECT  1.510 0.710 1.610 1.070 ;
        RECT  1.290 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.190 0.190 1.290 0.450 ;
        RECT  1.190 0.850 1.290 1.070 ;
        RECT  1.150 0.520 1.230 0.780 ;
        RECT  0.950 0.380 1.190 0.450 ;
        RECT  0.990 0.850 1.190 0.920 ;
        RECT  0.910 0.710 1.150 0.780 ;
        RECT  0.780 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.950 0.640 ;
        RECT  0.810 0.710 0.910 1.070 ;
        RECT  0.590 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.810 0.780 ;
        RECT  0.490 0.190 0.590 0.450 ;
        RECT  0.490 0.850 0.590 1.070 ;
        RECT  0.450 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.290 0.850 0.490 0.920 ;
        RECT  0.210 0.710 0.450 0.780 ;
        RECT  0.080 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GFILL4BWP

MACRO GFILLBWP
    CLASS CORE ;
    FOREIGN GFILLBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.700 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.700 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.490 0.190 0.600 0.450 ;
        RECT  0.490 0.850 0.600 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.490 0.450 ;
        RECT  0.290 0.850 0.490 0.920 ;
        RECT  0.210 0.710 0.445 0.780 ;
        RECT  0.080 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.100 0.710 0.210 1.070 ;
    END
END GFILLBWP

MACRO GINVD1BWP
    CLASS CORE ;
    FOREIGN GINVD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.210 0.290 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.530 0.765 ;
        RECT  0.265 0.675 0.435 0.765 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.700 0.115 ;
        RECT  0.500 -0.115 0.580 0.320 ;
        RECT  0.390 -0.115 0.500 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.700 1.375 ;
        RECT  0.500 0.850 0.580 1.375 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.000 1.145 0.500 1.375 ;
        END
    END VDD
END GINVD1BWP

MACRO GINVD2BWP
    CLASS CORE ;
    FOREIGN GINVD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.315 0.775 0.385 0.955 ;
        RECT  0.105 0.775 0.315 0.845 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.845 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.525 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.700 0.115 ;
        RECT  0.500 -0.115 0.580 0.320 ;
        RECT  0.220 -0.115 0.500 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.700 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.220 1.145 0.500 1.375 ;
        RECT  0.100 0.970 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
END GINVD2BWP

MACRO GINVD3BWP
    CLASS CORE ;
    FOREIGN GINVD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.190 0.910 0.425 ;
        RECT  0.810 0.805 0.910 1.070 ;
        RECT  0.400 0.355 0.810 0.425 ;
        RECT  0.400 0.805 0.810 0.875 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.300 0.805 0.400 0.955 ;
        RECT  0.105 0.355 0.300 0.425 ;
        RECT  0.105 0.805 0.300 0.875 ;
        RECT  0.035 0.355 0.105 0.875 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 1.295 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.320 ;
        RECT  1.090 -0.115 1.200 0.115 ;
        RECT  1.010 -0.115 1.090 0.320 ;
        RECT  0.600 -0.115 1.010 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 1.145 1.400 1.375 ;
        RECT  1.205 0.850 1.275 1.375 ;
        RECT  0.990 0.850 1.205 0.920 ;
        RECT  0.580 1.145 1.205 1.375 ;
        RECT  0.500 0.960 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.960 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
END GINVD3BWP

MACRO GINVD4BWP
    CLASS CORE ;
    FOREIGN GINVD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2304 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  1.000 0.805 1.085 0.955 ;
        RECT  0.400 0.355 1.000 0.425 ;
        RECT  0.400 0.805 1.000 0.875 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.300 0.805 0.400 0.955 ;
        RECT  0.105 0.355 0.300 0.425 ;
        RECT  0.105 0.805 0.300 0.875 ;
        RECT  0.035 0.355 0.105 0.875 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 1.225 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.320 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.960 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.960 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.960 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
END GINVD4BWP

MACRO GINVD8BWP
    CLASS CORE ;
    FOREIGN GINVD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4608 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.400 0.190 2.500 0.425 ;
        RECT  2.400 0.805 2.485 0.955 ;
        RECT  1.800 0.355 2.400 0.425 ;
        RECT  1.800 0.805 2.400 0.875 ;
        RECT  1.700 0.190 1.800 0.425 ;
        RECT  1.700 0.805 1.800 0.955 ;
        RECT  1.100 0.355 1.700 0.425 ;
        RECT  1.100 0.805 1.700 0.875 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  1.000 0.805 1.100 0.955 ;
        RECT  0.400 0.355 1.000 0.425 ;
        RECT  0.400 0.805 1.000 0.875 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.300 0.805 0.400 0.955 ;
        RECT  0.105 0.355 0.300 0.425 ;
        RECT  0.105 0.805 0.300 0.875 ;
        RECT  0.035 0.355 0.105 0.875 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 2.625 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 -0.115 2.800 0.115 ;
        RECT  2.600 -0.115 2.680 0.320 ;
        RECT  2.320 -0.115 2.600 0.115 ;
        RECT  2.200 -0.115 2.320 0.280 ;
        RECT  2.000 -0.115 2.200 0.115 ;
        RECT  1.880 -0.115 2.000 0.280 ;
        RECT  1.620 -0.115 1.880 0.115 ;
        RECT  1.500 -0.115 1.620 0.280 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.280 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.280 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 1.145 2.800 1.375 ;
        RECT  2.600 0.940 2.680 1.375 ;
        RECT  2.300 1.145 2.600 1.375 ;
        RECT  2.220 0.960 2.300 1.375 ;
        RECT  1.980 1.145 2.220 1.375 ;
        RECT  1.900 0.960 1.980 1.375 ;
        RECT  1.600 1.145 1.900 1.375 ;
        RECT  1.520 0.960 1.600 1.375 ;
        RECT  1.280 1.145 1.520 1.375 ;
        RECT  1.200 0.960 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.960 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.960 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.960 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
END GINVD8BWP

MACRO GMUX2D1BWP
    CLASS CORE ;
    FOREIGN GMUX2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.215 0.290 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.815 0.665 1.975 0.735 ;
        LAYER M1 ;
        RECT  1.835 0.495 1.925 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.665 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.670 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.145 2.100 1.375 ;
        RECT  1.740 0.835 1.810 1.375 ;
        RECT  1.700 0.835 1.740 0.935 ;
        RECT  0.410 1.145 1.740 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.995 0.355 2.065 1.070 ;
        RECT  1.890 0.190 1.995 0.425 ;
        RECT  1.890 0.970 1.995 1.070 ;
        RECT  1.225 0.355 1.890 0.425 ;
        RECT  1.180 0.200 1.620 0.275 ;
        RECT  1.510 0.775 1.610 1.075 ;
        RECT  1.190 0.775 1.290 1.075 ;
        RECT  1.155 0.355 1.225 0.660 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.425 ;
        RECT  0.335 0.355 1.000 0.425 ;
        RECT  0.855 0.495 0.945 0.765 ;
        RECT  0.480 0.200 0.920 0.275 ;
        RECT  0.810 0.845 0.910 1.075 ;
        RECT  0.490 0.775 0.590 1.070 ;
        RECT  0.265 0.355 0.335 0.640 ;
        RECT  0.175 0.520 0.265 0.640 ;
        LAYER VIA1 ;
        RECT  1.855 0.665 1.925 0.735 ;
        RECT  1.530 0.945 1.600 1.015 ;
        RECT  1.205 0.805 1.275 0.875 ;
        RECT  0.865 0.665 0.935 0.735 ;
        RECT  0.825 0.945 0.895 1.015 ;
        RECT  0.505 0.805 0.575 0.875 ;
        LAYER M2 ;
        RECT  0.775 0.945 1.650 1.015 ;
        RECT  0.455 0.805 1.325 0.875 ;
    END
END GMUX2D1BWP

MACRO GMUX2D2BWP
    CLASS CORE ;
    FOREIGN GMUX2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 0.420 0.920 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.665 2.675 0.735 ;
        LAYER M1 ;
        RECT  2.535 0.495 2.625 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.250 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.370 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.600 -0.115 0.990 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.280 1.145 2.440 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.220 1.145 0.500 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.695 0.355 2.765 1.070 ;
        RECT  2.590 0.190 2.695 0.425 ;
        RECT  2.590 0.970 2.695 1.070 ;
        RECT  1.925 0.355 2.590 0.425 ;
        RECT  1.880 0.200 2.320 0.275 ;
        RECT  2.210 0.775 2.310 1.075 ;
        RECT  1.890 0.775 1.990 1.075 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.560 0.495 1.645 0.765 ;
        RECT  1.250 0.200 1.620 0.275 ;
        RECT  1.510 0.845 1.610 1.075 ;
        RECT  1.180 0.200 1.250 0.415 ;
        RECT  0.910 0.345 1.180 0.415 ;
        RECT  1.000 0.775 1.100 1.045 ;
        RECT  0.810 0.190 0.910 0.415 ;
        RECT  0.485 0.355 0.555 0.640 ;
        RECT  0.175 0.495 0.485 0.640 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.230 0.945 2.300 1.015 ;
        RECT  1.905 0.805 1.975 0.875 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.015 0.805 1.085 0.875 ;
        RECT  0.485 0.385 0.555 0.455 ;
        LAYER M2 ;
        RECT  1.475 0.945 2.350 1.015 ;
        RECT  0.965 0.805 2.025 0.875 ;
        RECT  0.435 0.385 1.835 0.455 ;
    END
END GMUX2D2BWP

MACRO GMUX2ND1BWP
    CLASS CORE ;
    FOREIGN GMUX2ND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.210 0.290 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.665 2.675 0.735 ;
        LAYER M1 ;
        RECT  2.535 0.495 2.625 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.250 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.370 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.390 -0.115 0.990 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.280 1.145 2.440 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.410 1.145 0.820 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.695 0.355 2.765 1.070 ;
        RECT  2.590 0.190 2.695 0.425 ;
        RECT  2.590 0.970 2.695 1.070 ;
        RECT  1.925 0.355 2.590 0.425 ;
        RECT  1.880 0.200 2.320 0.275 ;
        RECT  2.210 0.775 2.310 1.075 ;
        RECT  1.890 0.775 1.990 1.075 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.560 0.495 1.645 0.765 ;
        RECT  1.250 0.200 1.620 0.275 ;
        RECT  1.510 0.845 1.610 1.075 ;
        RECT  1.180 0.200 1.250 0.415 ;
        RECT  0.910 0.345 1.180 0.415 ;
        RECT  1.000 0.775 1.100 1.045 ;
        RECT  0.810 0.190 0.910 0.415 ;
        RECT  0.635 0.355 0.705 0.615 ;
        RECT  0.430 0.545 0.635 0.615 ;
        RECT  0.555 0.185 0.595 0.290 ;
        RECT  0.560 0.970 0.595 1.070 ;
        RECT  0.490 0.695 0.560 1.070 ;
        RECT  0.485 0.185 0.555 0.440 ;
        RECT  0.245 0.695 0.490 0.765 ;
        RECT  0.245 0.370 0.485 0.440 ;
        RECT  0.175 0.370 0.245 0.765 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.230 0.945 2.300 1.015 ;
        RECT  1.905 0.805 1.975 0.875 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.015 0.805 1.085 0.875 ;
        RECT  0.635 0.385 0.705 0.455 ;
        LAYER M2 ;
        RECT  1.475 0.945 2.350 1.015 ;
        RECT  0.965 0.805 2.025 0.875 ;
        RECT  0.585 0.385 1.835 0.455 ;
    END
END GMUX2ND1BWP

MACRO GMUX2ND2BWP
    CLASS CORE ;
    FOREIGN GMUX2ND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 0.420 0.920 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.300 0.190 0.385 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.515 0.665 2.675 0.735 ;
        LAYER M1 ;
        RECT  2.535 0.495 2.625 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.365 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.370 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.580 -0.115 0.990 0.115 ;
        RECT  0.500 -0.115 0.580 0.300 ;
        RECT  0.220 -0.115 0.500 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.110 1.145 2.440 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.580 1.145 0.990 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.220 1.145 0.500 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.695 0.355 2.765 1.070 ;
        RECT  2.590 0.190 2.695 0.425 ;
        RECT  2.590 0.970 2.695 1.070 ;
        RECT  1.925 0.355 2.590 0.425 ;
        RECT  1.880 0.200 2.320 0.275 ;
        RECT  2.210 0.775 2.310 1.075 ;
        RECT  1.890 0.775 1.990 1.075 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.425 ;
        RECT  1.035 0.355 1.700 0.425 ;
        RECT  1.555 0.495 1.645 0.765 ;
        RECT  1.180 0.200 1.620 0.275 ;
        RECT  1.510 0.845 1.610 1.075 ;
        RECT  1.190 0.775 1.290 1.070 ;
        RECT  0.965 0.355 1.035 0.615 ;
        RECT  0.830 0.545 0.965 0.615 ;
        RECT  0.875 0.185 0.915 0.290 ;
        RECT  0.875 0.970 0.910 1.070 ;
        RECT  0.805 0.185 0.875 0.445 ;
        RECT  0.805 0.695 0.875 1.070 ;
        RECT  0.525 0.375 0.805 0.445 ;
        RECT  0.525 0.695 0.805 0.765 ;
        RECT  0.455 0.375 0.525 0.765 ;
        RECT  0.245 0.695 0.455 0.765 ;
        RECT  0.175 0.500 0.245 0.765 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.230 0.945 2.300 1.015 ;
        RECT  1.905 0.805 1.975 0.875 ;
        RECT  1.565 0.665 1.635 0.735 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.205 0.805 1.275 0.875 ;
        LAYER M2 ;
        RECT  1.475 0.945 2.350 1.015 ;
        RECT  1.155 0.805 2.025 0.875 ;
    END
END GMUX2ND2BWP

MACRO GND2D1BWP
    CLASS CORE ;
    FOREIGN GND2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1183 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.190 0.665 0.920 ;
        RECT  0.490 0.190 0.595 0.290 ;
        RECT  0.280 0.850 0.595 0.920 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.220 -0.115 0.700 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.700 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.200 1.145 0.480 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.190 0.400 0.410 ;
    END
END GND2D1BWP

MACRO GND2D2BWP
    CLASS CORE ;
    FOREIGN GND2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2366 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.850 1.130 0.920 ;
        RECT  0.805 0.205 0.920 0.275 ;
        RECT  0.735 0.205 0.805 0.920 ;
        RECT  0.480 0.205 0.735 0.275 ;
        RECT  0.270 0.850 0.735 0.920 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.125 0.385 1.275 0.455 ;
        LAYER M1 ;
        RECT  0.175 0.355 0.245 0.675 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.405 0.665 0.995 0.735 ;
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.220 -0.115 1.180 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.200 1.145 0.480 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.355 1.230 0.675 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.605 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.455 0.445 0.530 0.765 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.605 ;
        RECT  0.300 0.190 0.315 0.290 ;
        LAYER VIA1 ;
        RECT  1.155 0.385 1.225 0.455 ;
        RECT  0.875 0.665 0.945 0.735 ;
        RECT  0.455 0.665 0.525 0.735 ;
        RECT  0.175 0.385 0.245 0.455 ;
    END
END GND2D2BWP

MACRO GND2D3BWP
    CLASS CORE ;
    FOREIGN GND2D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3549 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.060 0.245 0.630 0.315 ;
        LAYER M1 ;
        RECT  0.105 0.845 1.820 0.915 ;
        RECT  0.105 0.190 0.220 0.315 ;
        RECT  0.035 0.190 0.105 0.915 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.645 0.695 1.855 0.765 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.225 0.695 1.575 0.765 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.525 0.695 0.875 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.245 0.695 0.455 0.765 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 -0.115 2.100 0.115 ;
        RECT  1.900 -0.115 1.980 0.320 ;
        RECT  1.620 -0.115 1.900 0.115 ;
        RECT  1.500 -0.115 1.620 0.275 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.000 -0.115 1.180 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.145 2.100 1.375 ;
        RECT  1.880 0.985 2.000 1.375 ;
        RECT  1.620 1.145 1.880 1.375 ;
        RECT  1.500 0.985 1.620 1.375 ;
        RECT  1.300 1.145 1.500 1.375 ;
        RECT  1.180 0.985 1.300 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.220 1.145 0.480 1.375 ;
        RECT  0.100 0.985 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.505 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.505 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.480 0.200 0.920 0.315 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.505 ;
        RECT  0.300 0.190 0.315 0.290 ;
        LAYER VIA1 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.510 0.245 0.580 0.315 ;
        RECT  0.315 0.385 0.385 0.455 ;
        RECT  0.110 0.245 0.180 0.315 ;
        LAYER M2 ;
        RECT  0.265 0.385 1.835 0.455 ;
    END
END GND2D3BWP

MACRO GND2D4BWP
    CLASS CORE ;
    FOREIGN GND2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4732 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.060 0.245 0.630 0.315 ;
        LAYER M1 ;
        RECT  1.365 0.845 2.520 0.915 ;
        RECT  1.295 0.205 1.365 0.915 ;
        RECT  1.180 0.205 1.295 0.275 ;
        RECT  0.105 0.845 1.295 0.915 ;
        RECT  0.105 0.190 0.220 0.315 ;
        RECT  0.035 0.190 0.105 0.915 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.625 0.765 ;
        RECT  2.345 0.695 2.555 0.765 ;
        RECT  2.275 0.495 2.345 0.765 ;
        RECT  1.925 0.695 2.275 0.765 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.645 0.695 1.855 0.765 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  0.945 0.695 1.155 0.765 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.525 0.695 0.875 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.245 0.695 0.455 0.765 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.680 -0.115 2.800 0.115 ;
        RECT  2.600 -0.115 2.680 0.320 ;
        RECT  2.320 -0.115 2.600 0.115 ;
        RECT  2.200 -0.115 2.320 0.275 ;
        RECT  2.000 -0.115 2.200 0.115 ;
        RECT  1.880 -0.115 2.000 0.275 ;
        RECT  1.620 -0.115 1.880 0.115 ;
        RECT  1.500 -0.115 1.620 0.275 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.145 2.800 1.375 ;
        RECT  2.580 0.985 2.700 1.375 ;
        RECT  2.320 1.145 2.580 1.375 ;
        RECT  2.200 0.985 2.320 1.375 ;
        RECT  2.000 1.145 2.200 1.375 ;
        RECT  1.880 0.985 2.000 1.375 ;
        RECT  1.620 1.145 1.880 1.375 ;
        RECT  1.500 0.985 1.620 1.375 ;
        RECT  1.300 1.145 1.500 1.375 ;
        RECT  1.180 0.985 1.300 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.220 1.145 0.480 1.375 ;
        RECT  0.100 0.985 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.190 2.500 0.290 ;
        RECT  2.415 0.190 2.485 0.505 ;
        RECT  2.400 0.190 2.415 0.290 ;
        RECT  1.015 0.190 1.085 0.505 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.480 0.200 0.920 0.315 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.505 ;
        RECT  0.300 0.190 0.315 0.290 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.505 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.085 0.190 1.100 0.290 ;
        LAYER VIA1 ;
        RECT  2.415 0.385 2.485 0.455 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.510 0.245 0.580 0.315 ;
        RECT  0.315 0.385 0.385 0.455 ;
        RECT  0.110 0.245 0.180 0.315 ;
        LAYER M2 ;
        RECT  0.265 0.385 2.535 0.455 ;
    END
END GND2D4BWP

MACRO GND3D1BWP
    CLASS CORE ;
    FOREIGN GND3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1839 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 1.110 0.920 ;
        RECT  0.105 0.190 0.210 0.290 ;
        RECT  0.035 0.190 0.105 0.920 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.495 0.665 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.495 1.235 0.765 ;
        RECT  0.960 0.695 1.145 0.765 ;
        RECT  0.865 0.495 0.960 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.320 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.220 1.145 0.480 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.590 0.345 1.000 0.415 ;
        RECT  0.490 0.190 0.590 0.415 ;
        RECT  0.300 0.190 0.400 0.410 ;
    END
END GND3D1BWP

MACRO GND3D2BWP
    CLASS CORE ;
    FOREIGN GND3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.3022 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.075 0.245 2.040 0.315 ;
        LAYER M1 ;
        RECT  1.995 0.190 2.065 0.920 ;
        RECT  1.890 0.190 1.995 0.345 ;
        RECT  0.270 0.850 1.995 0.920 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.225 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.645 0.640 ;
        RECT  0.525 0.355 1.575 0.425 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.780 ;
        RECT  0.245 0.710 1.855 0.780 ;
        RECT  0.175 0.495 0.245 0.780 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 2.100 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.000 -0.115 0.990 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.145 2.100 1.375 ;
        RECT  1.880 0.990 2.000 1.375 ;
        RECT  1.620 1.145 1.880 1.375 ;
        RECT  1.500 0.990 1.620 1.375 ;
        RECT  1.300 1.145 1.500 1.375 ;
        RECT  1.180 0.990 1.300 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.220 1.145 0.480 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.190 1.810 0.410 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.180 0.200 1.620 0.275 ;
        RECT  0.480 0.200 0.920 0.275 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.290 0.190 0.385 0.410 ;
        RECT  0.100 0.190 0.210 0.410 ;
        LAYER VIA1 ;
        RECT  1.920 0.245 1.990 0.315 ;
        RECT  0.125 0.245 0.195 0.315 ;
    END
END GND3D2BWP

MACRO GNR2D1BWP
    CLASS CORE ;
    FOREIGN GNR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1193 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.490 0.970 0.595 1.070 ;
        RECT  0.300 0.190 0.400 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 -0.115 0.700 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.145 0.700 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.850 0.410 1.070 ;
    END
END GNR2D1BWP

MACRO GNR2D2BWP
    CLASS CORE ;
    FOREIGN GNR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2386 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.365 1.070 ;
        RECT  1.100 0.345 1.295 0.415 ;
        RECT  1.190 0.970 1.295 1.070 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.400 0.345 1.000 0.415 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.345 0.105 1.070 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.780 ;
        RECT  0.245 0.710 1.155 0.780 ;
        RECT  0.175 0.495 0.245 0.780 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.495 0.970 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.145 1.400 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.600 1.145 0.800 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.000 1.145 0.480 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.850 1.110 1.060 ;
        RECT  0.290 0.850 0.410 1.060 ;
    END
END GNR2D2BWP

MACRO GNR3D1BWP
    CLASS CORE ;
    FOREIGN GNR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1689 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  0.400 0.355 1.000 0.425 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.105 0.355 0.300 0.425 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.355 0.105 1.070 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 1.250 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.320 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.400 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.000 1.145 0.800 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.850 1.120 0.920 ;
        RECT  0.640 0.850 0.720 1.055 ;
        RECT  0.480 0.985 0.640 1.055 ;
        RECT  0.300 0.835 0.400 1.055 ;
    END
END GNR3D1BWP

MACRO GNR3D2BWP
    CLASS CORE ;
    FOREIGN GNR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2882 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.190 1.800 0.415 ;
        RECT  1.100 0.345 1.700 0.415 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.400 0.345 1.000 0.415 ;
        RECT  0.105 0.990 0.600 1.060 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 1.060 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.930 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 1.230 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.530 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.100 0.115 ;
        RECT  1.890 -0.115 2.000 0.290 ;
        RECT  1.620 -0.115 1.890 0.115 ;
        RECT  1.500 -0.115 1.620 0.275 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.145 2.100 1.375 ;
        RECT  1.900 0.940 1.980 1.375 ;
        RECT  1.620 1.145 1.900 1.375 ;
        RECT  1.500 0.990 1.620 1.375 ;
        RECT  0.000 1.145 1.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.970 0.850 1.810 0.920 ;
        RECT  0.805 0.990 1.320 1.060 ;
        RECT  0.735 0.850 0.805 1.060 ;
        RECT  0.270 0.850 0.735 0.920 ;
    END
END GNR3D2BWP

MACRO GOAI21D1BWP
    CLASS CORE ;
    FOREIGN GOAI21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.2407 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.075 0.245 0.715 0.315 ;
        LAYER M1 ;
        RECT  0.665 0.850 1.130 0.920 ;
        RECT  0.595 0.190 0.665 1.055 ;
        RECT  0.490 0.190 0.595 0.290 ;
        RECT  0.480 0.985 0.595 1.055 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.230 0.765 ;
        RECT  0.945 0.685 1.155 0.765 ;
        RECT  0.855 0.495 0.945 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.445 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.280 0.320 ;
        RECT  0.900 -0.115 1.200 0.115 ;
        RECT  0.820 -0.115 0.900 0.320 ;
        RECT  0.000 -0.115 0.820 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 1.145 1.400 1.375 ;
        RECT  1.205 0.940 1.275 1.375 ;
        RECT  0.920 1.145 1.205 1.375 ;
        RECT  0.800 0.990 0.920 1.375 ;
        RECT  0.200 1.145 0.800 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.485 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.290 0.850 0.410 1.060 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.485 ;
        RECT  0.300 0.190 0.315 0.290 ;
        RECT  0.100 0.190 0.210 0.415 ;
        LAYER VIA1 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.595 0.245 0.665 0.315 ;
        RECT  0.315 0.385 0.385 0.455 ;
        RECT  0.125 0.245 0.195 0.315 ;
        LAYER M2 ;
        RECT  0.265 0.385 1.135 0.455 ;
    END
END GOAI21D1BWP

MACRO GOAI21D2BWP
    CLASS CORE ;
    FOREIGN GOAI21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.4158 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.620 0.245 2.040 0.315 ;
        LAYER M1 ;
        RECT  1.995 0.190 2.065 1.070 ;
        RECT  1.890 0.190 1.995 0.345 ;
        RECT  1.890 0.970 1.995 1.070 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        RECT  0.245 0.695 0.455 0.765 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.645 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.500 1.925 0.780 ;
        RECT  0.945 0.710 1.855 0.780 ;
        RECT  0.875 0.495 0.945 0.780 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 2.100 0.115 ;
        RECT  0.500 -0.115 0.580 0.320 ;
        RECT  0.210 -0.115 0.500 0.115 ;
        RECT  0.100 -0.115 0.210 0.290 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.145 2.100 1.375 ;
        RECT  1.520 0.940 1.600 1.375 ;
        RECT  1.280 1.145 1.520 1.375 ;
        RECT  1.200 0.940 1.280 1.375 ;
        RECT  0.600 1.145 1.200 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.200 1.145 0.480 1.375 ;
        RECT  0.120 0.935 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.850 1.810 1.060 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.485 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.180 0.205 1.620 0.315 ;
        RECT  0.990 0.850 1.110 1.060 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.485 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.740 0.190 0.910 0.290 ;
        RECT  0.810 0.850 0.910 1.070 ;
        RECT  0.740 0.850 0.810 0.920 ;
        RECT  0.670 0.190 0.740 0.920 ;
        RECT  0.270 0.850 0.670 0.920 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.485 ;
        RECT  0.300 0.190 0.315 0.290 ;
        LAYER VIA1 ;
        RECT  1.920 0.245 1.990 0.315 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.365 0.245 1.435 0.315 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.670 0.245 0.740 0.315 ;
        RECT  0.315 0.385 0.385 0.455 ;
        LAYER M2 ;
        RECT  0.265 0.385 1.835 0.455 ;
    END
END GOAI21D2BWP

MACRO GOR2D1BWP
    CLASS CORE ;
    FOREIGN GOR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.190 1.365 1.070 ;
        RECT  1.190 0.190 1.295 0.290 ;
        RECT  1.190 0.970 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.895 -0.115 1.010 0.115 ;
        RECT  0.825 -0.115 0.895 0.300 ;
        RECT  0.600 -0.115 0.825 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.145 1.400 1.375 ;
        RECT  0.895 0.850 1.130 0.920 ;
        RECT  0.825 0.850 0.895 1.375 ;
        RECT  0.200 1.145 0.825 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.500 1.225 0.780 ;
        RECT  0.945 0.710 1.155 0.780 ;
        RECT  0.875 0.500 0.945 0.780 ;
        RECT  0.665 0.710 0.875 0.780 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.490 0.970 0.595 1.070 ;
        RECT  0.290 0.845 0.410 1.055 ;
        RECT  0.300 0.190 0.400 0.415 ;
    END
END GOR2D1BWP

MACRO GOR2D2BWP
    CLASS CORE ;
    FOREIGN GOR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.365 0.920 ;
        RECT  1.100 0.345 1.295 0.415 ;
        RECT  0.980 0.850 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.415 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.180 -0.115 1.300 0.275 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.600 -0.115 0.800 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.400 1.375 ;
        RECT  1.180 0.990 1.300 1.375 ;
        RECT  0.900 1.145 1.180 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.200 1.145 0.820 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.145 0.500 1.225 0.780 ;
        RECT  0.945 0.710 1.145 0.780 ;
        RECT  0.875 0.500 0.945 0.780 ;
        RECT  0.665 0.710 0.875 0.780 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.490 0.970 0.595 1.070 ;
        RECT  0.290 0.845 0.410 1.055 ;
        RECT  0.300 0.190 0.400 0.415 ;
    END
END GOR2D2BWP

MACRO GSDFCNQD1BWP
    CLASS CORE ;
    FOREIGN GSDFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN SI
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.405 0.545 0.970 0.615 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.195 0.205 6.265 1.055 ;
        RECT  6.080 0.205 6.195 0.275 ;
        RECT  6.080 0.985 6.195 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.645 0.685 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.805 0.385 2.675 0.455 ;
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.640 ;
        RECT  1.715 0.495 1.855 0.640 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  3.795 0.665 5.475 0.735 ;
        RECT  3.725 0.525 3.795 0.735 ;
        RECT  3.340 0.525 3.725 0.595 ;
        LAYER M1 ;
        RECT  5.355 0.355 5.425 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.010 -0.115 6.300 0.115 ;
        RECT  5.890 -0.115 6.010 0.270 ;
        RECT  5.100 -0.115 5.890 0.115 ;
        RECT  5.015 -0.115 5.100 0.315 ;
        RECT  3.895 -0.115 5.015 0.115 ;
        RECT  3.820 -0.115 3.895 0.315 ;
        RECT  3.400 -0.115 3.820 0.115 ;
        RECT  3.310 -0.115 3.400 0.310 ;
        RECT  1.810 -0.115 3.310 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.390 -0.115 1.690 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.010 1.145 6.300 1.375 ;
        RECT  5.920 0.805 6.010 1.375 ;
        RECT  5.290 1.145 5.920 1.375 ;
        RECT  5.215 0.820 5.290 1.375 ;
        RECT  3.910 1.145 5.215 1.375 ;
        RECT  3.790 0.850 3.910 1.375 ;
        RECT  3.210 1.145 3.790 1.375 ;
        RECT  3.090 0.850 3.210 1.375 ;
        RECT  1.810 1.145 3.090 1.375 ;
        RECT  1.690 0.850 1.810 1.375 ;
        RECT  0.410 1.145 1.690 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.845 0.520 6.125 0.640 ;
        RECT  5.775 0.520 5.845 0.905 ;
        RECT  5.705 0.205 5.820 0.275 ;
        RECT  5.705 0.985 5.820 1.055 ;
        RECT  5.635 0.205 5.705 1.055 ;
        RECT  5.495 0.205 5.565 1.055 ;
        RECT  5.380 0.205 5.495 0.275 ;
        RECT  5.380 0.985 5.495 1.055 ;
        RECT  5.285 0.195 5.310 0.290 ;
        RECT  5.180 0.195 5.285 0.475 ;
        RECT  4.935 0.545 5.220 0.615 ;
        RECT  5.010 0.770 5.110 1.070 ;
        RECT  4.915 0.385 5.055 0.455 ;
        RECT  4.865 0.545 4.935 0.780 ;
        RECT  4.845 0.200 4.915 0.455 ;
        RECT  4.585 0.710 4.865 0.780 ;
        RECT  4.675 0.200 4.845 0.280 ;
        RECT  4.690 0.850 4.790 1.070 ;
        RECT  4.655 0.385 4.745 0.640 ;
        RECT  4.585 0.185 4.605 0.315 ;
        RECT  4.515 0.185 4.585 0.965 ;
        RECT  4.375 0.185 4.445 0.370 ;
        RECT  4.375 0.520 4.445 0.905 ;
        RECT  4.305 0.985 4.415 1.055 ;
        RECT  4.235 0.185 4.375 0.275 ;
        RECT  4.235 0.355 4.305 1.055 ;
        RECT  4.095 0.205 4.165 1.055 ;
        RECT  3.980 0.205 4.095 0.275 ;
        RECT  3.980 0.985 4.095 1.055 ;
        RECT  3.955 0.485 4.025 0.765 ;
        RECT  2.625 0.695 3.955 0.765 ;
        RECT  3.745 0.545 3.795 0.615 ;
        RECT  3.675 0.345 3.745 0.615 ;
        RECT  3.560 0.190 3.725 0.270 ;
        RECT  3.610 0.850 3.710 1.070 ;
        RECT  3.650 0.545 3.675 0.615 ;
        RECT  3.200 0.515 3.570 0.615 ;
        RECT  3.490 0.190 3.560 0.365 ;
        RECT  3.290 0.850 3.390 1.070 ;
        RECT  3.090 0.185 3.210 0.395 ;
        RECT  2.905 0.515 3.095 0.615 ;
        RECT  2.580 0.205 3.020 0.275 ;
        RECT  2.910 0.850 3.010 1.070 ;
        RECT  2.835 0.355 2.905 0.615 ;
        RECT  2.590 0.850 2.690 1.070 ;
        RECT  2.555 0.355 2.625 0.765 ;
        RECT  2.485 0.190 2.500 0.290 ;
        RECT  2.415 0.190 2.485 0.965 ;
        RECT  2.400 0.190 2.415 0.290 ;
        RECT  2.090 0.520 2.340 0.640 ;
        RECT  2.210 0.190 2.310 0.410 ;
        RECT  2.210 0.775 2.310 1.070 ;
        RECT  2.020 0.205 2.090 1.055 ;
        RECT  1.880 0.205 2.020 0.275 ;
        RECT  1.880 0.985 2.020 1.055 ;
        RECT  1.505 0.205 1.620 0.275 ;
        RECT  1.505 0.985 1.620 1.055 ;
        RECT  1.435 0.205 1.505 1.055 ;
        RECT  1.180 0.205 1.435 0.275 ;
        RECT  1.190 0.850 1.290 1.070 ;
        RECT  1.060 0.495 1.270 0.625 ;
        RECT  1.000 0.775 1.120 1.070 ;
        RECT  1.000 0.190 1.100 0.410 ;
        RECT  0.760 0.190 0.910 0.410 ;
        RECT  0.800 0.685 0.910 1.070 ;
        RECT  0.475 0.190 0.605 0.455 ;
        RECT  0.490 0.775 0.590 1.070 ;
        RECT  0.100 0.190 0.210 0.425 ;
        RECT  0.100 0.850 0.210 1.070 ;
        LAYER VIA1 ;
        RECT  5.775 0.805 5.845 0.875 ;
        RECT  5.635 0.245 5.705 0.315 ;
        RECT  5.635 0.945 5.705 1.015 ;
        RECT  5.495 0.805 5.565 0.875 ;
        RECT  5.355 0.665 5.425 0.735 ;
        RECT  5.025 0.805 5.095 0.875 ;
        RECT  4.935 0.385 5.005 0.455 ;
        RECT  4.705 0.945 4.775 1.015 ;
        RECT  4.655 0.525 4.725 0.595 ;
        RECT  4.375 0.245 4.445 0.315 ;
        RECT  4.375 0.805 4.445 0.875 ;
        RECT  4.235 0.385 4.305 0.455 ;
        RECT  4.235 0.945 4.305 1.015 ;
        RECT  4.095 0.805 4.165 0.875 ;
        RECT  3.955 0.525 4.025 0.595 ;
        RECT  3.675 0.385 3.745 0.455 ;
        RECT  3.625 0.945 3.695 1.015 ;
        RECT  3.490 0.245 3.560 0.315 ;
        RECT  3.395 0.525 3.465 0.595 ;
        RECT  3.305 0.945 3.375 1.015 ;
        RECT  2.925 0.945 2.995 1.015 ;
        RECT  2.835 0.385 2.905 0.455 ;
        RECT  2.605 0.945 2.675 1.015 ;
        RECT  2.555 0.385 2.625 0.455 ;
        RECT  2.415 0.525 2.485 0.595 ;
        RECT  2.225 0.245 2.295 0.315 ;
        RECT  2.225 0.805 2.295 0.875 ;
        RECT  1.855 0.385 1.925 0.455 ;
        RECT  1.435 0.665 1.505 0.735 ;
        RECT  1.205 0.945 1.275 1.015 ;
        RECT  1.095 0.525 1.165 0.595 ;
        RECT  1.050 0.805 1.120 0.875 ;
        RECT  1.030 0.245 1.100 0.315 ;
        RECT  0.830 0.755 0.900 0.825 ;
        RECT  0.760 0.245 0.830 0.315 ;
        RECT  0.505 0.385 0.575 0.455 ;
        RECT  0.505 0.805 0.575 0.875 ;
        RECT  0.125 0.245 0.195 0.315 ;
        RECT  0.125 0.945 0.195 1.015 ;
        LAYER M2 ;
        RECT  4.975 0.805 5.895 0.875 ;
        RECT  4.325 0.245 5.755 0.315 ;
        RECT  4.655 0.945 5.755 1.015 ;
        RECT  4.025 0.385 5.055 0.455 ;
        RECT  3.905 0.525 4.775 0.595 ;
        RECT  4.045 0.805 4.495 0.875 ;
        RECT  3.575 0.945 4.355 1.015 ;
        RECT  3.955 0.245 4.025 0.455 ;
        RECT  3.045 0.245 3.955 0.315 ;
        RECT  3.185 0.385 3.795 0.455 ;
        RECT  2.905 0.945 3.425 1.015 ;
        RECT  3.115 0.385 3.185 0.595 ;
        RECT  2.365 0.525 3.115 0.595 ;
        RECT  2.975 0.245 3.045 0.455 ;
        RECT  2.785 0.385 2.975 0.455 ;
        RECT  2.835 0.805 2.905 1.015 ;
        RECT  2.175 0.805 2.835 0.875 ;
        RECT  2.065 0.945 2.725 1.015 ;
        RECT  0.980 0.245 2.345 0.315 ;
        RECT  1.995 0.805 2.065 1.015 ;
        RECT  1.000 0.805 1.995 0.875 ;
        RECT  0.900 0.665 1.555 0.735 ;
        RECT  0.075 0.945 1.325 1.015 ;
        RECT  0.665 0.525 1.215 0.595 ;
        RECT  0.830 0.665 0.900 0.875 ;
        RECT  0.075 0.245 0.880 0.315 ;
        RECT  0.595 0.385 0.665 0.875 ;
        RECT  0.455 0.385 0.595 0.455 ;
        RECT  0.455 0.805 0.595 0.875 ;
    END
END GSDFCNQD1BWP

MACRO GTIEHBWP
    CLASS CORE ;
    FOREIGN GTIEHBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.0656 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.775 0.390 1.065 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.700 0.115 ;
        RECT  0.500 -0.115 0.580 0.320 ;
        RECT  0.200 -0.115 0.500 0.115 ;
        RECT  0.120 -0.115 0.200 0.320 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.700 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.400 0.545 0.550 0.615 ;
        RECT  0.300 0.190 0.400 0.615 ;
        RECT  0.140 0.545 0.300 0.615 ;
    END
END GTIEHBWP

MACRO GTIELBWP
    CLASS CORE ;
    FOREIGN GTIELBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.0496 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.485 ;
        RECT  0.300 0.190 0.315 0.290 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 -0.115 0.700 0.115 ;
        RECT  0.500 -0.115 0.580 0.320 ;
        RECT  0.200 -0.115 0.500 0.115 ;
        RECT  0.120 -0.115 0.200 0.320 ;
        RECT  0.000 -0.115 0.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.700 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.200 1.145 0.500 1.375 ;
        RECT  0.120 0.940 0.200 1.375 ;
        RECT  0.000 1.145 0.120 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.455 0.500 0.530 0.765 ;
        RECT  0.390 0.695 0.455 0.765 ;
        RECT  0.310 0.695 0.390 0.965 ;
        RECT  0.245 0.695 0.310 0.765 ;
        RECT  0.170 0.500 0.245 0.765 ;
    END
END GTIELBWP

MACRO GXNR2D1BWP
    CLASS CORE ;
    FOREIGN GXNR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.215 0.290 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.815 0.665 1.975 0.735 ;
        LAYER M1 ;
        RECT  1.835 0.495 1.925 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.145 2.100 1.375 ;
        RECT  1.740 0.835 1.810 1.375 ;
        RECT  1.700 0.835 1.740 0.935 ;
        RECT  0.410 1.145 1.740 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.995 0.355 2.065 1.070 ;
        RECT  1.890 0.190 1.995 0.425 ;
        RECT  1.890 0.970 1.995 1.070 ;
        RECT  1.225 0.355 1.890 0.425 ;
        RECT  1.365 0.545 1.670 0.615 ;
        RECT  1.180 0.200 1.620 0.275 ;
        RECT  1.510 0.775 1.610 1.075 ;
        RECT  1.295 0.545 1.365 1.055 ;
        RECT  1.180 0.985 1.295 1.055 ;
        RECT  1.155 0.355 1.225 0.660 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.855 0.495 0.945 0.765 ;
        RECT  0.675 0.200 0.920 0.275 ;
        RECT  0.810 0.845 0.910 1.075 ;
        RECT  0.605 0.200 0.675 1.055 ;
        RECT  0.480 0.200 0.605 0.275 ;
        RECT  0.480 0.985 0.605 1.055 ;
        RECT  0.265 0.355 0.335 0.640 ;
        RECT  0.175 0.520 0.265 0.640 ;
        LAYER VIA1 ;
        RECT  1.855 0.665 1.925 0.735 ;
        RECT  1.530 0.945 1.600 1.015 ;
        RECT  1.295 0.805 1.365 0.875 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.865 0.665 0.935 0.735 ;
        RECT  0.825 0.945 0.895 1.015 ;
        RECT  0.605 0.805 0.675 0.875 ;
        RECT  0.265 0.385 0.335 0.455 ;
        LAYER M2 ;
        RECT  0.775 0.945 1.650 1.015 ;
        RECT  0.555 0.805 1.415 0.875 ;
        RECT  0.215 0.385 1.135 0.455 ;
    END
END GXNR2D1BWP

MACRO GXNR2D2BWP
    CLASS CORE ;
    FOREIGN GXNR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 0.420 0.920 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.250 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.665 2.675 0.735 ;
        LAYER M1 ;
        RECT  2.535 0.495 2.625 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.600 -0.115 0.990 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.300 1.145 2.440 1.375 ;
        RECT  1.180 0.985 1.300 1.375 ;
        RECT  0.900 1.145 1.180 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.220 1.145 0.500 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.695 0.355 2.765 1.070 ;
        RECT  2.590 0.190 2.695 0.425 ;
        RECT  2.590 0.970 2.695 1.070 ;
        RECT  1.925 0.355 2.590 0.425 ;
        RECT  2.135 0.545 2.370 0.615 ;
        RECT  1.880 0.200 2.320 0.275 ;
        RECT  2.210 0.775 2.310 1.075 ;
        RECT  2.065 0.545 2.135 1.055 ;
        RECT  1.870 0.985 2.065 1.055 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.560 0.495 1.645 0.765 ;
        RECT  1.435 0.200 1.620 0.275 ;
        RECT  1.510 0.845 1.610 1.075 ;
        RECT  1.365 0.200 1.435 0.875 ;
        RECT  1.250 0.200 1.365 0.275 ;
        RECT  1.090 0.805 1.365 0.875 ;
        RECT  1.180 0.200 1.250 0.415 ;
        RECT  0.910 0.345 1.180 0.415 ;
        RECT  1.010 0.805 1.090 0.965 ;
        RECT  0.810 0.190 0.910 0.415 ;
        RECT  0.485 0.355 0.555 0.640 ;
        RECT  0.175 0.495 0.485 0.640 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.230 0.945 2.300 1.015 ;
        RECT  2.065 0.805 2.135 0.875 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.315 0.805 1.385 0.875 ;
        RECT  0.485 0.385 0.555 0.455 ;
        LAYER M2 ;
        RECT  1.475 0.945 2.350 1.015 ;
        RECT  1.265 0.805 2.185 0.875 ;
        RECT  0.435 0.385 1.835 0.455 ;
    END
END GXNR2D2BWP

MACRO GXOR2D1BWP
    CLASS CORE ;
    FOREIGN GXOR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1224 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.205 0.220 0.275 ;
        RECT  0.105 0.970 0.210 1.070 ;
        RECT  0.035 0.205 0.105 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.550 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.640 ;
        RECT  1.225 0.355 1.855 0.425 ;
        RECT  1.155 0.355 1.225 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 1.145 2.100 1.375 ;
        RECT  1.715 0.805 1.785 1.375 ;
        RECT  0.410 1.145 1.715 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.995 0.205 2.065 0.880 ;
        RECT  1.880 0.205 1.995 0.275 ;
        RECT  1.990 0.800 1.995 0.880 ;
        RECT  1.890 0.800 1.990 1.070 ;
        RECT  1.440 0.545 1.670 0.615 ;
        RECT  1.180 0.200 1.620 0.275 ;
        RECT  1.510 0.855 1.610 1.075 ;
        RECT  1.360 0.545 1.440 1.055 ;
        RECT  1.180 0.985 1.360 1.055 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.875 0.495 0.945 0.875 ;
        RECT  0.665 0.945 0.920 1.055 ;
        RECT  0.815 0.805 0.875 0.875 ;
        RECT  0.665 0.200 0.735 0.875 ;
        RECT  0.480 0.200 0.665 0.275 ;
        RECT  0.590 0.805 0.665 0.875 ;
        RECT  0.490 0.805 0.590 1.070 ;
        RECT  0.175 0.355 0.245 0.675 ;
        RECT  0.735 0.200 0.920 0.275 ;
        LAYER VIA1 ;
        RECT  1.925 0.805 1.995 0.875 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.365 0.665 1.435 0.735 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.845 0.805 0.915 0.875 ;
        RECT  0.695 0.945 0.765 1.015 ;
        RECT  0.665 0.665 0.735 0.735 ;
        RECT  0.175 0.385 0.245 0.455 ;
        LAYER M2 ;
        RECT  0.795 0.805 2.045 0.875 ;
        RECT  0.645 0.945 1.645 1.015 ;
        RECT  0.615 0.665 1.485 0.735 ;
        RECT  0.125 0.385 1.135 0.455 ;
    END
END GXOR2D1BWP

MACRO GXOR2D2BWP
    CLASS CORE ;
    FOREIGN GXOR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 0.420 0.920 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.250 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.640 ;
        RECT  1.925 0.355 2.555 0.425 ;
        RECT  1.855 0.355 1.925 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.600 -0.115 0.990 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.220 -0.115 0.480 0.115 ;
        RECT  0.100 -0.115 0.220 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.485 1.145 2.800 1.375 ;
        RECT  2.415 0.805 2.485 1.375 ;
        RECT  1.280 1.145 2.415 1.375 ;
        RECT  1.200 0.950 1.280 1.375 ;
        RECT  0.900 1.145 1.200 1.375 ;
        RECT  0.820 0.940 0.900 1.375 ;
        RECT  0.580 1.145 0.820 1.375 ;
        RECT  0.500 0.940 0.580 1.375 ;
        RECT  0.220 1.145 0.500 1.375 ;
        RECT  0.100 0.990 0.220 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.695 0.205 2.765 0.880 ;
        RECT  2.580 0.205 2.695 0.275 ;
        RECT  2.690 0.800 2.695 0.880 ;
        RECT  2.590 0.800 2.690 1.070 ;
        RECT  2.140 0.545 2.370 0.615 ;
        RECT  1.880 0.200 2.320 0.275 ;
        RECT  2.210 0.855 2.310 1.075 ;
        RECT  2.060 0.545 2.140 1.055 ;
        RECT  1.880 0.985 2.060 1.055 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.575 0.495 1.645 0.875 ;
        RECT  1.435 0.200 1.620 0.275 ;
        RECT  1.350 0.945 1.620 1.055 ;
        RECT  1.515 0.805 1.575 0.875 ;
        RECT  1.365 0.200 1.435 0.870 ;
        RECT  1.250 0.200 1.365 0.275 ;
        RECT  1.090 0.800 1.365 0.870 ;
        RECT  1.180 0.200 1.250 0.415 ;
        RECT  0.910 0.345 1.180 0.415 ;
        RECT  1.010 0.800 1.090 0.965 ;
        RECT  0.810 0.190 0.910 0.415 ;
        RECT  0.485 0.355 0.555 0.640 ;
        RECT  0.175 0.495 0.485 0.640 ;
        LAYER VIA1 ;
        RECT  2.625 0.805 2.695 0.875 ;
        RECT  2.225 0.945 2.295 1.015 ;
        RECT  2.065 0.665 2.135 0.735 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.545 0.805 1.615 0.875 ;
        RECT  1.395 0.945 1.465 1.015 ;
        RECT  1.365 0.665 1.435 0.735 ;
        RECT  0.485 0.385 0.555 0.455 ;
        LAYER M2 ;
        RECT  1.495 0.805 2.745 0.875 ;
        RECT  1.345 0.945 2.345 1.015 ;
        RECT  1.315 0.665 2.185 0.735 ;
        RECT  0.435 0.385 1.835 0.455 ;
    END
END GXOR2D2BWP

MACRO HA1D0BWP
    CLASS CORE ;
    FOREIGN HA1D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.200 2.345 0.905 ;
        RECT  2.260 0.200 2.275 0.320 ;
        RECT  2.260 0.715 2.275 0.905 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.305 ;
        RECT  0.105 0.930 0.125 1.060 ;
        RECT  0.035 0.185 0.105 1.060 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.985 1.970 1.075 ;
        RECT  1.225 0.985 1.850 1.055 ;
        RECT  1.155 0.870 1.225 1.055 ;
        RECT  0.665 0.870 1.155 0.940 ;
        RECT  0.595 0.705 0.665 0.940 ;
        RECT  0.530 0.705 0.595 0.775 ;
        RECT  0.455 0.495 0.530 0.775 ;
        RECT  0.370 0.495 0.455 0.640 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.625 ;
        RECT  0.660 0.545 0.715 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 -0.115 2.380 0.115 ;
        RECT  2.015 -0.115 2.085 0.445 ;
        RECT  1.080 -0.115 2.015 0.115 ;
        RECT  0.960 -0.115 1.080 0.135 ;
        RECT  0.340 -0.115 0.960 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.145 2.380 1.375 ;
        RECT  0.960 1.010 1.080 1.375 ;
        RECT  0.710 1.145 0.960 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.520 2.190 0.915 ;
        RECT  1.470 0.845 2.120 0.915 ;
        RECT  1.815 0.185 1.885 0.775 ;
        RECT  1.750 0.500 1.815 0.620 ;
        RECT  1.605 0.205 1.680 0.775 ;
        RECT  1.070 0.205 1.605 0.275 ;
        RECT  1.550 0.705 1.605 0.775 ;
        RECT  1.470 0.345 1.525 0.415 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.330 0.845 1.400 0.915 ;
        RECT  1.200 0.355 1.270 0.800 ;
        RECT  1.150 0.355 1.200 0.425 ;
        RECT  1.150 0.730 1.200 0.800 ;
        RECT  1.070 0.520 1.130 0.640 ;
        RECT  1.000 0.205 1.070 0.800 ;
        RECT  0.880 0.205 1.000 0.285 ;
        RECT  0.770 0.730 1.000 0.800 ;
        RECT  0.770 0.185 0.880 0.285 ;
        RECT  0.600 0.185 0.700 0.285 ;
        RECT  0.535 0.210 0.600 0.285 ;
        RECT  0.465 0.210 0.535 0.415 ;
        RECT  0.435 0.845 0.505 1.025 ;
        RECT  0.265 0.345 0.465 0.415 ;
        RECT  0.265 0.845 0.435 0.915 ;
        RECT  0.195 0.345 0.265 0.915 ;
        RECT  0.175 0.520 0.195 0.640 ;
    END
END HA1D0BWP

MACRO HA1D1BWP
    CLASS CORE ;
    FOREIGN HA1D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.045 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.735 2.415 1.045 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.725 0.125 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.0720 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 0.995 2.060 1.075 ;
        RECT  0.945 0.995 1.920 1.065 ;
        RECT  0.875 0.870 0.945 1.065 ;
        RECT  0.665 0.870 0.875 0.940 ;
        RECT  0.595 0.545 0.665 0.940 ;
        RECT  0.340 0.545 0.595 0.615 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.545 0.900 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.260 0.140 ;
        RECT  1.245 -0.115 2.140 0.115 ;
        RECT  1.135 -0.115 1.245 0.265 ;
        RECT  0.870 -0.115 1.135 0.115 ;
        RECT  0.790 -0.115 0.870 0.270 ;
        RECT  0.335 -0.115 0.790 0.115 ;
        RECT  0.215 -0.115 0.335 0.275 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.145 2.520 1.375 ;
        RECT  2.160 0.710 2.240 1.375 ;
        RECT  1.180 1.145 2.160 1.375 ;
        RECT  1.060 1.135 1.180 1.375 ;
        RECT  0.740 1.145 1.060 1.375 ;
        RECT  0.620 1.010 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.860 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 0.520 2.320 0.640 ;
        RECT  2.190 0.210 2.260 0.640 ;
        RECT  1.585 0.210 2.190 0.280 ;
        RECT  1.955 0.350 2.025 0.925 ;
        RECT  1.810 0.520 1.955 0.600 ;
        RECT  1.740 0.855 1.830 0.925 ;
        RECT  1.740 0.350 1.810 0.420 ;
        RECT  1.670 0.350 1.740 0.925 ;
        RECT  1.170 0.855 1.670 0.925 ;
        RECT  1.510 0.210 1.585 0.785 ;
        RECT  1.360 0.215 1.430 0.785 ;
        RECT  1.335 0.215 1.360 0.335 ;
        RECT  1.270 0.715 1.360 0.785 ;
        RECT  1.170 0.510 1.290 0.630 ;
        RECT  1.100 0.410 1.170 0.925 ;
        RECT  1.045 0.410 1.100 0.480 ;
        RECT  0.830 0.730 1.100 0.800 ;
        RECT  0.975 0.220 1.045 0.480 ;
        RECT  0.540 0.205 0.710 0.275 ;
        RECT  0.470 0.205 0.540 0.415 ;
        RECT  0.435 0.710 0.505 1.000 ;
        RECT  0.265 0.345 0.470 0.415 ;
        RECT  0.265 0.710 0.435 0.780 ;
        RECT  0.195 0.345 0.265 0.780 ;
        RECT  0.180 0.520 0.195 0.640 ;
    END
END HA1D1BWP

MACRO HA1D2BWP
    CLASS CORE ;
    FOREIGN HA1D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.565 0.355 2.625 0.805 ;
        RECT  2.555 0.185 2.565 1.035 ;
        RECT  2.495 0.185 2.555 0.465 ;
        RECT  2.495 0.735 2.555 1.035 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.185 0.300 0.465 ;
        RECT  0.245 0.735 0.300 1.035 ;
        RECT  0.230 0.185 0.245 1.035 ;
        RECT  0.175 0.355 0.230 0.900 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.0718 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.985 2.205 1.075 ;
        RECT  0.870 0.985 2.060 1.055 ;
        RECT  0.800 0.705 0.870 1.055 ;
        RECT  0.665 0.705 0.800 0.775 ;
        RECT  0.595 0.495 0.665 0.775 ;
        RECT  0.520 0.495 0.595 0.640 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.545 1.040 0.625 ;
        RECT  0.875 0.355 0.945 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.300 ;
        RECT  2.400 -0.115 2.670 0.115 ;
        RECT  2.280 -0.115 2.400 0.135 ;
        RECT  1.410 -0.115 2.280 0.115 ;
        RECT  1.290 -0.115 1.410 0.265 ;
        RECT  1.030 -0.115 1.290 0.115 ;
        RECT  0.950 -0.115 1.030 0.275 ;
        RECT  0.510 -0.115 0.950 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.390 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.895 2.750 1.375 ;
        RECT  2.360 1.145 2.670 1.375 ;
        RECT  2.280 0.735 2.360 1.375 ;
        RECT  1.340 1.145 2.280 1.375 ;
        RECT  1.220 1.130 1.340 1.375 ;
        RECT  0.520 1.145 1.220 1.375 ;
        RECT  0.400 1.000 0.520 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.970 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.360 0.545 2.480 0.615 ;
        RECT  2.290 0.205 2.360 0.615 ;
        RECT  1.745 0.205 2.290 0.275 ;
        RECT  2.145 0.345 2.185 0.580 ;
        RECT  2.115 0.345 2.145 0.820 ;
        RECT  2.075 0.510 2.115 0.820 ;
        RECT  2.000 0.510 2.075 0.630 ;
        RECT  1.930 0.345 1.990 0.415 ;
        RECT  1.930 0.845 1.990 0.915 ;
        RECT  1.860 0.345 1.930 0.915 ;
        RECT  1.205 0.845 1.860 0.915 ;
        RECT  1.745 0.695 1.790 0.765 ;
        RECT  1.670 0.205 1.745 0.765 ;
        RECT  1.520 0.205 1.590 0.765 ;
        RECT  1.495 0.205 1.520 0.325 ;
        RECT  1.430 0.695 1.520 0.765 ;
        RECT  1.205 0.500 1.450 0.620 ;
        RECT  1.135 0.210 1.205 0.915 ;
        RECT  1.000 0.845 1.135 0.915 ;
        RECT  0.685 0.205 0.870 0.275 ;
        RECT  0.615 0.205 0.685 0.415 ;
        RECT  0.615 0.850 0.685 1.000 ;
        RECT  0.440 0.345 0.615 0.415 ;
        RECT  0.440 0.850 0.615 0.920 ;
        RECT  0.370 0.345 0.440 0.920 ;
        RECT  0.320 0.545 0.370 0.615 ;
    END
END HA1D2BWP

MACRO HA1D4BWP
    CLASS CORE ;
    FOREIGN HA1D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.465 ;
        RECT  3.955 0.700 3.965 1.075 ;
        RECT  3.895 0.185 3.955 1.075 ;
        RECT  3.745 0.345 3.895 0.905 ;
        RECT  3.605 0.345 3.745 0.465 ;
        RECT  3.605 0.700 3.745 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.700 3.605 1.075 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.700 0.665 1.075 ;
        RECT  0.455 0.345 0.595 0.465 ;
        RECT  0.455 0.700 0.595 0.905 ;
        RECT  0.305 0.345 0.455 0.905 ;
        RECT  0.245 0.185 0.305 1.075 ;
        RECT  0.235 0.185 0.245 0.465 ;
        RECT  0.235 0.700 0.245 1.075 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.155 0.990 3.275 1.075 ;
        RECT  1.925 0.990 3.155 1.060 ;
        RECT  1.855 0.870 1.925 1.060 ;
        RECT  1.560 0.870 1.855 0.940 ;
        RECT  1.490 0.730 1.560 0.940 ;
        RECT  1.455 0.730 1.490 0.800 ;
        RECT  1.385 0.515 1.455 0.800 ;
        RECT  0.960 0.730 1.385 0.800 ;
        RECT  0.875 0.495 0.960 0.800 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.1440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.605 0.495 1.785 0.625 ;
        RECT  1.535 0.355 1.605 0.625 ;
        RECT  1.225 0.355 1.535 0.425 ;
        RECT  1.155 0.355 1.225 0.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 -0.115 4.200 0.115 ;
        RECT  4.075 -0.115 4.145 0.465 ;
        RECT  3.810 -0.115 4.075 0.115 ;
        RECT  3.690 -0.115 3.810 0.265 ;
        RECT  3.440 -0.115 3.690 0.115 ;
        RECT  3.320 -0.115 3.440 0.135 ;
        RECT  2.490 -0.115 3.320 0.115 ;
        RECT  2.370 -0.115 2.490 0.235 ;
        RECT  1.925 -0.115 2.370 0.115 ;
        RECT  1.855 -0.115 1.925 0.275 ;
        RECT  1.565 -0.115 1.855 0.115 ;
        RECT  1.495 -0.115 1.565 0.275 ;
        RECT  0.845 -0.115 1.495 0.115 ;
        RECT  0.775 -0.115 0.845 0.270 ;
        RECT  0.510 -0.115 0.775 0.115 ;
        RECT  0.390 -0.115 0.510 0.265 ;
        RECT  0.125 -0.115 0.390 0.115 ;
        RECT  0.055 -0.115 0.125 0.475 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 1.145 4.200 1.375 ;
        RECT  4.075 0.700 4.145 1.375 ;
        RECT  3.810 1.145 4.075 1.375 ;
        RECT  3.690 0.985 3.810 1.375 ;
        RECT  3.425 1.145 3.690 1.375 ;
        RECT  3.355 0.695 3.425 1.375 ;
        RECT  2.520 1.145 3.355 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  1.960 1.145 2.400 1.375 ;
        RECT  1.840 1.130 1.960 1.375 ;
        RECT  1.590 1.145 1.840 1.375 ;
        RECT  1.470 1.010 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.010 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.010 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.125 1.145 0.390 1.375 ;
        RECT  0.055 0.680 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.345 3.675 0.465 ;
        RECT  3.605 0.700 3.675 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.700 3.605 1.075 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.700 0.665 1.075 ;
        RECT  0.525 0.345 0.595 0.465 ;
        RECT  0.525 0.700 0.595 0.905 ;
        RECT  3.430 0.545 3.635 0.615 ;
        RECT  3.360 0.205 3.430 0.615 ;
        RECT  2.845 0.205 3.360 0.275 ;
        RECT  3.175 0.345 3.245 0.885 ;
        RECT  3.155 0.345 3.175 0.640 ;
        RECT  3.090 0.520 3.155 0.640 ;
        RECT  3.020 0.850 3.090 0.920 ;
        RECT  3.020 0.355 3.070 0.435 ;
        RECT  2.950 0.355 3.020 0.920 ;
        RECT  2.125 0.850 2.950 0.920 ;
        RECT  2.845 0.680 2.880 0.780 ;
        RECT  2.770 0.205 2.845 0.780 ;
        RECT  2.645 0.395 2.685 0.780 ;
        RECT  2.615 0.200 2.645 0.780 ;
        RECT  2.575 0.200 2.615 0.460 ;
        RECT  2.210 0.710 2.615 0.780 ;
        RECT  2.285 0.380 2.575 0.460 ;
        RECT  2.125 0.545 2.500 0.615 ;
        RECT  2.215 0.200 2.285 0.460 ;
        RECT  2.105 0.545 2.125 0.920 ;
        RECT  2.055 0.200 2.105 0.920 ;
        RECT  2.035 0.200 2.055 0.800 ;
        RECT  1.745 0.345 2.035 0.415 ;
        RECT  1.640 0.730 2.035 0.800 ;
        RECT  1.675 0.230 1.745 0.415 ;
        RECT  0.805 0.870 1.410 0.940 ;
        RECT  1.030 0.215 1.240 0.285 ;
        RECT  0.960 0.215 1.030 0.410 ;
        RECT  0.805 0.340 0.960 0.410 ;
        RECT  0.735 0.340 0.805 0.940 ;
        RECT  0.630 0.545 0.735 0.615 ;
    END
END HA1D4BWP

MACRO HCOSCIND1BWP
    CLASS CORE ;
    FOREIGN HCOSCIND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.185 4.445 1.045 ;
        RECT  4.355 0.185 4.375 0.465 ;
        RECT  4.355 0.750 4.375 1.045 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.465 0.765 ;
        RECT  3.325 0.635 3.395 0.765 ;
        END
    END CS
    PIN CO
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.730 0.125 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 2.905 0.765 ;
        RECT  2.760 0.495 2.835 0.635 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.1440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.625 ;
        RECT  0.625 0.545 0.875 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 -0.115 4.480 0.115 ;
        RECT  4.155 -0.115 4.245 0.440 ;
        RECT  3.340 -0.115 4.155 0.115 ;
        RECT  3.220 -0.115 3.340 0.135 ;
        RECT  2.940 -0.115 3.220 0.115 ;
        RECT  2.820 -0.115 2.940 0.130 ;
        RECT  2.640 -0.115 2.820 0.115 ;
        RECT  2.520 -0.115 2.640 0.130 ;
        RECT  1.660 -0.115 2.520 0.115 ;
        RECT  1.540 -0.115 1.660 0.130 ;
        RECT  1.260 -0.115 1.540 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.340 -0.115 1.140 0.115 ;
        RECT  0.220 -0.115 0.340 0.255 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.145 4.480 1.375 ;
        RECT  4.140 1.065 4.260 1.375 ;
        RECT  2.930 1.145 4.140 1.375 ;
        RECT  2.850 0.890 2.930 1.375 ;
        RECT  1.590 1.145 2.850 1.375 ;
        RECT  1.470 1.030 1.590 1.375 ;
        RECT  1.160 1.145 1.470 1.375 ;
        RECT  1.040 1.030 1.160 1.375 ;
        RECT  0.740 1.145 1.040 1.375 ;
        RECT  0.620 1.030 0.740 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 0.995 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.275 0.520 4.290 0.640 ;
        RECT  4.205 0.520 4.275 0.995 ;
        RECT  3.670 0.925 4.205 0.995 ;
        RECT  3.975 0.340 4.045 0.845 ;
        RECT  3.910 0.520 3.975 0.640 ;
        RECT  3.825 0.205 3.890 0.275 ;
        RECT  3.825 0.765 3.890 0.835 ;
        RECT  3.755 0.205 3.825 0.835 ;
        RECT  2.550 0.205 3.755 0.275 ;
        RECT  3.595 0.345 3.670 0.995 ;
        RECT  3.105 0.345 3.510 0.415 ;
        RECT  3.390 0.845 3.510 1.060 ;
        RECT  3.105 0.845 3.390 0.925 ;
        RECT  3.035 0.345 3.105 1.070 ;
        RECT  3.020 0.345 3.035 0.415 ;
        RECT  2.690 0.345 2.790 0.415 ;
        RECT  2.690 0.730 2.740 0.850 ;
        RECT  2.620 0.345 2.690 1.055 ;
        RECT  1.750 0.980 2.620 1.055 ;
        RECT  2.480 0.205 2.550 0.910 ;
        RECT  1.980 0.840 2.480 0.910 ;
        RECT  2.330 0.325 2.400 0.770 ;
        RECT  2.280 0.510 2.330 0.770 ;
        RECT  2.250 0.510 2.280 0.630 ;
        RECT  2.180 0.365 2.250 0.435 ;
        RECT  2.110 0.205 2.180 0.770 ;
        RECT  1.175 0.205 2.110 0.275 ;
        RECT  2.060 0.690 2.110 0.770 ;
        RECT  1.980 0.345 2.040 0.465 ;
        RECT  1.910 0.345 1.980 0.910 ;
        RECT  1.850 0.840 1.910 0.910 ;
        RECT  1.710 0.345 1.780 0.815 ;
        RECT  1.680 0.890 1.750 1.055 ;
        RECT  1.330 0.345 1.710 0.415 ;
        RECT  1.270 0.745 1.710 0.815 ;
        RECT  0.725 0.890 1.680 0.960 ;
        RECT  1.175 0.545 1.415 0.615 ;
        RECT  1.105 0.205 1.175 0.815 ;
        RECT  0.950 0.205 1.105 0.275 ;
        RECT  0.840 0.745 1.105 0.815 ;
        RECT  0.645 0.705 0.725 0.960 ;
        RECT  0.610 0.190 0.690 0.450 ;
        RECT  0.445 0.705 0.645 0.775 ;
        RECT  0.280 0.380 0.610 0.450 ;
        RECT  0.410 0.845 0.530 1.055 ;
        RECT  0.370 0.520 0.445 0.775 ;
        RECT  0.280 0.845 0.410 0.915 ;
        RECT  0.210 0.380 0.280 0.915 ;
        RECT  0.175 0.520 0.210 0.640 ;
    END
END HCOSCIND1BWP

MACRO HCOSCIND2BWP
    CLASS CORE ;
    FOREIGN HCOSCIND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.665 0.355 4.725 0.780 ;
        RECT  4.655 0.185 4.665 1.035 ;
        RECT  4.595 0.185 4.655 0.465 ;
        RECT  4.595 0.710 4.655 1.035 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.510 0.495 3.605 0.765 ;
        END
    END CS
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.185 0.300 0.465 ;
        RECT  0.245 0.770 0.300 1.050 ;
        RECT  0.230 0.185 0.245 1.050 ;
        RECT  0.175 0.355 0.230 0.840 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.355 3.185 0.630 ;
        RECT  2.960 0.495 3.115 0.630 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.1440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.350 1.085 0.625 ;
        RECT  0.765 0.545 1.015 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.115 4.900 0.115 ;
        RECT  4.770 -0.115 4.850 0.300 ;
        RECT  4.460 -0.115 4.770 0.115 ;
        RECT  4.380 -0.115 4.460 0.460 ;
        RECT  3.540 -0.115 4.380 0.115 ;
        RECT  3.420 -0.115 3.540 0.135 ;
        RECT  3.140 -0.115 3.420 0.115 ;
        RECT  3.020 -0.115 3.140 0.130 ;
        RECT  2.840 -0.115 3.020 0.115 ;
        RECT  2.720 -0.115 2.840 0.130 ;
        RECT  1.840 -0.115 2.720 0.115 ;
        RECT  1.720 -0.115 1.840 0.130 ;
        RECT  1.440 -0.115 1.720 0.115 ;
        RECT  1.320 -0.115 1.440 0.135 ;
        RECT  0.520 -0.115 1.320 0.115 ;
        RECT  0.400 -0.115 0.520 0.260 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 1.145 4.900 1.375 ;
        RECT  4.770 0.850 4.850 1.375 ;
        RECT  3.130 1.145 4.770 1.375 ;
        RECT  3.050 0.750 3.130 1.375 ;
        RECT  1.790 1.145 3.050 1.375 ;
        RECT  1.670 1.030 1.790 1.375 ;
        RECT  1.360 1.145 1.670 1.375 ;
        RECT  1.240 1.030 1.360 1.375 ;
        RECT  0.960 1.145 1.240 1.375 ;
        RECT  0.840 1.030 0.960 1.375 ;
        RECT  0.520 1.145 0.840 1.375 ;
        RECT  0.440 0.995 0.520 1.375 ;
        RECT  0.130 1.145 0.440 1.375 ;
        RECT  0.050 0.910 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.465 0.545 4.585 0.615 ;
        RECT  4.395 0.545 4.465 0.960 ;
        RECT  3.870 0.890 4.395 0.960 ;
        RECT  4.175 0.335 4.245 0.810 ;
        RECT  4.105 0.520 4.175 0.640 ;
        RECT  4.025 0.205 4.090 0.275 ;
        RECT  4.025 0.740 4.090 0.810 ;
        RECT  3.955 0.205 4.025 0.810 ;
        RECT  2.750 0.205 3.955 0.275 ;
        RECT  3.795 0.345 3.870 0.960 ;
        RECT  3.330 0.345 3.710 0.415 ;
        RECT  3.590 0.845 3.710 1.060 ;
        RECT  3.330 0.845 3.590 0.925 ;
        RECT  3.305 0.345 3.330 0.925 ;
        RECT  3.260 0.345 3.305 1.035 ;
        RECT  3.235 0.750 3.260 1.035 ;
        RECT  2.890 0.345 2.990 0.415 ;
        RECT  2.890 0.725 2.940 0.845 ;
        RECT  2.820 0.345 2.890 1.055 ;
        RECT  1.950 0.980 2.820 1.055 ;
        RECT  2.680 0.205 2.750 0.910 ;
        RECT  2.180 0.840 2.680 0.910 ;
        RECT  2.530 0.325 2.600 0.770 ;
        RECT  2.480 0.510 2.530 0.770 ;
        RECT  2.450 0.510 2.480 0.630 ;
        RECT  2.380 0.365 2.450 0.435 ;
        RECT  2.310 0.205 2.380 0.770 ;
        RECT  1.350 0.205 2.310 0.275 ;
        RECT  2.260 0.690 2.310 0.770 ;
        RECT  2.180 0.345 2.240 0.465 ;
        RECT  2.110 0.345 2.180 0.910 ;
        RECT  2.050 0.840 2.110 0.910 ;
        RECT  1.910 0.345 1.980 0.815 ;
        RECT  1.880 0.890 1.950 1.055 ;
        RECT  1.510 0.345 1.910 0.415 ;
        RECT  1.470 0.745 1.910 0.815 ;
        RECT  0.945 0.890 1.880 0.960 ;
        RECT  1.350 0.545 1.595 0.615 ;
        RECT  1.280 0.205 1.350 0.815 ;
        RECT  1.130 0.205 1.280 0.275 ;
        RECT  1.050 0.745 1.280 0.815 ;
        RECT  0.865 0.705 0.945 0.960 ;
        RECT  0.795 0.190 0.865 0.450 ;
        RECT  0.625 0.705 0.865 0.775 ;
        RECT  0.440 0.380 0.795 0.450 ;
        RECT  0.630 0.845 0.750 1.055 ;
        RECT  0.440 0.845 0.630 0.915 ;
        RECT  0.550 0.520 0.625 0.775 ;
        RECT  0.370 0.380 0.440 0.915 ;
        RECT  0.315 0.545 0.370 0.615 ;
    END
END HCOSCIND2BWP

MACRO HCOSCOND1BWP
    CLASS CORE ;
    FOREIGN HCOSCOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.750 3.955 1.045 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.640 2.975 0.765 ;
        RECT  2.835 0.495 2.905 0.765 ;
        END
    END CS
    PIN CON
        ANTENNADIFFAREA 0.0997 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.510 0.285 ;
        RECT  0.310 0.215 0.385 0.770 ;
        RECT  0.210 0.700 0.310 0.770 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0560 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.985 2.290 1.055 ;
        RECT  1.480 0.870 1.550 1.055 ;
        RECT  0.510 0.870 1.480 0.940 ;
        RECT  0.440 0.845 0.510 0.940 ;
        RECT  0.105 0.845 0.440 0.915 ;
        RECT  0.105 0.495 0.210 0.630 ;
        RECT  0.035 0.495 0.105 0.915 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.1440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.740 -0.115 3.820 0.420 ;
        RECT  2.890 -0.115 3.740 0.115 ;
        RECT  2.770 -0.115 2.890 0.135 ;
        RECT  2.480 -0.115 2.770 0.115 ;
        RECT  2.360 -0.115 2.480 0.135 ;
        RECT  1.500 -0.115 2.360 0.115 ;
        RECT  1.380 -0.115 1.500 0.130 ;
        RECT  1.080 -0.115 1.380 0.115 ;
        RECT  0.960 -0.115 1.080 0.135 ;
        RECT  0.670 -0.115 0.960 0.115 ;
        RECT  0.590 -0.115 0.670 0.420 ;
        RECT  0.130 -0.115 0.590 0.115 ;
        RECT  0.050 -0.115 0.130 0.345 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 1.145 4.060 1.375 ;
        RECT  3.720 1.075 3.840 1.375 ;
        RECT  2.870 1.145 3.720 1.375 ;
        RECT  2.750 1.010 2.870 1.375 ;
        RECT  2.490 1.145 2.750 1.375 ;
        RECT  2.370 1.000 2.490 1.375 ;
        RECT  1.390 1.145 2.370 1.375 ;
        RECT  1.270 1.010 1.390 1.375 ;
        RECT  0.950 1.145 1.270 1.375 ;
        RECT  0.830 1.010 0.950 1.375 ;
        RECT  0.560 1.145 0.830 1.375 ;
        RECT  0.440 1.010 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.990 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.855 0.520 3.870 0.640 ;
        RECT  3.785 0.520 3.855 0.995 ;
        RECT  3.250 0.925 3.785 0.995 ;
        RECT  3.555 0.340 3.625 0.845 ;
        RECT  3.490 0.520 3.555 0.640 ;
        RECT  3.405 0.770 3.470 0.840 ;
        RECT  3.405 0.205 3.460 0.275 ;
        RECT  3.335 0.205 3.405 0.840 ;
        RECT  2.450 0.205 3.335 0.275 ;
        RECT  3.180 0.345 3.250 0.995 ;
        RECT  3.155 0.345 3.180 0.465 ;
        RECT  2.970 0.860 3.090 1.070 ;
        RECT  2.655 0.345 3.070 0.415 ;
        RECT  2.655 0.860 2.970 0.930 ;
        RECT  2.585 0.345 2.655 1.070 ;
        RECT  2.370 0.205 2.450 0.915 ;
        RECT  1.725 0.845 2.370 0.915 ;
        RECT  2.225 0.335 2.265 0.600 ;
        RECT  2.195 0.335 2.225 0.775 ;
        RECT  2.155 0.515 2.195 0.775 ;
        RECT  2.090 0.515 2.155 0.640 ;
        RECT  2.020 0.360 2.100 0.430 ;
        RECT  1.950 0.205 2.020 0.775 ;
        RECT  0.845 0.205 1.950 0.275 ;
        RECT  1.890 0.705 1.950 0.775 ;
        RECT  1.810 0.360 1.880 0.625 ;
        RECT  1.725 0.555 1.810 0.625 ;
        RECT  1.655 0.555 1.725 0.915 ;
        RECT  1.265 0.345 1.660 0.415 ;
        RECT  1.265 0.730 1.570 0.800 ;
        RECT  1.195 0.345 1.265 0.800 ;
        RECT  1.060 0.730 1.195 0.800 ;
        RECT  0.850 0.520 1.100 0.640 ;
        RECT  0.845 0.520 0.850 0.790 ;
        RECT  0.775 0.205 0.845 0.790 ;
        RECT  0.640 0.720 0.775 0.790 ;
    END
END HCOSCOND1BWP

MACRO HCOSCOND2BWP
    CLASS CORE ;
    FOREIGN HCOSCOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.355 4.445 0.790 ;
        RECT  4.305 0.185 4.375 0.465 ;
        RECT  4.305 0.720 4.375 1.035 ;
        END
    END S
    PIN CS
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 0.495 3.325 0.765 ;
        END
    END CS
    PIN CON
        ANTENNADIFFAREA 0.1644 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.700 0.730 0.770 ;
        RECT  0.385 0.205 0.540 0.275 ;
        RECT  0.310 0.205 0.385 0.770 ;
        RECT  0.230 0.700 0.310 0.770 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0848 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 0.985 2.610 1.055 ;
        RECT  1.800 0.870 1.870 1.055 ;
        RECT  0.880 0.870 1.800 0.940 ;
        RECT  0.810 0.495 0.880 0.940 ;
        RECT  0.710 0.495 0.810 0.625 ;
        RECT  0.365 0.870 0.810 0.940 ;
        RECT  0.295 0.840 0.365 0.940 ;
        RECT  0.105 0.840 0.295 0.910 ;
        RECT  0.105 0.495 0.230 0.630 ;
        RECT  0.035 0.495 0.105 0.910 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.1728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.355 1.085 0.640 ;
        RECT  0.555 0.355 1.005 0.425 ;
        RECT  0.455 0.355 0.555 0.630 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.300 ;
        RECT  4.180 -0.115 4.490 0.115 ;
        RECT  4.100 -0.115 4.180 0.450 ;
        RECT  3.210 -0.115 4.100 0.115 ;
        RECT  3.090 -0.115 3.210 0.135 ;
        RECT  2.800 -0.115 3.090 0.115 ;
        RECT  2.680 -0.115 2.800 0.135 ;
        RECT  1.790 -0.115 2.680 0.115 ;
        RECT  1.670 -0.115 1.790 0.135 ;
        RECT  0.890 -0.115 1.670 0.115 ;
        RECT  0.810 -0.115 0.890 0.275 ;
        RECT  0.140 -0.115 0.810 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.865 4.570 1.375 ;
        RECT  4.200 1.145 4.490 1.375 ;
        RECT  4.080 1.030 4.200 1.375 ;
        RECT  3.190 1.145 4.080 1.375 ;
        RECT  3.070 1.005 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 1.000 2.810 1.375 ;
        RECT  1.710 1.145 2.690 1.375 ;
        RECT  1.590 1.015 1.710 1.375 ;
        RECT  1.270 1.145 1.590 1.375 ;
        RECT  1.150 1.010 1.270 1.375 ;
        RECT  0.910 1.145 1.150 1.375 ;
        RECT  0.790 1.010 0.910 1.375 ;
        RECT  0.540 1.145 0.790 1.375 ;
        RECT  0.420 1.010 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.990 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.150 0.545 4.305 0.615 ;
        RECT  4.080 0.545 4.150 0.960 ;
        RECT  3.575 0.890 4.080 0.960 ;
        RECT  3.875 0.335 3.945 0.810 ;
        RECT  3.785 0.510 3.875 0.630 ;
        RECT  3.715 0.740 3.790 0.810 ;
        RECT  3.715 0.205 3.780 0.275 ;
        RECT  3.645 0.205 3.715 0.810 ;
        RECT  2.770 0.205 3.645 0.275 ;
        RECT  3.570 0.890 3.575 1.060 ;
        RECT  3.500 0.345 3.570 1.060 ;
        RECT  3.475 0.345 3.500 0.465 ;
        RECT  3.290 0.865 3.410 1.075 ;
        RECT  2.980 0.345 3.390 0.415 ;
        RECT  2.980 0.865 3.290 0.935 ;
        RECT  2.900 0.345 2.980 1.070 ;
        RECT  2.690 0.205 2.770 0.915 ;
        RECT  2.045 0.845 2.690 0.915 ;
        RECT  2.545 0.335 2.585 0.600 ;
        RECT  2.515 0.335 2.545 0.775 ;
        RECT  2.475 0.515 2.515 0.775 ;
        RECT  2.410 0.515 2.475 0.640 ;
        RECT  2.340 0.360 2.410 0.430 ;
        RECT  2.270 0.205 2.340 0.775 ;
        RECT  1.265 0.205 2.270 0.275 ;
        RECT  2.210 0.705 2.270 0.775 ;
        RECT  2.130 0.360 2.200 0.625 ;
        RECT  2.045 0.555 2.130 0.625 ;
        RECT  1.975 0.555 2.045 0.915 ;
        RECT  1.730 0.345 1.970 0.415 ;
        RECT  1.730 0.730 1.890 0.800 ;
        RECT  1.660 0.345 1.730 0.800 ;
        RECT  1.420 0.345 1.660 0.415 ;
        RECT  1.380 0.730 1.660 0.800 ;
        RECT  1.265 0.545 1.525 0.615 ;
        RECT  1.195 0.205 1.265 0.790 ;
        RECT  0.990 0.205 1.195 0.275 ;
        RECT  0.970 0.720 1.195 0.790 ;
    END
END HCOSCOND2BWP

MACRO HICIND1BWP
    CLASS CORE ;
    FOREIGN HICIND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.765 1.045 ;
        RECT  2.675 0.185 2.695 0.465 ;
        RECT  2.675 0.735 2.695 1.045 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.735 0.125 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.670 0.765 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.545 0.910 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 -0.115 2.800 0.115 ;
        RECT  2.480 -0.115 2.560 0.420 ;
        RECT  1.650 -0.115 2.480 0.115 ;
        RECT  1.530 -0.115 1.650 0.135 ;
        RECT  1.260 -0.115 1.530 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.865 -0.115 1.140 0.115 ;
        RECT  0.795 -0.115 0.865 0.280 ;
        RECT  0.340 -0.115 0.795 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.145 2.800 1.375 ;
        RECT  2.460 1.010 2.580 1.375 ;
        RECT  1.590 1.145 2.460 1.375 ;
        RECT  1.470 1.125 1.590 1.375 ;
        RECT  1.180 1.145 1.470 1.375 ;
        RECT  1.060 1.010 1.180 1.375 ;
        RECT  0.740 1.145 1.060 1.375 ;
        RECT  0.620 1.010 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.520 2.620 0.640 ;
        RECT  2.480 0.520 2.550 0.940 ;
        RECT  2.235 0.870 2.480 0.940 ;
        RECT  2.295 0.185 2.365 0.790 ;
        RECT  2.200 0.515 2.295 0.635 ;
        RECT  2.165 0.845 2.235 0.940 ;
        RECT  2.130 0.705 2.190 0.775 ;
        RECT  2.130 0.205 2.185 0.330 ;
        RECT  1.980 0.845 2.165 0.915 ;
        RECT  2.060 0.205 2.130 0.775 ;
        RECT  1.960 0.985 2.080 1.065 ;
        RECT  1.045 0.205 2.060 0.275 ;
        RECT  1.910 0.345 1.980 0.915 ;
        RECT  1.365 0.985 1.960 1.055 ;
        RECT  1.760 0.345 1.830 0.915 ;
        RECT  1.330 0.345 1.760 0.415 ;
        RECT  1.505 0.845 1.760 0.915 ;
        RECT  1.435 0.730 1.505 0.915 ;
        RECT  1.260 0.730 1.435 0.800 ;
        RECT  1.295 0.870 1.365 1.055 ;
        RECT  1.160 0.545 1.360 0.615 ;
        RECT  0.715 0.870 1.295 0.940 ;
        RECT  1.090 0.415 1.160 0.800 ;
        RECT  1.045 0.415 1.090 0.485 ;
        RECT  0.840 0.730 1.090 0.800 ;
        RECT  0.975 0.205 1.045 0.485 ;
        RECT  0.645 0.705 0.715 0.940 ;
        RECT  0.535 0.210 0.710 0.280 ;
        RECT  0.435 0.705 0.645 0.775 ;
        RECT  0.465 0.210 0.535 0.415 ;
        RECT  0.435 0.845 0.505 1.000 ;
        RECT  0.275 0.345 0.465 0.415 ;
        RECT  0.365 0.520 0.435 0.775 ;
        RECT  0.275 0.845 0.435 0.915 ;
        RECT  0.205 0.345 0.275 0.915 ;
        RECT  0.180 0.520 0.205 0.640 ;
    END
END HICIND1BWP

MACRO HICIND2BWP
    CLASS CORE ;
    FOREIGN HICIND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.355 3.045 0.805 ;
        RECT  2.975 0.185 2.985 1.035 ;
        RECT  2.915 0.185 2.975 0.465 ;
        RECT  2.915 0.735 2.975 1.035 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.185 0.300 0.465 ;
        RECT  0.230 0.735 0.300 1.035 ;
        RECT  0.105 0.355 0.230 0.425 ;
        RECT  0.105 0.735 0.230 0.805 ;
        RECT  0.035 0.355 0.105 0.805 ;
        END
    END CO
    PIN CIN
        ANTENNAGATEAREA 0.0488 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 1.840 0.660 ;
        RECT  1.710 0.495 1.785 0.765 ;
        END
    END CIN
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.625 ;
        RECT  0.900 0.540 1.155 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.300 ;
        RECT  2.780 -0.115 3.090 0.115 ;
        RECT  2.700 -0.115 2.780 0.465 ;
        RECT  1.810 -0.115 2.700 0.115 ;
        RECT  1.690 -0.115 1.810 0.135 ;
        RECT  1.420 -0.115 1.690 0.115 ;
        RECT  1.300 -0.115 1.420 0.135 ;
        RECT  1.025 -0.115 1.300 0.115 ;
        RECT  0.955 -0.115 1.025 0.420 ;
        RECT  0.510 -0.115 0.955 0.115 ;
        RECT  0.390 -0.115 0.510 0.280 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.280 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.875 3.170 1.375 ;
        RECT  2.800 1.145 3.090 1.375 ;
        RECT  2.680 1.020 2.800 1.375 ;
        RECT  1.750 1.145 2.680 1.375 ;
        RECT  1.630 1.125 1.750 1.375 ;
        RECT  1.340 1.145 1.630 1.375 ;
        RECT  1.220 1.125 1.340 1.375 ;
        RECT  0.920 1.145 1.220 1.375 ;
        RECT  0.800 1.010 0.920 1.375 ;
        RECT  0.520 1.145 0.800 1.375 ;
        RECT  0.400 1.010 0.520 1.375 ;
        RECT  0.125 1.145 0.400 1.375 ;
        RECT  0.055 0.905 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.830 0.545 2.900 0.615 ;
        RECT  2.760 0.545 2.830 0.950 ;
        RECT  2.415 0.880 2.760 0.950 ;
        RECT  2.495 0.185 2.565 0.810 ;
        RECT  2.370 0.470 2.495 0.590 ;
        RECT  2.345 0.845 2.415 0.950 ;
        RECT  2.300 0.205 2.370 0.275 ;
        RECT  2.300 0.705 2.370 0.775 ;
        RECT  2.145 0.845 2.345 0.915 ;
        RECT  2.230 0.205 2.300 0.775 ;
        RECT  2.160 0.985 2.280 1.065 ;
        RECT  1.365 0.205 2.230 0.275 ;
        RECT  1.290 0.985 2.160 1.055 ;
        RECT  2.075 0.345 2.145 0.915 ;
        RECT  1.920 0.355 1.990 0.915 ;
        RECT  1.490 0.355 1.920 0.425 ;
        RECT  1.420 0.845 1.920 0.915 ;
        RECT  1.365 0.545 1.570 0.615 ;
        RECT  1.295 0.205 1.365 0.800 ;
        RECT  1.110 0.205 1.295 0.275 ;
        RECT  1.010 0.730 1.295 0.800 ;
        RECT  1.220 0.870 1.290 1.055 ;
        RECT  0.905 0.870 1.220 0.940 ;
        RECT  0.835 0.720 0.905 0.940 ;
        RECT  0.775 0.190 0.845 0.465 ;
        RECT  0.580 0.720 0.835 0.790 ;
        RECT  0.440 0.370 0.775 0.440 ;
        RECT  0.615 0.870 0.685 1.030 ;
        RECT  0.440 0.870 0.615 0.940 ;
        RECT  0.510 0.520 0.580 0.790 ;
        RECT  0.370 0.370 0.440 0.940 ;
        RECT  0.270 0.545 0.370 0.615 ;
    END
END HICIND2BWP

MACRO HICOND1BWP
    CLASS CORE ;
    FOREIGN HICOND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.045 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.735 2.415 1.045 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.0997 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.235 0.735 0.305 1.035 ;
        RECT  0.105 0.735 0.235 0.805 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.035 0.185 0.105 0.805 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.0724 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.995 2.120 1.075 ;
        RECT  0.710 0.995 2.000 1.065 ;
        RECT  0.640 0.880 0.710 1.065 ;
        RECT  0.525 0.880 0.640 0.950 ;
        RECT  0.455 0.520 0.525 0.950 ;
        RECT  0.360 0.520 0.455 0.640 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.345 0.670 0.640 ;
        RECT  0.280 0.345 0.595 0.415 ;
        RECT  0.210 0.345 0.280 0.640 ;
        RECT  0.180 0.520 0.210 0.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.115 2.520 0.115 ;
        RECT  2.180 -0.115 2.300 0.140 ;
        RECT  1.350 -0.115 2.180 0.115 ;
        RECT  1.270 -0.115 1.350 0.280 ;
        RECT  0.980 -0.115 1.270 0.115 ;
        RECT  0.860 -0.115 0.980 0.130 ;
        RECT  0.540 -0.115 0.860 0.115 ;
        RECT  0.460 -0.115 0.540 0.265 ;
        RECT  0.000 -0.115 0.460 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.200 0.735 2.280 1.375 ;
        RECT  1.340 1.145 2.200 1.375 ;
        RECT  1.220 1.135 1.340 1.375 ;
        RECT  0.925 1.145 1.220 1.375 ;
        RECT  0.805 1.135 0.925 1.375 ;
        RECT  0.540 1.145 0.805 1.375 ;
        RECT  0.420 1.020 0.540 1.375 ;
        RECT  0.125 1.145 0.420 1.375 ;
        RECT  0.055 0.920 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.290 0.520 2.340 0.640 ;
        RECT  2.220 0.210 2.290 0.640 ;
        RECT  1.730 0.210 2.220 0.280 ;
        RECT  2.015 0.350 2.085 0.865 ;
        RECT  1.950 0.520 2.015 0.640 ;
        RECT  1.880 0.365 1.930 0.435 ;
        RECT  1.880 0.855 1.930 0.925 ;
        RECT  1.810 0.365 1.880 0.925 ;
        RECT  0.880 0.855 1.810 0.925 ;
        RECT  1.660 0.210 1.730 0.775 ;
        RECT  1.610 0.705 1.660 0.775 ;
        RECT  1.455 0.200 1.525 0.785 ;
        RECT  1.190 0.360 1.455 0.430 ;
        RECT  1.010 0.715 1.455 0.785 ;
        RECT  0.880 0.545 1.350 0.615 ;
        RECT  1.070 0.220 1.190 0.430 ;
        RECT  0.810 0.205 0.880 0.925 ;
        RECT  0.640 0.205 0.810 0.275 ;
        RECT  0.610 0.740 0.810 0.810 ;
    END
END HICOND1BWP

MACRO HICOND2BWP
    CLASS CORE ;
    FOREIGN HICOND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.845 0.355 2.905 0.805 ;
        RECT  2.835 0.185 2.845 1.035 ;
        RECT  2.775 0.185 2.835 0.465 ;
        RECT  2.775 0.735 2.835 1.035 ;
        END
    END S
    PIN CON
        ANTENNADIFFAREA 0.1664 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 0.870 0.710 0.940 ;
        RECT  0.415 0.215 0.530 0.285 ;
        RECT  0.345 0.215 0.415 0.410 ;
        RECT  0.105 0.340 0.345 0.410 ;
        RECT  0.210 0.820 0.285 0.940 ;
        RECT  0.105 0.820 0.210 0.890 ;
        RECT  0.035 0.340 0.105 0.890 ;
        END
    END CON
    PIN CI
        ANTENNAGATEAREA 0.1012 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 0.990 2.480 1.075 ;
        RECT  1.045 0.990 2.340 1.060 ;
        RECT  0.975 0.870 1.045 1.060 ;
        RECT  0.865 0.870 0.975 0.940 ;
        RECT  0.805 0.720 0.865 0.940 ;
        RECT  0.795 0.495 0.805 0.940 ;
        RECT  0.715 0.495 0.795 0.790 ;
        RECT  0.430 0.720 0.715 0.790 ;
        RECT  0.360 0.650 0.430 0.790 ;
        RECT  0.265 0.650 0.360 0.720 ;
        RECT  0.175 0.495 0.265 0.720 ;
        END
    END CI
    PIN A
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.520 0.995 0.645 ;
        RECT  0.875 0.355 0.955 0.645 ;
        RECT  0.635 0.355 0.875 0.425 ;
        RECT  0.565 0.355 0.635 0.630 ;
        RECT  0.500 0.530 0.565 0.630 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.300 ;
        RECT  2.660 -0.115 2.950 0.115 ;
        RECT  2.540 -0.115 2.660 0.135 ;
        RECT  1.260 -0.115 2.540 0.115 ;
        RECT  1.140 -0.115 1.260 0.140 ;
        RECT  0.865 -0.115 1.140 0.115 ;
        RECT  0.795 -0.115 0.865 0.280 ;
        RECT  0.140 -0.115 0.795 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.875 3.030 1.375 ;
        RECT  2.640 1.145 2.950 1.375 ;
        RECT  2.560 0.735 2.640 1.375 ;
        RECT  1.640 1.145 2.560 1.375 ;
        RECT  1.520 1.130 1.640 1.375 ;
        RECT  1.270 1.145 1.520 1.375 ;
        RECT  1.150 1.130 1.270 1.375 ;
        RECT  0.890 1.145 1.150 1.375 ;
        RECT  0.770 1.010 0.890 1.375 ;
        RECT  0.530 1.145 0.770 1.375 ;
        RECT  0.410 1.010 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.970 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.675 0.545 2.760 0.615 ;
        RECT  2.605 0.205 2.675 0.615 ;
        RECT  2.015 0.205 2.605 0.275 ;
        RECT  2.355 0.345 2.425 0.920 ;
        RECT  2.265 0.520 2.355 0.640 ;
        RECT  2.180 0.850 2.250 0.920 ;
        RECT  2.180 0.355 2.240 0.425 ;
        RECT  2.110 0.355 2.180 0.920 ;
        RECT  1.220 0.850 2.110 0.920 ;
        RECT  1.925 0.205 2.015 0.775 ;
        RECT  1.735 0.195 1.805 0.780 ;
        RECT  1.450 0.360 1.735 0.430 ;
        RECT  1.330 0.710 1.735 0.780 ;
        RECT  1.220 0.545 1.620 0.615 ;
        RECT  1.330 0.220 1.450 0.430 ;
        RECT  1.150 0.210 1.220 0.920 ;
        RECT  0.950 0.210 1.150 0.280 ;
        RECT  0.950 0.730 1.150 0.800 ;
    END
END HICOND2BWP

MACRO IAO21D0BWP
    CLASS CORE ;
    FOREIGN IAO21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 1.045 ;
        RECT  0.735 0.355 0.875 0.425 ;
        RECT  0.845 0.915 0.875 1.045 ;
        RECT  0.665 0.185 0.735 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.400 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.820 -0.115 0.940 0.275 ;
        RECT  0.550 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.160 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.160 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.980 1.375 ;
        RECT  0.430 0.990 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.525 0.345 0.595 0.915 ;
        RECT  0.320 0.345 0.525 0.415 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.240 0.185 0.320 0.415 ;
        RECT  0.060 0.845 0.140 1.040 ;
    END
END IAO21D0BWP

MACRO IAO21D1BWP
    CLASS CORE ;
    FOREIGN IAO21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0885 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 1.075 ;
        RECT  0.735 0.355 0.875 0.425 ;
        RECT  0.830 0.835 0.875 1.075 ;
        RECT  0.665 0.245 0.735 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.400 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.820 -0.115 0.940 0.280 ;
        RECT  0.550 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.160 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.160 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.980 1.375 ;
        RECT  0.430 1.000 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.525 0.345 0.595 0.915 ;
        RECT  0.320 0.345 0.525 0.415 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.240 0.185 0.320 0.415 ;
        RECT  0.060 0.845 0.140 1.055 ;
    END
END IAO21D1BWP

MACRO IAO21D2BWP
    CLASS CORE ;
    FOREIGN IAO21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.235 1.025 0.405 ;
        RECT  0.805 0.335 0.955 0.405 ;
        RECT  0.805 0.855 0.870 0.925 ;
        RECT  0.735 0.335 0.805 0.925 ;
        RECT  0.665 0.335 0.735 0.405 ;
        RECT  0.595 0.235 0.665 0.405 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.440 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.265 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.265 ;
        RECT  0.150 -0.115 0.390 0.115 ;
        RECT  0.035 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.145 1.260 1.375 ;
        RECT  1.130 0.970 1.225 1.375 ;
        RECT  0.510 1.145 1.130 1.375 ;
        RECT  0.390 1.030 0.510 1.375 ;
        RECT  0.000 1.145 0.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.065 0.520 1.135 0.900 ;
        RECT  1.060 0.830 1.065 0.900 ;
        RECT  0.990 0.830 1.060 1.065 ;
        RECT  0.660 0.995 0.990 1.065 ;
        RECT  0.590 0.890 0.660 1.065 ;
        RECT  0.525 0.545 0.620 0.615 ;
        RECT  0.525 0.890 0.590 0.960 ;
        RECT  0.455 0.345 0.525 0.960 ;
        RECT  0.305 0.345 0.455 0.415 ;
        RECT  0.130 0.890 0.455 0.960 ;
        RECT  0.235 0.235 0.305 0.415 ;
        RECT  0.050 0.730 0.130 1.030 ;
    END
END IAO21D2BWP

MACRO IAO21D4BWP
    CLASS CORE ;
    FOREIGN IAO21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2884 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.005 0.470 ;
        RECT  1.995 0.775 2.005 0.905 ;
        RECT  1.930 0.185 1.995 0.905 ;
        RECT  1.785 0.355 1.930 0.905 ;
        RECT  1.650 0.355 1.785 0.425 ;
        RECT  1.575 0.775 1.785 0.905 ;
        RECT  1.570 0.195 1.650 0.425 ;
        RECT  1.290 0.355 1.570 0.425 ;
        RECT  1.210 0.195 1.290 0.425 ;
        RECT  0.930 0.355 1.210 0.425 ;
        RECT  0.850 0.265 0.930 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.650 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.185 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.185 0.465 ;
        RECT  1.830 -0.115 2.110 0.115 ;
        RECT  1.750 -0.115 1.830 0.285 ;
        RECT  1.470 -0.115 1.750 0.115 ;
        RECT  1.390 -0.115 1.470 0.285 ;
        RECT  1.110 -0.115 1.390 0.115 ;
        RECT  1.030 -0.115 1.110 0.285 ;
        RECT  0.750 -0.115 1.030 0.115 ;
        RECT  0.675 -0.115 0.750 0.465 ;
        RECT  0.560 -0.115 0.675 0.115 ;
        RECT  0.460 -0.115 0.560 0.275 ;
        RECT  0.200 -0.115 0.460 0.115 ;
        RECT  0.100 -0.115 0.200 0.275 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 1.145 2.240 1.375 ;
        RECT  1.215 0.835 1.285 1.375 ;
        RECT  0.925 1.145 1.215 1.375 ;
        RECT  0.855 0.835 0.925 1.375 ;
        RECT  0.190 1.145 0.855 1.375 ;
        RECT  0.115 0.745 0.190 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.650 0.355 1.715 0.425 ;
        RECT  1.575 0.775 1.715 0.905 ;
        RECT  1.570 0.195 1.650 0.425 ;
        RECT  1.290 0.355 1.570 0.425 ;
        RECT  1.210 0.195 1.290 0.425 ;
        RECT  0.930 0.355 1.210 0.425 ;
        RECT  2.115 0.740 2.185 1.055 ;
        RECT  1.465 0.985 2.115 1.055 ;
        RECT  1.395 0.695 1.465 1.055 ;
        RECT  1.105 0.695 1.395 0.765 ;
        RECT  0.570 0.545 1.290 0.615 ;
        RECT  1.035 0.695 1.105 1.030 ;
        RECT  0.745 0.695 1.035 0.765 ;
        RECT  0.675 0.695 0.745 1.030 ;
        RECT  0.500 0.355 0.570 1.025 ;
        RECT  0.365 0.355 0.500 0.425 ;
        RECT  0.480 0.745 0.500 1.025 ;
        RECT  0.295 0.255 0.365 0.425 ;
        RECT  0.850 0.265 0.930 0.425 ;
    END
END IAO21D4BWP

MACRO IAO22D0BWP
    CLASS CORE ;
    FOREIGN IAO22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.205 0.870 0.275 ;
        RECT  0.735 0.205 0.805 0.775 ;
        RECT  0.665 0.700 0.735 0.775 ;
        RECT  0.595 0.700 0.665 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.625 ;
        RECT  1.040 0.540 1.155 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.260 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.665 -0.115 1.120 0.115 ;
        RECT  0.595 -0.115 0.665 0.280 ;
        RECT  0.485 -0.115 0.595 0.115 ;
        RECT  0.415 -0.115 0.485 0.280 ;
        RECT  0.130 -0.115 0.415 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.260 1.375 ;
        RECT  0.930 0.990 1.050 1.375 ;
        RECT  0.130 1.145 0.930 1.375 ;
        RECT  0.050 0.940 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.845 1.205 1.065 ;
        RECT  0.845 0.845 1.135 0.915 ;
        RECT  0.775 0.845 0.845 1.065 ;
        RECT  0.525 0.540 0.665 0.620 ;
        RECT  0.455 0.355 0.525 1.045 ;
        RECT  0.310 0.355 0.455 0.425 ;
        RECT  0.390 0.975 0.455 1.045 ;
        RECT  0.230 0.185 0.310 0.425 ;
    END
END IAO22D0BWP

MACRO IAO22D1BWP
    CLASS CORE ;
    FOREIGN IAO22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0885 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.185 0.860 0.425 ;
        RECT  0.735 0.185 0.805 0.775 ;
        RECT  0.665 0.700 0.735 0.775 ;
        RECT  0.595 0.700 0.665 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.625 ;
        RECT  1.040 0.545 1.155 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.260 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.665 -0.115 1.120 0.115 ;
        RECT  0.595 -0.115 0.665 0.430 ;
        RECT  0.130 -0.115 0.595 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.260 1.375 ;
        RECT  0.930 0.985 1.050 1.375 ;
        RECT  0.130 1.145 0.930 1.375 ;
        RECT  0.050 0.935 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.845 1.205 0.965 ;
        RECT  0.750 0.845 1.135 0.915 ;
        RECT  0.525 0.540 0.645 0.620 ;
        RECT  0.455 0.345 0.525 1.050 ;
        RECT  0.310 0.345 0.455 0.415 ;
        RECT  0.390 0.980 0.455 1.050 ;
        RECT  0.230 0.185 0.310 0.415 ;
    END
END IAO22D1BWP

MACRO IAO22D2BWP
    CLASS CORE ;
    FOREIGN IAO22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.195 1.085 0.810 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.905 ;
        RECT  1.485 0.495 1.575 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.680 0.115 ;
        RECT  1.160 -0.115 1.280 0.285 ;
        RECT  0.890 -0.115 1.160 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.340 -0.115 0.810 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.985 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 1.030 1.280 1.375 ;
        RECT  0.910 1.145 1.160 1.375 ;
        RECT  0.790 1.025 0.910 1.375 ;
        RECT  0.710 1.145 0.790 1.375 ;
        RECT  0.590 1.025 0.710 1.375 ;
        RECT  0.130 1.145 0.590 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.185 1.640 0.425 ;
        RECT  1.225 0.355 1.540 0.425 ;
        RECT  1.225 0.885 1.470 0.955 ;
        RECT  1.155 0.355 1.225 0.955 ;
        RECT  0.670 0.885 1.155 0.955 ;
        RECT  0.845 0.370 0.915 0.640 ;
        RECT  0.685 0.370 0.845 0.440 ;
        RECT  0.615 0.205 0.685 0.440 ;
        RECT  0.600 0.520 0.670 0.955 ;
        RECT  0.525 0.370 0.615 0.440 ;
        RECT  0.130 0.215 0.530 0.285 ;
        RECT  0.455 0.370 0.525 0.990 ;
        RECT  0.420 0.750 0.455 0.990 ;
        RECT  0.050 0.215 0.130 0.385 ;
    END
END IAO22D2BWP

MACRO IAO22D4BWP
    CLASS CORE ;
    FOREIGN IAO22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.920 0.465 ;
        RECT  1.855 0.700 1.920 0.820 ;
        RECT  1.850 0.185 1.855 0.820 ;
        RECT  1.645 0.350 1.850 0.820 ;
        RECT  1.575 0.350 1.645 0.465 ;
        RECT  1.480 0.700 1.645 0.820 ;
        RECT  1.495 0.185 1.575 0.465 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.485 0.905 ;
        RECT  2.325 0.495 2.415 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.225 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.805 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.270 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.115 2.520 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.750 -0.115 2.010 0.115 ;
        RECT  1.670 -0.115 1.750 0.280 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.300 ;
        RECT  0.670 -0.115 1.310 0.115 ;
        RECT  0.590 -0.115 0.670 0.285 ;
        RECT  0.310 -0.115 0.590 0.115 ;
        RECT  0.230 -0.115 0.310 0.285 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.985 2.480 1.375 ;
        RECT  2.130 1.145 2.380 1.375 ;
        RECT  2.010 1.030 2.130 1.375 ;
        RECT  1.770 1.145 2.010 1.375 ;
        RECT  1.650 1.030 1.770 1.375 ;
        RECT  1.410 1.145 1.650 1.375 ;
        RECT  1.290 1.030 1.410 1.375 ;
        RECT  1.030 1.145 1.290 1.375 ;
        RECT  0.950 0.975 1.030 1.375 ;
        RECT  0.310 1.145 0.950 1.375 ;
        RECT  0.230 0.835 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.495 0.185 1.575 0.465 ;
        RECT  1.480 0.700 1.575 0.820 ;
        RECT  2.380 0.185 2.480 0.425 ;
        RECT  2.060 0.355 2.380 0.425 ;
        RECT  2.210 0.890 2.290 1.040 ;
        RECT  2.060 0.890 2.210 0.960 ;
        RECT  1.990 0.355 2.060 0.960 ;
        RECT  1.380 0.890 1.990 0.960 ;
        RECT  1.375 0.540 1.540 0.610 ;
        RECT  1.310 0.680 1.380 0.960 ;
        RECT  1.305 0.370 1.375 0.610 ;
        RECT  1.225 0.680 1.310 0.750 ;
        RECT  1.025 0.370 1.305 0.440 ;
        RECT  0.850 0.215 1.230 0.285 ;
        RECT  1.155 0.520 1.225 0.750 ;
        RECT  1.120 0.835 1.220 1.075 ;
        RECT  1.025 0.835 1.120 0.905 ;
        RECT  0.955 0.370 1.025 0.905 ;
        RECT  0.680 0.835 0.955 0.905 ;
        RECT  0.490 0.695 0.870 0.765 ;
        RECT  0.770 0.215 0.850 0.425 ;
        RECT  0.130 0.355 0.770 0.425 ;
        RECT  0.580 0.835 0.680 1.075 ;
        RECT  0.410 0.695 0.490 1.025 ;
        RECT  0.130 0.695 0.410 0.765 ;
        RECT  0.050 0.265 0.130 0.425 ;
        RECT  0.050 0.695 0.130 1.025 ;
    END
END IAO22D4BWP

MACRO IIND4D0BWP
    CLASS CORE ;
    FOREIGN IIND4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0827 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.185 1.130 0.275 ;
        RECT  0.875 0.185 0.945 1.045 ;
        RECT  0.845 0.855 0.875 1.045 ;
        RECT  0.535 0.855 0.845 0.925 ;
        RECT  0.455 0.855 0.535 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.620 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.520 1.435 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 -0.115 1.540 0.115 ;
        RECT  1.380 -0.115 1.480 0.275 ;
        RECT  0.340 -0.115 1.380 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.145 1.540 1.375 ;
        RECT  1.390 0.920 1.470 1.375 ;
        RECT  1.110 1.145 1.390 1.375 ;
        RECT  1.030 0.920 1.110 1.375 ;
        RECT  0.740 1.145 1.030 1.375 ;
        RECT  0.620 0.995 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.045 ;
        RECT  1.015 0.540 1.210 0.620 ;
        RECT  0.315 0.345 0.385 0.925 ;
        RECT  0.125 0.345 0.315 0.415 ;
        RECT  0.125 0.855 0.315 0.925 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.855 0.125 1.045 ;
    END
END IIND4D0BWP

MACRO IIND4D1BWP
    CLASS CORE ;
    FOREIGN IIND4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1653 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.100 0.445 ;
        RECT  0.945 0.355 1.015 0.445 ;
        RECT  0.875 0.355 0.945 0.915 ;
        RECT  0.525 0.845 0.875 0.915 ;
        RECT  0.455 0.745 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.495 1.435 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 -0.115 1.540 0.115 ;
        RECT  1.380 -0.115 1.480 0.275 ;
        RECT  0.340 -0.115 1.380 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.145 1.540 1.375 ;
        RECT  1.390 0.930 1.470 1.375 ;
        RECT  1.110 1.145 1.390 1.375 ;
        RECT  1.030 0.840 1.110 1.375 ;
        RECT  0.740 1.145 1.030 1.375 ;
        RECT  0.620 0.995 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.055 ;
        RECT  1.015 0.540 1.210 0.620 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.195 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END IIND4D1BWP

MACRO IIND4D2BWP
    CLASS CORE ;
    FOREIGN IIND4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2730 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.720 2.170 0.790 ;
        RECT  0.875 0.355 0.945 0.790 ;
        RECT  0.790 0.355 0.875 0.455 ;
        RECT  0.790 0.720 0.875 0.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.810 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.225 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.415 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.150 -0.115 2.380 0.115 ;
        RECT  2.070 -0.115 2.150 0.305 ;
        RECT  0.315 -0.115 2.070 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.145 2.380 1.375 ;
        RECT  2.240 1.000 2.340 1.375 ;
        RECT  1.965 1.145 2.240 1.375 ;
        RECT  1.895 1.000 1.965 1.375 ;
        RECT  1.620 1.145 1.895 1.375 ;
        RECT  1.520 1.000 1.620 1.375 ;
        RECT  1.425 1.145 1.520 1.375 ;
        RECT  1.355 1.000 1.425 1.375 ;
        RECT  1.065 1.145 1.355 1.375 ;
        RECT  0.995 1.000 1.065 1.375 ;
        RECT  0.705 1.145 0.995 1.375 ;
        RECT  0.635 1.000 0.705 1.375 ;
        RECT  0.315 1.145 0.635 1.375 ;
        RECT  0.245 1.000 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.255 0.205 2.325 0.465 ;
        RECT  2.250 0.545 2.320 0.930 ;
        RECT  1.965 0.395 2.255 0.465 ;
        RECT  2.050 0.545 2.250 0.615 ;
        RECT  0.140 0.860 2.250 0.930 ;
        RECT  1.895 0.205 1.965 0.465 ;
        RECT  1.620 0.205 1.895 0.285 ;
        RECT  1.150 0.355 1.815 0.425 ;
        RECT  1.510 0.185 1.620 0.285 ;
        RECT  1.340 0.185 1.440 0.285 ;
        RECT  0.710 0.205 1.340 0.285 ;
        RECT  0.555 0.545 0.805 0.615 ;
        RECT  0.640 0.205 0.710 0.465 ;
        RECT  0.485 0.195 0.555 0.790 ;
        RECT  0.410 0.195 0.485 0.275 ;
        RECT  0.410 0.720 0.485 0.790 ;
        RECT  0.105 0.860 0.140 0.960 ;
        RECT  0.105 0.195 0.130 0.315 ;
        RECT  0.035 0.195 0.105 0.960 ;
    END
END IIND4D2BWP

MACRO IIND4D4BWP
    CLASS CORE ;
    FOREIGN IIND4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.345 3.965 0.465 ;
        RECT  3.955 0.700 3.965 1.035 ;
        RECT  3.895 0.345 3.955 1.035 ;
        RECT  3.745 0.345 3.895 0.820 ;
        RECT  3.510 0.345 3.745 0.465 ;
        RECT  3.605 0.700 3.745 0.820 ;
        RECT  3.535 0.700 3.605 1.035 ;
        RECT  3.080 0.835 3.535 0.905 ;
        RECT  2.980 0.835 3.080 1.075 ;
        RECT  2.720 0.835 2.980 0.905 ;
        RECT  2.620 0.835 2.720 1.075 ;
        RECT  2.360 0.835 2.620 0.905 ;
        RECT  2.260 0.835 2.360 1.075 ;
        RECT  2.000 0.835 2.260 0.905 ;
        RECT  1.900 0.835 2.000 1.075 ;
        RECT  1.460 0.835 1.900 0.905 ;
        RECT  1.360 0.835 1.460 1.075 ;
        RECT  1.100 0.835 1.360 0.905 ;
        RECT  1.000 0.835 1.100 1.075 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.495 2.350 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.535 0.495 0.620 0.640 ;
        RECT  0.455 0.495 0.535 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.535 0.230 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 4.200 0.115 ;
        RECT  1.550 -0.115 1.630 0.280 ;
        RECT  1.270 -0.115 1.550 0.115 ;
        RECT  1.190 -0.115 1.270 0.280 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.830 -0.115 0.910 0.455 ;
        RECT  0.550 -0.115 0.830 0.115 ;
        RECT  0.470 -0.115 0.550 0.415 ;
        RECT  0.190 -0.115 0.470 0.115 ;
        RECT  0.110 -0.115 0.190 0.285 ;
        RECT  0.000 -0.115 0.110 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.680 4.150 1.375 ;
        RECT  3.790 1.145 4.070 1.375 ;
        RECT  3.710 0.890 3.790 1.375 ;
        RECT  3.430 1.145 3.710 1.375 ;
        RECT  3.350 0.975 3.430 1.375 ;
        RECT  3.250 1.145 3.350 1.375 ;
        RECT  3.170 0.975 3.250 1.375 ;
        RECT  2.890 1.145 3.170 1.375 ;
        RECT  2.810 0.975 2.890 1.375 ;
        RECT  2.530 1.145 2.810 1.375 ;
        RECT  2.450 0.975 2.530 1.375 ;
        RECT  2.170 1.145 2.450 1.375 ;
        RECT  2.090 0.975 2.170 1.375 ;
        RECT  1.810 1.145 2.090 1.375 ;
        RECT  1.730 0.975 1.810 1.375 ;
        RECT  1.630 1.145 1.730 1.375 ;
        RECT  1.550 0.975 1.630 1.375 ;
        RECT  1.270 1.145 1.550 1.375 ;
        RECT  1.190 0.975 1.270 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 1.010 0.930 1.375 ;
        RECT  0.570 1.145 0.810 1.375 ;
        RECT  0.450 1.010 0.570 1.375 ;
        RECT  0.200 1.145 0.450 1.375 ;
        RECT  0.100 0.700 0.200 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.510 0.345 3.675 0.465 ;
        RECT  3.605 0.700 3.675 0.820 ;
        RECT  3.535 0.700 3.605 1.035 ;
        RECT  3.080 0.835 3.535 0.905 ;
        RECT  2.980 0.835 3.080 1.075 ;
        RECT  2.720 0.835 2.980 0.905 ;
        RECT  2.620 0.835 2.720 1.075 ;
        RECT  2.360 0.835 2.620 0.905 ;
        RECT  2.260 0.835 2.360 1.075 ;
        RECT  2.000 0.835 2.260 0.905 ;
        RECT  1.900 0.835 2.000 1.075 ;
        RECT  1.460 0.835 1.900 0.905 ;
        RECT  1.360 0.835 1.460 1.075 ;
        RECT  1.100 0.835 1.360 0.905 ;
        RECT  1.000 0.835 1.100 1.075 ;
        RECT  4.070 0.205 4.150 0.485 ;
        RECT  3.430 0.205 4.070 0.275 ;
        RECT  3.340 0.545 3.655 0.615 ;
        RECT  3.350 0.205 3.430 0.460 ;
        RECT  2.610 0.205 3.350 0.275 ;
        RECT  3.270 0.545 3.340 0.765 ;
        RECT  2.530 0.345 3.270 0.415 ;
        RECT  0.900 0.695 3.270 0.765 ;
        RECT  2.450 0.205 2.530 0.415 ;
        RECT  1.710 0.205 2.450 0.275 ;
        RECT  1.445 0.350 2.370 0.420 ;
        RECT  0.760 0.545 1.510 0.615 ;
        RECT  1.375 0.185 1.445 0.420 ;
        RECT  1.085 0.350 1.375 0.420 ;
        RECT  1.015 0.185 1.085 0.450 ;
        RECT  0.830 0.695 0.900 0.940 ;
        RECT  0.370 0.870 0.830 0.940 ;
        RECT  0.690 0.185 0.760 0.790 ;
        RECT  0.640 0.185 0.690 0.425 ;
        RECT  0.630 0.720 0.690 0.790 ;
        RECT  0.300 0.190 0.370 1.070 ;
    END
END IIND4D4BWP

MACRO IINR4D0BWP
    CLASS CORE ;
    FOREIGN IINR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0967 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.185 1.085 0.425 ;
        RECT  0.685 0.355 0.980 0.425 ;
        RECT  0.615 0.185 0.685 0.425 ;
        RECT  0.530 0.355 0.615 0.425 ;
        RECT  0.455 0.355 0.530 1.065 ;
        RECT  0.410 0.985 0.455 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.110 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.355 1.365 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.115 1.540 0.115 ;
        RECT  1.170 -0.115 1.270 0.285 ;
        RECT  0.870 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.870 0.285 ;
        RECT  0.510 -0.115 0.790 0.115 ;
        RECT  0.430 -0.115 0.510 0.280 ;
        RECT  0.320 -0.115 0.430 0.115 ;
        RECT  0.220 -0.115 0.320 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.160 1.115 1.280 1.375 ;
        RECT  0.320 1.145 1.160 1.375 ;
        RECT  0.220 0.985 0.320 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.470 0.205 1.505 0.795 ;
        RECT  1.435 0.205 1.470 1.045 ;
        RECT  1.370 0.205 1.435 0.285 ;
        RECT  1.390 0.715 1.435 1.045 ;
        RECT  0.760 0.975 1.390 1.045 ;
        RECT  0.680 0.520 0.760 1.045 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.125 0.345 0.315 0.415 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.015 ;
    END
END IINR4D0BWP

MACRO IINR4D1BWP
    CLASS CORE ;
    FOREIGN IINR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1287 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.345 1.430 0.415 ;
        RECT  1.085 0.845 1.250 0.915 ;
        RECT  1.015 0.345 1.085 0.915 ;
        RECT  0.230 0.345 1.015 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.230 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.355 1.925 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.445 2.065 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.240 0.115 ;
        RECT  1.880 -0.115 2.000 0.280 ;
        RECT  1.580 -0.115 1.880 0.115 ;
        RECT  1.510 -0.115 1.580 0.460 ;
        RECT  1.210 -0.115 1.510 0.115 ;
        RECT  1.090 -0.115 1.210 0.275 ;
        RECT  0.570 -0.115 1.090 0.115 ;
        RECT  0.450 -0.115 0.570 0.275 ;
        RECT  0.150 -0.115 0.450 0.115 ;
        RECT  0.070 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 1.145 2.240 1.375 ;
        RECT  1.900 0.990 1.980 1.375 ;
        RECT  0.530 1.145 1.900 1.375 ;
        RECT  0.410 0.975 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.135 0.200 2.205 0.980 ;
        RECT  2.115 0.200 2.135 0.320 ;
        RECT  2.115 0.845 2.135 0.980 ;
        RECT  1.425 0.845 2.115 0.915 ;
        RECT  1.720 0.220 1.790 0.290 ;
        RECT  1.720 0.705 1.790 0.775 ;
        RECT  1.650 0.220 1.720 0.775 ;
        RECT  1.515 0.540 1.650 0.620 ;
        RECT  0.865 0.985 1.610 1.055 ;
        RECT  1.355 0.540 1.425 0.915 ;
        RECT  1.170 0.540 1.355 0.620 ;
        RECT  0.785 0.835 0.865 1.055 ;
        RECT  0.150 0.835 0.785 0.905 ;
        RECT  0.070 0.735 0.150 1.035 ;
    END
END IINR4D1BWP

MACRO IINR4D2BWP
    CLASS CORE ;
    FOREIGN IINR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3094 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.575 0.615 2.665 1.065 ;
        RECT  2.305 0.615 2.575 0.705 ;
        RECT  2.205 0.215 2.485 0.335 ;
        RECT  2.235 0.615 2.305 0.905 ;
        RECT  2.205 0.615 2.235 0.705 ;
        RECT  2.135 0.215 2.205 0.705 ;
        RECT  0.595 0.215 2.135 0.335 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.450 0.805 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.450 1.365 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.355 3.045 0.640 ;
        RECT  2.890 0.520 2.975 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 -0.115 3.080 0.115 ;
        RECT  2.940 -0.115 3.040 0.275 ;
        RECT  2.670 -0.115 2.940 0.115 ;
        RECT  2.590 -0.115 2.670 0.295 ;
        RECT  0.510 -0.115 2.590 0.115 ;
        RECT  0.430 -0.115 0.510 0.295 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.295 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.145 3.080 1.375 ;
        RECT  2.940 0.720 3.040 1.375 ;
        RECT  0.890 1.145 2.940 1.375 ;
        RECT  0.770 0.985 0.890 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.430 0.950 0.510 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.950 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.820 0.195 2.870 0.265 ;
        RECT  2.820 0.760 2.850 1.045 ;
        RECT  2.750 0.195 2.820 1.045 ;
        RECT  2.285 0.450 2.750 0.520 ;
        RECT  2.410 0.775 2.490 1.055 ;
        RECT  2.125 0.985 2.410 1.055 ;
        RECT  2.055 0.775 2.125 1.055 ;
        RECT  1.670 0.985 2.055 1.055 ;
        RECT  1.875 0.615 1.945 0.915 ;
        RECT  1.670 0.450 1.910 0.520 ;
        RECT  1.590 0.845 1.875 0.915 ;
        RECT  1.600 0.450 1.670 0.775 ;
        RECT  0.330 0.705 1.600 0.775 ;
        RECT  1.510 0.845 1.590 1.055 ;
        RECT  1.130 0.985 1.510 1.055 ;
        RECT  0.590 0.845 1.430 0.915 ;
        RECT  0.260 0.185 0.330 1.075 ;
    END
END IINR4D2BWP

MACRO IINR4D4BWP
    CLASS CORE ;
    FOREIGN IINR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5756 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.205 5.090 0.325 ;
        RECT  5.010 0.635 5.090 0.915 ;
        RECT  4.730 0.635 5.010 0.740 ;
        RECT  4.650 0.635 4.730 0.915 ;
        RECT  4.515 0.635 4.650 0.740 ;
        RECT  4.365 0.205 4.515 0.740 ;
        RECT  4.305 0.205 4.365 0.915 ;
        RECT  0.790 0.205 4.305 0.325 ;
        RECT  4.295 0.635 4.305 0.915 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.445 1.535 0.515 ;
        RECT  0.735 0.445 0.945 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.445 2.485 0.515 ;
        RECT  1.855 0.445 2.065 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.600 0.495 5.845 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.115 5.880 0.115 ;
        RECT  5.540 -0.115 5.660 0.275 ;
        RECT  5.270 -0.115 5.540 0.115 ;
        RECT  5.190 -0.115 5.270 0.320 ;
        RECT  0.690 -0.115 5.190 0.115 ;
        RECT  0.610 -0.115 0.690 0.320 ;
        RECT  0.510 -0.115 0.610 0.115 ;
        RECT  0.430 -0.115 0.510 0.425 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.425 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.640 1.145 5.880 1.375 ;
        RECT  5.560 0.835 5.640 1.375 ;
        RECT  1.610 1.145 5.560 1.375 ;
        RECT  1.490 0.985 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 0.985 1.250 1.375 ;
        RECT  0.890 1.145 1.130 1.375 ;
        RECT  0.770 0.985 0.890 1.375 ;
        RECT  0.510 1.145 0.770 1.375 ;
        RECT  0.430 0.845 0.510 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.835 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.205 5.090 0.325 ;
        RECT  5.010 0.635 5.090 0.915 ;
        RECT  4.730 0.635 5.010 0.740 ;
        RECT  4.650 0.635 4.730 0.915 ;
        RECT  4.585 0.635 4.650 0.740 ;
        RECT  0.790 0.205 4.235 0.325 ;
        RECT  5.750 0.190 5.830 0.415 ;
        RECT  5.750 0.695 5.830 1.030 ;
        RECT  5.450 0.345 5.750 0.415 ;
        RECT  5.450 0.695 5.750 0.765 ;
        RECT  5.370 0.190 5.450 1.030 ;
        RECT  4.685 0.445 5.370 0.515 ;
        RECT  5.190 0.610 5.270 1.065 ;
        RECT  4.910 0.995 5.190 1.065 ;
        RECT  4.830 0.810 4.910 1.065 ;
        RECT  4.545 0.995 4.830 1.065 ;
        RECT  4.475 0.810 4.545 1.065 ;
        RECT  4.185 0.995 4.475 1.065 ;
        RECT  4.115 0.625 4.185 1.065 ;
        RECT  3.830 0.995 4.115 1.065 ;
        RECT  3.930 0.615 4.010 0.905 ;
        RECT  2.690 0.445 4.000 0.515 ;
        RECT  3.650 0.615 3.930 0.685 ;
        RECT  3.750 0.765 3.830 1.065 ;
        RECT  3.470 0.995 3.750 1.065 ;
        RECT  3.570 0.615 3.650 0.905 ;
        RECT  3.290 0.615 3.570 0.685 ;
        RECT  3.390 0.765 3.470 1.065 ;
        RECT  3.110 0.995 3.390 1.065 ;
        RECT  3.210 0.615 3.290 0.905 ;
        RECT  2.840 0.615 3.210 0.685 ;
        RECT  3.030 0.765 3.110 1.065 ;
        RECT  1.770 0.985 2.870 1.055 ;
        RECT  2.770 0.615 2.840 0.915 ;
        RECT  1.850 0.845 2.770 0.915 ;
        RECT  2.620 0.445 2.690 0.775 ;
        RECT  0.330 0.705 2.620 0.775 ;
        RECT  1.690 0.845 1.770 1.055 ;
        RECT  1.410 0.845 1.690 0.915 ;
        RECT  1.330 0.845 1.410 1.075 ;
        RECT  1.050 0.845 1.330 0.915 ;
        RECT  0.970 0.845 1.050 1.075 ;
        RECT  0.690 0.845 0.970 0.915 ;
        RECT  0.610 0.845 0.690 1.045 ;
        RECT  0.260 0.190 0.330 1.070 ;
    END
END IINR4D4BWP

MACRO IND2D0BWP
    CLASS CORE ;
    FOREIGN IND2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0551 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 0.845 ;
        RECT  0.630 0.215 0.735 0.285 ;
        RECT  0.550 0.775 0.735 0.845 ;
        RECT  0.470 0.775 0.550 1.065 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.665 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.115 0.840 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.640 0.985 0.740 1.375 ;
        RECT  0.350 1.145 0.640 1.375 ;
        RECT  0.250 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.390 0.545 0.460 0.615 ;
        RECT  0.320 0.345 0.390 0.915 ;
        RECT  0.130 0.345 0.320 0.415 ;
        RECT  0.130 0.845 0.320 0.915 ;
        RECT  0.055 0.185 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.065 ;
    END
END IND2D0BWP

MACRO IND2D1BWP
    CLASS CORE ;
    FOREIGN IND2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1101 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 0.780 ;
        RECT  0.630 0.215 0.735 0.285 ;
        RECT  0.550 0.710 0.735 0.780 ;
        RECT  0.470 0.710 0.550 1.040 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.665 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.115 0.840 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.640 0.985 0.740 1.375 ;
        RECT  0.350 1.145 0.640 1.375 ;
        RECT  0.250 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.390 0.545 0.460 0.615 ;
        RECT  0.320 0.345 0.390 0.915 ;
        RECT  0.130 0.345 0.320 0.415 ;
        RECT  0.130 0.845 0.320 0.915 ;
        RECT  0.055 0.185 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.070 ;
    END
END IND2D1BWP

MACRO IND2D2BWP
    CLASS CORE ;
    FOREIGN IND2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1582 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 0.775 0.865 1.065 ;
        RECT  0.790 0.775 0.795 0.920 ;
        RECT  0.720 0.345 0.790 0.920 ;
        RECT  0.590 0.345 0.720 0.415 ;
        RECT  0.525 0.850 0.720 0.920 ;
        RECT  0.435 0.850 0.525 1.065 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.495 1.085 0.625 ;
        RECT  0.860 0.205 0.930 0.625 ;
        RECT  0.480 0.205 0.860 0.275 ;
        RECT  0.410 0.205 0.480 0.640 ;
        RECT  0.370 0.520 0.410 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.355 0.265 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.115 1.120 0.115 ;
        RECT  1.000 -0.115 1.070 0.350 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.250 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.120 1.375 ;
        RECT  0.970 0.705 1.050 1.375 ;
        RECT  0.700 1.145 0.970 1.375 ;
        RECT  0.600 0.990 0.700 1.375 ;
        RECT  0.330 1.145 0.600 1.375 ;
        RECT  0.250 0.850 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.520 0.650 0.780 ;
        RECT  0.120 0.710 0.560 0.780 ;
        RECT  0.105 0.205 0.170 0.285 ;
        RECT  0.105 0.710 0.120 1.035 ;
        RECT  0.035 0.205 0.105 1.035 ;
    END
END IND2D2BWP

MACRO IND2D4BWP
    CLASS CORE ;
    FOREIGN IND2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3164 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.915 0.345 1.995 1.065 ;
        RECT  1.785 0.345 1.915 0.785 ;
        RECT  1.530 0.345 1.785 0.425 ;
        RECT  1.625 0.695 1.785 0.785 ;
        RECT  1.555 0.695 1.625 1.015 ;
        RECT  1.265 0.695 1.555 0.785 ;
        RECT  1.195 0.695 1.265 1.015 ;
        RECT  0.905 0.695 1.195 0.785 ;
        RECT  0.835 0.695 0.905 1.015 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.650 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.115 2.240 0.115 ;
        RECT  1.190 -0.115 1.270 0.285 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.830 -0.115 0.910 0.285 ;
        RECT  0.510 -0.115 0.830 0.115 ;
        RECT  0.430 -0.115 0.510 0.465 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.425 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.145 2.240 1.375 ;
        RECT  2.090 0.685 2.170 1.375 ;
        RECT  1.810 1.145 2.090 1.375 ;
        RECT  1.730 0.855 1.810 1.375 ;
        RECT  1.450 1.145 1.730 1.375 ;
        RECT  1.370 0.855 1.450 1.375 ;
        RECT  1.090 1.145 1.370 1.375 ;
        RECT  1.010 0.855 1.090 1.375 ;
        RECT  0.730 1.145 1.010 1.375 ;
        RECT  0.650 0.685 0.730 1.375 ;
        RECT  0.510 1.145 0.650 1.375 ;
        RECT  0.430 0.685 0.510 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.345 1.715 0.425 ;
        RECT  1.625 0.695 1.715 0.785 ;
        RECT  1.555 0.695 1.625 1.015 ;
        RECT  1.265 0.695 1.555 0.785 ;
        RECT  1.195 0.695 1.265 1.015 ;
        RECT  0.905 0.695 1.195 0.785 ;
        RECT  0.835 0.695 0.905 1.015 ;
        RECT  2.090 0.205 2.165 0.465 ;
        RECT  1.450 0.205 2.090 0.275 ;
        RECT  1.370 0.205 1.450 0.425 ;
        RECT  1.090 0.355 1.370 0.425 ;
        RECT  0.330 0.545 1.195 0.615 ;
        RECT  1.010 0.190 1.090 0.425 ;
        RECT  0.740 0.355 1.010 0.425 ;
        RECT  0.640 0.185 0.740 0.425 ;
        RECT  0.260 0.185 0.330 1.065 ;
    END
END IND2D4BWP

MACRO IND3D0BWP
    CLASS CORE ;
    FOREIGN IND3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0755 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.215 0.945 0.920 ;
        RECT  0.875 0.215 0.910 1.045 ;
        RECT  0.810 0.215 0.875 0.290 ;
        RECT  0.830 0.850 0.875 1.045 ;
        RECT  0.540 0.850 0.830 0.920 ;
        RECT  0.455 0.850 0.540 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.640 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.115 0.980 0.115 ;
        RECT  0.240 -0.115 0.360 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.145 0.980 1.375 ;
        RECT  0.630 0.990 0.750 1.375 ;
        RECT  0.360 1.145 0.630 1.375 ;
        RECT  0.240 0.990 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.125 0.345 0.315 0.415 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.045 ;
    END
END IND3D0BWP

MACRO IND3D1BWP
    CLASS CORE ;
    FOREIGN IND3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1510 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.195 0.945 0.425 ;
        RECT  0.835 0.845 0.905 1.045 ;
        RECT  0.520 0.195 0.840 0.265 ;
        RECT  0.545 0.845 0.835 0.915 ;
        RECT  0.520 0.740 0.545 1.045 ;
        RECT  0.450 0.195 0.520 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.765 ;
        RECT  0.740 0.545 0.855 0.615 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.345 0.665 0.660 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 -0.115 0.980 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.145 0.980 1.375 ;
        RECT  0.630 1.020 0.750 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.260 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.310 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.310 0.415 ;
        RECT  0.130 0.845 0.310 0.915 ;
        RECT  0.050 0.195 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.065 ;
    END
END IND3D1BWP

MACRO IND3D2BWP
    CLASS CORE ;
    FOREIGN IND3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2156 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.345 1.440 0.415 ;
        RECT  1.340 0.700 1.420 1.055 ;
        RECT  1.225 0.700 1.340 0.780 ;
        RECT  1.155 0.345 1.225 0.780 ;
        RECT  1.060 0.700 1.155 0.780 ;
        RECT  0.980 0.700 1.060 1.055 ;
        RECT  0.525 0.700 0.980 0.780 ;
        RECT  0.445 0.700 0.525 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.645 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.980 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.200 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.620 -0.115 0.700 0.265 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.145 1.680 1.375 ;
        RECT  1.520 0.700 1.600 1.375 ;
        RECT  1.250 1.145 1.520 1.375 ;
        RECT  1.150 0.860 1.250 1.375 ;
        RECT  0.880 1.145 1.150 1.375 ;
        RECT  0.800 0.850 0.880 1.375 ;
        RECT  0.700 1.145 0.800 1.375 ;
        RECT  0.620 0.850 0.700 1.375 ;
        RECT  0.360 1.145 0.620 1.375 ;
        RECT  0.240 0.985 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.520 0.195 1.600 0.385 ;
        RECT  0.780 0.195 1.520 0.265 ;
        RECT  0.530 0.335 1.080 0.425 ;
        RECT  0.340 0.545 0.550 0.615 ;
        RECT  0.430 0.185 0.530 0.425 ;
        RECT  0.270 0.355 0.340 0.915 ;
        RECT  0.170 0.355 0.270 0.425 ;
        RECT  0.160 0.845 0.270 0.915 ;
        RECT  0.070 0.185 0.170 0.425 ;
        RECT  0.080 0.845 0.160 0.985 ;
    END
END IND3D2BWP

MACRO IND3D4BWP
    CLASS CORE ;
    FOREIGN IND3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4312 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.345 2.730 0.465 ;
        RECT  2.635 0.695 2.705 1.035 ;
        RECT  2.415 0.695 2.635 0.800 ;
        RECT  2.345 0.345 2.415 0.800 ;
        RECT  2.275 0.345 2.345 1.035 ;
        RECT  2.205 0.345 2.275 0.800 ;
        RECT  1.985 0.695 2.205 0.800 ;
        RECT  1.915 0.695 1.985 1.035 ;
        RECT  1.625 0.695 1.915 0.800 ;
        RECT  1.555 0.695 1.625 1.035 ;
        RECT  1.085 0.695 1.555 0.800 ;
        RECT  1.015 0.695 1.085 1.035 ;
        RECT  0.725 0.695 1.015 0.800 ;
        RECT  0.655 0.695 0.725 1.035 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.815 0.355 2.905 0.625 ;
        RECT  2.505 0.545 2.815 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 0.495 2.015 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.200 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.115 2.940 0.115 ;
        RECT  1.190 -0.115 1.270 0.285 ;
        RECT  0.905 -0.115 1.190 0.115 ;
        RECT  0.835 -0.115 0.905 0.285 ;
        RECT  0.550 -0.115 0.835 0.115 ;
        RECT  0.470 -0.115 0.550 0.465 ;
        RECT  0.190 -0.115 0.470 0.115 ;
        RECT  0.110 -0.115 0.190 0.425 ;
        RECT  0.000 -0.115 0.110 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.715 2.900 1.375 ;
        RECT  2.540 1.145 2.800 1.375 ;
        RECT  2.440 0.870 2.540 1.375 ;
        RECT  2.180 1.145 2.440 1.375 ;
        RECT  2.080 0.870 2.180 1.375 ;
        RECT  1.820 1.145 2.080 1.375 ;
        RECT  1.720 0.870 1.820 1.375 ;
        RECT  1.460 1.145 1.720 1.375 ;
        RECT  1.360 0.870 1.460 1.375 ;
        RECT  1.280 1.145 1.360 1.375 ;
        RECT  1.180 0.870 1.280 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.820 0.870 0.920 1.375 ;
        RECT  0.550 1.145 0.820 1.375 ;
        RECT  0.470 0.700 0.550 1.375 ;
        RECT  0.190 1.145 0.470 1.375 ;
        RECT  0.110 0.835 0.190 1.375 ;
        RECT  0.000 1.145 0.110 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.345 2.730 0.465 ;
        RECT  2.635 0.695 2.705 1.035 ;
        RECT  2.485 0.695 2.635 0.800 ;
        RECT  1.985 0.695 2.135 0.800 ;
        RECT  1.915 0.695 1.985 1.035 ;
        RECT  1.625 0.695 1.915 0.800 ;
        RECT  1.555 0.695 1.625 1.035 ;
        RECT  1.085 0.695 1.555 0.800 ;
        RECT  1.015 0.695 1.085 1.035 ;
        RECT  0.725 0.695 1.015 0.800 ;
        RECT  0.655 0.695 0.725 1.035 ;
        RECT  2.800 0.185 2.900 0.285 ;
        RECT  1.350 0.205 2.800 0.275 ;
        RECT  1.085 0.355 2.010 0.425 ;
        RECT  0.370 0.545 1.120 0.615 ;
        RECT  1.015 0.185 1.085 0.425 ;
        RECT  0.740 0.355 1.015 0.425 ;
        RECT  0.640 0.185 0.740 0.425 ;
        RECT  0.290 0.185 0.370 1.075 ;
    END
END IND3D4BWP

MACRO IND4D0BWP
    CLASS CORE ;
    FOREIGN IND4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0775 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.200 1.085 0.840 ;
        RECT  0.950 0.200 1.015 0.275 ;
        RECT  0.865 0.770 1.015 0.840 ;
        RECT  0.795 0.770 0.865 1.060 ;
        RECT  0.525 0.770 0.795 0.840 ;
        RECT  0.440 0.770 0.525 1.060 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.670 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.215 0.805 0.485 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 1.120 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.120 1.375 ;
        RECT  0.970 0.920 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.920 0.690 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.345 0.370 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.060 ;
    END
END IND4D0BWP

MACRO IND4D1BWP
    CLASS CORE ;
    FOREIGN IND4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1551 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.195 1.085 0.855 ;
        RECT  0.950 0.195 1.015 0.275 ;
        RECT  0.870 0.775 1.015 0.855 ;
        RECT  0.790 0.775 0.870 1.055 ;
        RECT  0.525 0.775 0.790 0.855 ;
        RECT  0.440 0.775 0.525 1.055 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.670 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 0.640 ;
        RECT  0.705 0.520 0.735 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 -0.115 1.120 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.120 1.375 ;
        RECT  0.970 0.935 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.935 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.985 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.345 0.370 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.075 ;
    END
END IND4D1BWP

MACRO IND4D2BWP
    CLASS CORE ;
    FOREIGN IND4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.185 2.205 0.905 ;
        RECT  2.100 0.185 2.135 0.425 ;
        RECT  2.005 0.835 2.135 0.905 ;
        RECT  1.730 0.355 2.100 0.425 ;
        RECT  1.935 0.835 2.005 1.075 ;
        RECT  1.425 0.835 1.935 0.905 ;
        RECT  1.355 0.835 1.425 1.075 ;
        RECT  1.065 0.835 1.355 0.905 ;
        RECT  0.995 0.835 1.065 1.075 ;
        RECT  0.500 0.835 0.995 0.905 ;
        RECT  0.400 0.835 0.500 1.075 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.495 0.670 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 1.090 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.510 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.670 -0.115 2.240 0.115 ;
        RECT  0.590 -0.115 0.670 0.285 ;
        RECT  0.330 -0.115 0.590 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.145 2.240 1.375 ;
        RECT  2.100 0.975 2.200 1.375 ;
        RECT  1.840 1.145 2.100 1.375 ;
        RECT  1.740 0.975 1.840 1.375 ;
        RECT  1.260 1.145 1.740 1.375 ;
        RECT  1.160 0.975 1.260 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.800 0.975 0.900 1.375 ;
        RECT  0.680 1.145 0.800 1.375 ;
        RECT  0.580 0.975 0.680 1.375 ;
        RECT  0.320 1.145 0.580 1.375 ;
        RECT  0.220 0.975 0.320 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.205 2.030 0.275 ;
        RECT  1.920 0.530 2.020 0.765 ;
        RECT  0.330 0.695 1.920 0.765 ;
        RECT  1.250 0.345 1.630 0.415 ;
        RECT  1.170 0.205 1.250 0.415 ;
        RECT  0.790 0.205 1.170 0.275 ;
        RECT  0.500 0.355 1.090 0.425 ;
        RECT  0.400 0.185 0.500 0.425 ;
        RECT  0.260 0.345 0.330 0.905 ;
        RECT  0.130 0.345 0.260 0.415 ;
        RECT  0.130 0.835 0.260 0.905 ;
        RECT  0.050 0.265 0.130 0.415 ;
        RECT  0.050 0.835 0.130 1.005 ;
    END
END IND4D2BWP

MACRO IND4D4BWP
    CLASS CORE ;
    FOREIGN IND4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.345 3.560 0.455 ;
        RECT  3.535 0.750 3.545 1.050 ;
        RECT  3.475 0.345 3.535 1.050 ;
        RECT  3.325 0.345 3.475 0.915 ;
        RECT  3.090 0.345 3.325 0.455 ;
        RECT  3.185 0.750 3.325 0.915 ;
        RECT  3.115 0.750 3.185 1.050 ;
        RECT  0.570 0.845 3.115 0.915 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 1.090 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.925 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.765 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.200 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 3.780 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.860 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.860 0.275 ;
        RECT  0.490 -0.115 0.760 0.115 ;
        RECT  0.410 -0.115 0.490 0.445 ;
        RECT  0.150 -0.115 0.410 0.115 ;
        RECT  0.035 -0.115 0.150 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.675 3.730 1.375 ;
        RECT  3.380 1.145 3.650 1.375 ;
        RECT  3.280 0.990 3.380 1.375 ;
        RECT  3.020 1.145 3.280 1.375 ;
        RECT  2.920 0.990 3.020 1.375 ;
        RECT  2.480 1.145 2.920 1.375 ;
        RECT  2.380 0.990 2.480 1.375 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.020 0.990 2.120 1.375 ;
        RECT  1.760 1.145 2.020 1.375 ;
        RECT  1.660 0.990 1.760 1.375 ;
        RECT  1.220 1.145 1.660 1.375 ;
        RECT  1.120 0.990 1.220 1.375 ;
        RECT  0.860 1.145 1.120 1.375 ;
        RECT  0.760 0.990 0.860 1.375 ;
        RECT  0.490 1.145 0.760 1.375 ;
        RECT  0.410 0.845 0.490 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.090 0.345 3.255 0.455 ;
        RECT  3.185 0.750 3.255 0.915 ;
        RECT  3.115 0.750 3.185 1.050 ;
        RECT  0.570 0.845 3.115 0.915 ;
        RECT  3.650 0.205 3.730 0.465 ;
        RECT  3.010 0.205 3.650 0.275 ;
        RECT  3.000 0.545 3.245 0.615 ;
        RECT  2.930 0.205 3.010 0.465 ;
        RECT  2.930 0.545 3.000 0.775 ;
        RECT  2.190 0.205 2.930 0.275 ;
        RECT  0.340 0.705 2.930 0.775 ;
        RECT  2.110 0.345 2.850 0.415 ;
        RECT  2.030 0.195 2.110 0.415 ;
        RECT  1.290 0.195 2.030 0.265 ;
        RECT  1.025 0.355 1.950 0.425 ;
        RECT  0.955 0.190 1.025 0.425 ;
        RECT  0.680 0.355 0.955 0.425 ;
        RECT  0.580 0.185 0.680 0.425 ;
        RECT  0.310 0.190 0.340 0.775 ;
        RECT  0.270 0.190 0.310 1.015 ;
        RECT  0.235 0.190 0.270 0.450 ;
        RECT  0.230 0.705 0.270 1.015 ;
    END
END IND4D4BWP

MACRO INR2D0BWP
    CLASS CORE ;
    FOREIGN INR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0536 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.915 0.805 1.045 ;
        RECT  0.525 0.915 0.715 0.985 ;
        RECT  0.525 0.210 0.600 0.280 ;
        RECT  0.455 0.210 0.525 0.985 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.620 0.545 0.735 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.805 -0.115 0.840 0.115 ;
        RECT  0.690 -0.115 0.805 0.275 ;
        RECT  0.360 -0.115 0.690 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.840 1.375 ;
        RECT  0.240 0.985 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END INR2D0BWP

MACRO INR2D1BWP
    CLASS CORE ;
    FOREIGN INR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1071 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.825 0.805 1.065 ;
        RECT  0.525 0.825 0.700 0.905 ;
        RECT  0.525 0.195 0.590 0.435 ;
        RECT  0.455 0.195 0.525 0.905 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.620 0.540 0.735 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.805 -0.115 0.840 0.115 ;
        RECT  0.690 -0.115 0.805 0.275 ;
        RECT  0.360 -0.115 0.690 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.840 1.375 ;
        RECT  0.240 0.985 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.055 ;
    END
END INR2D1BWP

MACRO INR2D2BWP
    CLASS CORE ;
    FOREIGN INR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.910 0.275 ;
        RECT  0.525 0.715 0.710 0.785 ;
        RECT  0.440 0.205 0.525 0.785 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.685 0.520 0.735 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 -0.115 1.120 0.115 ;
        RECT  0.995 -0.115 1.065 0.450 ;
        RECT  0.720 -0.115 0.995 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.950 1.010 1.070 1.375 ;
        RECT  0.340 1.145 0.950 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.545 1.000 0.615 ;
        RECT  0.875 0.545 0.945 0.935 ;
        RECT  0.370 0.865 0.875 0.935 ;
        RECT  0.300 0.345 0.370 0.935 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.125 0.865 0.300 0.935 ;
        RECT  0.050 0.265 0.130 0.415 ;
        RECT  0.055 0.865 0.125 0.985 ;
    END
END INR2D2BWP

MACRO INR2D4BWP
    CLASS CORE ;
    FOREIGN INR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2884 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.210 1.890 0.420 ;
        RECT  1.670 0.210 1.740 0.795 ;
        RECT  1.515 0.210 1.670 0.420 ;
        RECT  1.570 0.710 1.670 0.795 ;
        RECT  0.860 0.210 1.515 0.285 ;
        RECT  0.860 0.710 0.910 0.790 ;
        RECT  0.790 0.210 0.860 0.790 ;
        RECT  0.690 0.210 0.790 0.285 ;
        RECT  0.610 0.210 0.690 0.470 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.520 1.600 0.640 ;
        RECT  1.365 0.355 1.435 0.640 ;
        RECT  1.085 0.355 1.365 0.425 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.930 0.520 1.015 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.465 ;
        RECT  1.700 -0.115 1.970 0.115 ;
        RECT  1.580 -0.115 1.700 0.140 ;
        RECT  1.300 -0.115 1.580 0.115 ;
        RECT  1.180 -0.115 1.300 0.140 ;
        RECT  0.900 -0.115 1.180 0.115 ;
        RECT  0.780 -0.115 0.900 0.140 ;
        RECT  0.510 -0.115 0.780 0.115 ;
        RECT  0.430 -0.115 0.510 0.460 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.145 2.100 1.375 ;
        RECT  1.950 0.700 2.030 1.375 ;
        RECT  1.300 1.145 1.950 1.375 ;
        RECT  1.180 1.005 1.300 1.375 ;
        RECT  0.510 1.145 1.180 1.375 ;
        RECT  0.430 0.700 0.510 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.420 1.740 0.795 ;
        RECT  1.570 0.710 1.670 0.795 ;
        RECT  0.860 0.210 1.515 0.285 ;
        RECT  0.860 0.710 0.910 0.790 ;
        RECT  0.790 0.210 0.860 0.790 ;
        RECT  0.690 0.210 0.790 0.285 ;
        RECT  0.610 0.210 0.690 0.470 ;
        RECT  1.880 0.545 2.000 0.615 ;
        RECT  1.810 0.545 1.880 0.935 ;
        RECT  1.275 0.865 1.810 0.935 ;
        RECT  1.205 0.520 1.275 0.935 ;
        RECT  0.715 0.865 1.205 0.935 ;
        RECT  0.645 0.545 0.715 0.935 ;
        RECT  0.330 0.545 0.645 0.615 ;
        RECT  0.260 0.200 0.330 1.025 ;
    END
END INR2D4BWP

MACRO INR2XD0BWP
    CLASS CORE ;
    FOREIGN INR2XD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0761 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.705 0.805 1.045 ;
        RECT  0.525 0.705 0.710 0.775 ;
        RECT  0.525 0.210 0.600 0.280 ;
        RECT  0.455 0.210 0.525 0.775 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.620 0.540 0.735 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.805 -0.115 0.840 0.115 ;
        RECT  0.695 -0.115 0.805 0.275 ;
        RECT  0.350 -0.115 0.695 0.115 ;
        RECT  0.250 -0.115 0.350 0.270 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.145 0.840 1.375 ;
        RECT  0.250 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.310 0.345 0.385 0.915 ;
        RECT  0.125 0.345 0.310 0.415 ;
        RECT  0.125 0.845 0.310 0.915 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.065 ;
    END
END INR2XD0BWP

MACRO INR2XD1BWP
    CLASS CORE ;
    FOREIGN INR2XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.910 0.275 ;
        RECT  0.525 0.715 0.710 0.785 ;
        RECT  0.455 0.205 0.525 0.785 ;
        RECT  0.410 0.205 0.455 0.275 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.685 0.520 0.735 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 -0.115 1.120 0.115 ;
        RECT  0.995 -0.115 1.065 0.300 ;
        RECT  0.720 -0.115 0.995 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.315 -0.115 0.600 0.115 ;
        RECT  0.245 -0.115 0.315 0.275 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.950 0.995 1.070 1.375 ;
        RECT  0.340 1.145 0.950 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.905 0.520 0.975 0.925 ;
        RECT  0.385 0.855 0.905 0.925 ;
        RECT  0.315 0.345 0.385 0.925 ;
        RECT  0.125 0.345 0.315 0.415 ;
        RECT  0.125 0.855 0.315 0.925 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  0.055 0.855 0.125 0.995 ;
    END
END INR2XD1BWP

MACRO INR2XD2BWP
    CLASS CORE ;
    FOREIGN INR2XD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2028 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.185 1.585 0.360 ;
        RECT  1.505 0.290 1.515 0.360 ;
        RECT  1.435 0.290 1.505 0.785 ;
        RECT  1.230 0.290 1.435 0.360 ;
        RECT  1.310 0.715 1.435 0.785 ;
        RECT  1.155 0.185 1.230 0.360 ;
        RECT  0.865 0.290 1.155 0.360 ;
        RECT  0.795 0.185 0.865 0.360 ;
        RECT  0.525 0.290 0.795 0.360 ;
        RECT  0.525 0.715 0.710 0.785 ;
        RECT  0.510 0.290 0.525 0.785 ;
        RECT  0.440 0.185 0.510 0.785 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.540 1.340 0.620 ;
        RECT  1.155 0.430 1.225 0.765 ;
        RECT  0.685 0.430 1.155 0.500 ;
        RECT  0.595 0.430 0.685 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.200 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.300 ;
        RECT  1.430 -0.115 1.690 0.115 ;
        RECT  1.310 -0.115 1.430 0.220 ;
        RECT  1.070 -0.115 1.310 0.115 ;
        RECT  0.950 -0.115 1.070 0.220 ;
        RECT  0.710 -0.115 0.950 0.115 ;
        RECT  0.590 -0.115 0.710 0.220 ;
        RECT  0.315 -0.115 0.590 0.115 ;
        RECT  0.245 -0.115 0.315 0.275 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.990 1.770 1.375 ;
        RECT  1.050 1.145 1.690 1.375 ;
        RECT  0.970 0.995 1.050 1.375 ;
        RECT  0.320 1.145 0.970 1.375 ;
        RECT  0.240 0.995 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.585 0.505 1.655 0.925 ;
        RECT  0.950 0.855 1.585 0.925 ;
        RECT  0.950 0.570 1.010 0.640 ;
        RECT  0.880 0.570 0.950 0.925 ;
        RECT  0.370 0.855 0.880 0.925 ;
        RECT  0.300 0.355 0.370 0.925 ;
        RECT  0.140 0.355 0.300 0.425 ;
        RECT  0.125 0.855 0.300 0.925 ;
        RECT  0.040 0.185 0.140 0.425 ;
        RECT  0.055 0.855 0.125 1.030 ;
    END
END INR2XD2BWP

MACRO INR2XD4BWP
    CLASS CORE ;
    FOREIGN INR2XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.775 2.870 0.880 ;
        RECT  2.400 0.185 2.500 0.425 ;
        RECT  2.135 0.350 2.400 0.425 ;
        RECT  1.945 0.350 2.135 0.880 ;
        RECT  1.925 0.185 1.945 0.880 ;
        RECT  1.855 0.185 1.925 0.425 ;
        RECT  1.680 0.775 1.925 0.880 ;
        RECT  1.405 0.350 1.855 0.425 ;
        RECT  1.335 0.195 1.405 0.425 ;
        RECT  1.045 0.350 1.335 0.425 ;
        RECT  0.975 0.195 1.045 0.425 ;
        RECT  0.685 0.350 0.975 0.425 ;
        RECT  0.615 0.195 0.685 0.425 ;
        RECT  0.325 0.350 0.615 0.425 ;
        RECT  0.255 0.195 0.325 0.425 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 1.440 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.605 0.765 ;
        RECT  3.450 0.495 3.535 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 -0.115 3.640 0.115 ;
        RECT  3.490 -0.115 3.570 0.425 ;
        RECT  3.210 -0.115 3.490 0.115 ;
        RECT  3.130 -0.115 3.210 0.465 ;
        RECT  2.670 -0.115 3.130 0.115 ;
        RECT  2.590 -0.115 2.670 0.465 ;
        RECT  2.320 -0.115 2.590 0.115 ;
        RECT  2.220 -0.115 2.320 0.270 ;
        RECT  2.140 -0.115 2.220 0.115 ;
        RECT  2.040 -0.115 2.140 0.270 ;
        RECT  1.780 -0.115 2.040 0.115 ;
        RECT  1.680 -0.115 1.780 0.270 ;
        RECT  1.600 -0.115 1.680 0.115 ;
        RECT  1.500 -0.115 1.600 0.270 ;
        RECT  1.230 -0.115 1.500 0.115 ;
        RECT  1.150 -0.115 1.230 0.270 ;
        RECT  0.870 -0.115 1.150 0.115 ;
        RECT  0.790 -0.115 0.870 0.270 ;
        RECT  0.510 -0.115 0.790 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.305 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.145 3.640 1.375 ;
        RECT  3.490 0.845 3.570 1.375 ;
        RECT  3.210 1.145 3.490 1.375 ;
        RECT  3.130 0.685 3.210 1.375 ;
        RECT  1.410 1.145 3.130 1.375 ;
        RECT  1.330 0.840 1.410 1.375 ;
        RECT  1.050 1.145 1.330 1.375 ;
        RECT  0.970 0.840 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.840 0.690 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.250 0.840 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.775 2.870 0.880 ;
        RECT  2.400 0.185 2.500 0.425 ;
        RECT  2.205 0.350 2.400 0.425 ;
        RECT  1.405 0.350 1.855 0.425 ;
        RECT  1.680 0.775 1.855 0.880 ;
        RECT  1.335 0.195 1.405 0.425 ;
        RECT  1.045 0.350 1.335 0.425 ;
        RECT  0.975 0.195 1.045 0.425 ;
        RECT  0.685 0.350 0.975 0.425 ;
        RECT  0.615 0.195 0.685 0.425 ;
        RECT  0.325 0.350 0.615 0.425 ;
        RECT  0.255 0.195 0.325 0.425 ;
        RECT  3.310 0.185 3.380 1.070 ;
        RECT  2.225 0.545 3.310 0.615 ;
        RECT  2.955 0.735 3.025 1.035 ;
        RECT  1.585 0.965 2.955 1.035 ;
        RECT  1.565 0.540 1.845 0.620 ;
        RECT  1.515 0.700 1.585 1.035 ;
        RECT  0.145 0.700 0.435 0.770 ;
        RECT  0.075 0.700 0.145 1.045 ;
        RECT  1.230 0.700 1.515 0.770 ;
        RECT  1.155 0.700 1.230 1.045 ;
        RECT  0.865 0.700 1.155 0.770 ;
        RECT  0.795 0.700 0.865 1.045 ;
        RECT  0.505 0.700 0.795 0.770 ;
        RECT  0.435 0.700 0.505 1.045 ;
    END
END INR2XD4BWP

MACRO INR3D0BWP
    CLASS CORE ;
    FOREIGN INR3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0869 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.205 0.945 1.045 ;
        RECT  0.855 0.205 0.875 0.345 ;
        RECT  0.850 0.885 0.875 1.045 ;
        RECT  0.440 0.205 0.855 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.810 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.640 ;
        RECT  0.545 0.520 0.595 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.135 ;
        RECT  0.360 -0.115 0.640 0.115 ;
        RECT  0.240 -0.115 0.360 0.280 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.980 1.375 ;
        RECT  0.260 0.975 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.320 0.350 0.390 0.905 ;
        RECT  0.145 0.350 0.320 0.420 ;
        RECT  0.160 0.835 0.320 0.905 ;
        RECT  0.060 0.835 0.160 1.075 ;
        RECT  0.075 0.185 0.145 0.420 ;
    END
END INR3D0BWP

MACRO INR3D1BWP
    CLASS CORE ;
    FOREIGN INR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1369 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.360 1.505 0.920 ;
        RECT  1.330 0.360 1.435 0.430 ;
        RECT  1.280 0.840 1.435 0.920 ;
        RECT  1.260 0.205 1.330 0.430 ;
        RECT  1.210 0.840 1.280 1.045 ;
        RECT  0.420 0.205 1.260 0.275 ;
        RECT  0.780 0.975 1.210 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.540 1.200 0.625 ;
        RECT  1.015 0.345 1.085 0.625 ;
        RECT  0.665 0.345 1.015 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        RECT  0.520 0.540 0.595 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.290 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.000 -0.115 1.120 0.135 ;
        RECT  0.740 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.320 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.320 0.285 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.145 1.540 1.375 ;
        RECT  1.360 0.990 1.460 1.375 ;
        RECT  0.340 1.145 1.360 1.375 ;
        RECT  0.220 0.975 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.290 0.510 1.365 0.770 ;
        RECT  1.140 0.700 1.290 0.770 ;
        RECT  1.070 0.700 1.140 0.905 ;
        RECT  0.400 0.835 1.070 0.905 ;
        RECT  0.325 0.355 0.400 0.905 ;
        RECT  0.140 0.355 0.325 0.425 ;
        RECT  0.140 0.835 0.325 0.905 ;
        RECT  0.040 0.185 0.140 0.425 ;
        RECT  0.040 0.835 0.140 1.075 ;
    END
END INR3D1BWP

MACRO INR3D2BWP
    CLASS CORE ;
    FOREIGN INR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2082 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.360 1.505 0.920 ;
        RECT  1.330 0.360 1.435 0.430 ;
        RECT  1.290 0.850 1.435 0.920 ;
        RECT  1.260 0.205 1.330 0.430 ;
        RECT  1.220 0.850 1.290 1.045 ;
        RECT  0.420 0.205 1.260 0.275 ;
        RECT  0.780 0.975 1.220 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.540 1.200 0.625 ;
        RECT  1.015 0.345 1.085 0.625 ;
        RECT  0.665 0.345 1.015 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        RECT  0.520 0.540 0.595 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.290 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.000 -0.115 1.120 0.135 ;
        RECT  0.740 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.320 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.320 0.285 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.145 1.540 1.375 ;
        RECT  1.360 0.990 1.460 1.375 ;
        RECT  0.340 1.145 1.360 1.375 ;
        RECT  0.220 0.975 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.290 0.510 1.365 0.780 ;
        RECT  1.150 0.710 1.290 0.780 ;
        RECT  1.080 0.710 1.150 0.905 ;
        RECT  0.400 0.835 1.080 0.905 ;
        RECT  0.325 0.355 0.400 0.905 ;
        RECT  0.140 0.355 0.325 0.425 ;
        RECT  0.140 0.835 0.325 0.905 ;
        RECT  0.040 0.185 0.140 0.425 ;
        RECT  0.040 0.835 0.140 1.075 ;
    END
END INR3D2BWP

MACRO INR3D4BWP
    CLASS CORE ;
    FOREIGN INR3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3752 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.710 2.710 0.915 ;
        RECT  2.615 0.190 2.685 0.450 ;
        RECT  2.415 0.355 2.615 0.450 ;
        RECT  2.345 0.355 2.415 0.915 ;
        RECT  2.260 0.190 2.345 0.915 ;
        RECT  2.205 0.355 2.260 0.915 ;
        RECT  1.965 0.355 2.205 0.425 ;
        RECT  1.895 0.190 1.965 0.425 ;
        RECT  1.605 0.355 1.895 0.425 ;
        RECT  1.535 0.190 1.605 0.425 ;
        RECT  1.065 0.355 1.535 0.425 ;
        RECT  0.995 0.190 1.065 0.425 ;
        RECT  0.720 0.355 0.995 0.425 ;
        RECT  0.620 0.185 0.720 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.625 ;
        RECT  2.710 0.540 2.835 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 0.495 1.970 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.870 -0.115 2.940 0.115 ;
        RECT  2.790 -0.115 2.870 0.275 ;
        RECT  2.510 -0.115 2.790 0.115 ;
        RECT  2.430 -0.115 2.510 0.285 ;
        RECT  2.150 -0.115 2.430 0.115 ;
        RECT  2.070 -0.115 2.150 0.285 ;
        RECT  1.790 -0.115 2.070 0.115 ;
        RECT  1.710 -0.115 1.790 0.285 ;
        RECT  1.430 -0.115 1.710 0.115 ;
        RECT  1.350 -0.115 1.430 0.285 ;
        RECT  1.250 -0.115 1.350 0.115 ;
        RECT  1.170 -0.115 1.250 0.285 ;
        RECT  0.890 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.890 0.285 ;
        RECT  0.520 -0.115 0.810 0.115 ;
        RECT  0.440 -0.115 0.520 0.450 ;
        RECT  0.150 -0.115 0.440 0.115 ;
        RECT  0.070 -0.115 0.150 0.425 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.145 2.940 1.375 ;
        RECT  1.170 0.835 1.250 1.375 ;
        RECT  0.890 1.145 1.170 1.375 ;
        RECT  0.810 0.835 0.890 1.375 ;
        RECT  0.520 1.145 0.810 1.375 ;
        RECT  0.440 0.740 0.520 1.375 ;
        RECT  0.150 1.145 0.440 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.710 2.710 0.915 ;
        RECT  2.615 0.190 2.685 0.450 ;
        RECT  2.485 0.355 2.615 0.450 ;
        RECT  1.965 0.355 2.135 0.425 ;
        RECT  1.895 0.190 1.965 0.425 ;
        RECT  1.605 0.355 1.895 0.425 ;
        RECT  1.535 0.190 1.605 0.425 ;
        RECT  1.065 0.355 1.535 0.425 ;
        RECT  0.995 0.190 1.065 0.425 ;
        RECT  0.720 0.355 0.995 0.425 ;
        RECT  0.620 0.185 0.720 0.425 ;
        RECT  2.790 0.765 2.870 1.065 ;
        RECT  1.785 0.995 2.790 1.065 ;
        RECT  1.890 0.695 1.970 0.905 ;
        RECT  1.610 0.695 1.890 0.765 ;
        RECT  1.715 0.835 1.785 1.065 ;
        RECT  1.450 0.995 1.715 1.065 ;
        RECT  1.530 0.695 1.610 0.905 ;
        RECT  1.065 0.695 1.530 0.765 ;
        RECT  1.330 0.835 1.450 1.065 ;
        RECT  0.330 0.545 1.070 0.615 ;
        RECT  0.995 0.695 1.065 1.025 ;
        RECT  0.705 0.695 0.995 0.765 ;
        RECT  0.635 0.695 0.705 1.025 ;
        RECT  0.260 0.190 0.330 1.075 ;
    END
END INR3D4BWP

MACRO INR4D0BWP
    CLASS CORE ;
    FOREIGN INR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1029 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 1.075 ;
        RECT  0.985 0.355 1.155 0.425 ;
        RECT  1.090 0.835 1.155 1.075 ;
        RECT  0.915 0.190 0.985 0.425 ;
        RECT  0.585 0.355 0.915 0.425 ;
        RECT  0.515 0.190 0.585 0.425 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.840 0.640 ;
        RECT  0.735 0.495 0.805 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.495 0.665 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0186 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.200 -0.115 1.260 0.115 ;
        RECT  1.080 -0.115 1.200 0.285 ;
        RECT  0.810 -0.115 1.080 0.115 ;
        RECT  0.690 -0.115 0.810 0.285 ;
        RECT  0.390 -0.115 0.690 0.115 ;
        RECT  0.270 -0.115 0.390 0.135 ;
        RECT  0.000 -0.115 0.270 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.145 1.260 1.375 ;
        RECT  0.290 0.835 0.370 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.205 0.435 0.765 ;
        RECT  0.060 0.205 0.365 0.275 ;
        RECT  0.155 0.695 0.365 0.765 ;
        RECT  0.085 0.695 0.155 1.075 ;
    END
END INR4D0BWP

MACRO INR4D1BWP
    CLASS CORE ;
    FOREIGN INR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1338 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.355 1.870 0.425 ;
        RECT  1.365 0.845 1.690 0.915 ;
        RECT  1.295 0.355 1.365 0.915 ;
        RECT  0.590 0.355 1.295 0.425 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.665 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.065 0.625 ;
        RECT  1.870 0.540 1.995 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.575 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.040 -0.115 2.100 0.115 ;
        RECT  1.940 -0.115 2.040 0.275 ;
        RECT  1.640 -0.115 1.940 0.115 ;
        RECT  1.520 -0.115 1.640 0.275 ;
        RECT  0.940 -0.115 1.520 0.115 ;
        RECT  0.820 -0.115 0.940 0.275 ;
        RECT  0.510 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.510 0.425 ;
        RECT  0.160 -0.115 0.430 0.115 ;
        RECT  0.060 -0.115 0.160 0.275 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.145 2.100 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.150 1.145 0.780 1.375 ;
        RECT  0.070 0.935 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.955 0.745 2.025 1.055 ;
        RECT  0.410 0.985 1.955 1.055 ;
        RECT  0.800 0.520 0.880 0.915 ;
        RECT  0.330 0.845 0.800 0.915 ;
        RECT  0.260 0.185 0.330 1.055 ;
    END
END INR4D1BWP

MACRO INR4D2BWP
    CLASS CORE ;
    FOREIGN INR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.845 2.730 0.915 ;
        RECT  2.345 0.215 2.490 0.345 ;
        RECT  2.275 0.215 2.345 0.915 ;
        RECT  0.590 0.215 2.275 0.345 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.625 ;
        RECT  2.415 0.445 2.695 0.515 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.445 2.005 0.515 ;
        RECT  1.715 0.445 1.925 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.445 1.440 0.515 ;
        RECT  1.155 0.445 1.365 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.490 -0.115 2.940 0.115 ;
        RECT  0.410 -0.115 0.490 0.320 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.145 2.940 1.375 ;
        RECT  0.770 0.765 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.950 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.950 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.810 0.910 2.890 1.065 ;
        RECT  2.170 0.995 2.810 1.065 ;
        RECT  2.090 0.625 2.170 1.065 ;
        RECT  1.830 0.995 2.090 1.065 ;
        RECT  1.600 0.695 2.010 0.765 ;
        RECT  1.710 0.855 1.830 1.065 ;
        RECT  1.520 0.625 1.600 1.065 ;
        RECT  1.230 0.855 1.520 0.925 ;
        RECT  1.030 0.695 1.410 0.765 ;
        RECT  1.110 0.855 1.230 1.065 ;
        RECT  0.950 0.625 1.030 1.065 ;
        RECT  0.670 0.625 0.950 0.695 ;
        RECT  0.340 0.445 0.870 0.515 ;
        RECT  0.590 0.625 0.670 1.065 ;
        RECT  0.270 0.215 0.340 1.045 ;
        RECT  0.210 0.215 0.270 0.285 ;
        RECT  0.210 0.975 0.270 1.045 ;
    END
END INR4D2BWP

MACRO INR4D4BWP
    CLASS CORE ;
    FOREIGN INR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4620 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.775 3.570 0.905 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.395 0.345 3.475 0.465 ;
        RECT  3.190 0.345 3.395 0.905 ;
        RECT  3.185 0.185 3.190 0.905 ;
        RECT  3.110 0.185 3.185 0.415 ;
        RECT  3.090 0.775 3.185 0.905 ;
        RECT  2.650 0.345 3.110 0.415 ;
        RECT  2.570 0.185 2.650 0.415 ;
        RECT  2.290 0.345 2.570 0.415 ;
        RECT  2.210 0.185 2.290 0.415 ;
        RECT  1.930 0.345 2.210 0.415 ;
        RECT  1.850 0.185 1.930 0.415 ;
        RECT  1.570 0.345 1.850 0.415 ;
        RECT  1.490 0.185 1.570 0.415 ;
        RECT  1.030 0.345 1.490 0.415 ;
        RECT  0.950 0.185 1.030 0.415 ;
        RECT  0.690 0.345 0.950 0.415 ;
        RECT  0.570 0.210 0.690 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.550 0.540 3.675 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.495 2.700 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.930 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.740 -0.115 3.780 0.115 ;
        RECT  3.640 -0.115 3.740 0.275 ;
        RECT  3.380 -0.115 3.640 0.115 ;
        RECT  3.280 -0.115 3.380 0.275 ;
        RECT  3.020 -0.115 3.280 0.115 ;
        RECT  2.920 -0.115 3.020 0.275 ;
        RECT  2.840 -0.115 2.920 0.115 ;
        RECT  2.740 -0.115 2.840 0.275 ;
        RECT  2.480 -0.115 2.740 0.115 ;
        RECT  2.380 -0.115 2.480 0.275 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.020 -0.115 2.120 0.275 ;
        RECT  1.760 -0.115 2.020 0.115 ;
        RECT  1.660 -0.115 1.760 0.275 ;
        RECT  1.400 -0.115 1.660 0.115 ;
        RECT  1.300 -0.115 1.400 0.275 ;
        RECT  1.220 -0.115 1.300 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.860 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.860 0.275 ;
        RECT  0.490 -0.115 0.760 0.115 ;
        RECT  0.410 -0.115 0.490 0.465 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 3.780 1.375 ;
        RECT  1.120 0.850 1.220 1.375 ;
        RECT  0.860 1.145 1.120 1.375 ;
        RECT  0.760 0.850 0.860 1.375 ;
        RECT  0.490 1.145 0.760 1.375 ;
        RECT  0.410 0.685 0.490 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.775 3.570 0.905 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.465 0.345 3.475 0.465 ;
        RECT  3.110 0.185 3.115 0.415 ;
        RECT  3.090 0.775 3.115 0.905 ;
        RECT  2.650 0.345 3.110 0.415 ;
        RECT  2.570 0.185 2.650 0.415 ;
        RECT  2.290 0.345 2.570 0.415 ;
        RECT  2.210 0.185 2.290 0.415 ;
        RECT  1.930 0.345 2.210 0.415 ;
        RECT  1.850 0.185 1.930 0.415 ;
        RECT  1.570 0.345 1.850 0.415 ;
        RECT  1.490 0.185 1.570 0.415 ;
        RECT  1.030 0.345 1.490 0.415 ;
        RECT  0.950 0.185 1.030 0.415 ;
        RECT  0.690 0.345 0.950 0.415 ;
        RECT  0.570 0.210 0.690 0.415 ;
        RECT  3.650 0.755 3.730 1.055 ;
        RECT  3.010 0.985 3.650 1.055 ;
        RECT  2.930 0.715 3.010 1.055 ;
        RECT  2.190 0.715 2.930 0.785 ;
        RECT  2.110 0.865 2.850 0.935 ;
        RECT  2.030 0.675 2.110 1.075 ;
        RECT  1.290 0.865 2.030 0.935 ;
        RECT  1.025 0.710 1.950 0.780 ;
        RECT  0.330 0.545 1.035 0.615 ;
        RECT  0.955 0.710 1.025 1.040 ;
        RECT  0.665 0.710 0.955 0.780 ;
        RECT  0.595 0.710 0.665 1.040 ;
        RECT  0.260 0.185 0.330 1.045 ;
        RECT  0.220 0.185 0.260 0.425 ;
        RECT  0.230 0.765 0.260 1.045 ;
    END
END INR4D4BWP

MACRO INVD0BWP
    CLASS CORE ;
    FOREIGN INVD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.215 0.385 1.045 ;
        RECT  0.240 0.215 0.315 0.295 ;
        RECT  0.240 0.965 0.315 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.160 -0.115 0.420 0.115 ;
        RECT  0.080 -0.115 0.160 0.325 ;
        RECT  0.000 -0.115 0.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.145 0.420 1.375 ;
        RECT  0.080 0.935 0.160 1.375 ;
        RECT  0.000 1.145 0.080 1.375 ;
        END
    END VDD
END INVD0BWP

MACRO INVD12BWP
    CLASS CORE ;
    FOREIGN INVD12BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6048 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.695 2.125 1.035 ;
        RECT  1.765 0.300 2.055 0.465 ;
        RECT  1.765 0.695 2.055 0.885 ;
        RECT  1.695 0.185 1.765 0.465 ;
        RECT  1.695 0.695 1.765 1.035 ;
        RECT  1.435 0.300 1.695 0.465 ;
        RECT  1.435 0.695 1.695 0.885 ;
        RECT  1.405 0.300 1.435 0.885 ;
        RECT  1.335 0.185 1.405 1.035 ;
        RECT  1.085 0.300 1.335 0.885 ;
        RECT  1.045 0.300 1.085 0.465 ;
        RECT  1.045 0.695 1.085 0.885 ;
        RECT  0.975 0.185 1.045 0.465 ;
        RECT  0.975 0.695 1.045 1.035 ;
        RECT  0.685 0.300 0.975 0.465 ;
        RECT  0.685 0.695 0.975 0.885 ;
        RECT  0.615 0.185 0.685 0.465 ;
        RECT  0.615 0.695 0.685 1.035 ;
        RECT  0.325 0.300 0.615 0.465 ;
        RECT  0.325 0.695 0.615 0.885 ;
        RECT  0.255 0.185 0.325 0.465 ;
        RECT  0.255 0.695 0.325 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.995 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.115 2.380 0.115 ;
        RECT  2.235 -0.115 2.305 0.465 ;
        RECT  1.970 -0.115 2.235 0.115 ;
        RECT  1.850 -0.115 1.970 0.230 ;
        RECT  1.610 -0.115 1.850 0.115 ;
        RECT  1.490 -0.115 1.610 0.230 ;
        RECT  1.250 -0.115 1.490 0.115 ;
        RECT  1.130 -0.115 1.250 0.230 ;
        RECT  0.890 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.890 0.230 ;
        RECT  0.530 -0.115 0.770 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.150 -0.115 0.410 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.145 2.380 1.375 ;
        RECT  2.230 0.685 2.310 1.375 ;
        RECT  1.970 1.145 2.230 1.375 ;
        RECT  1.850 0.955 1.970 1.375 ;
        RECT  1.610 1.145 1.850 1.375 ;
        RECT  1.490 0.955 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 0.955 1.250 1.375 ;
        RECT  0.890 1.145 1.130 1.375 ;
        RECT  0.770 0.955 0.890 1.375 ;
        RECT  0.530 1.145 0.770 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.150 1.145 0.410 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.695 2.125 1.035 ;
        RECT  1.765 0.300 2.055 0.465 ;
        RECT  1.765 0.695 2.055 0.885 ;
        RECT  1.695 0.185 1.765 0.465 ;
        RECT  1.695 0.695 1.765 1.035 ;
        RECT  1.505 0.300 1.695 0.465 ;
        RECT  1.505 0.695 1.695 0.885 ;
        RECT  0.975 0.185 1.015 0.465 ;
        RECT  0.975 0.695 1.015 1.035 ;
        RECT  0.685 0.300 0.975 0.465 ;
        RECT  0.685 0.695 0.975 0.885 ;
        RECT  0.615 0.185 0.685 0.465 ;
        RECT  0.615 0.695 0.685 1.035 ;
        RECT  0.325 0.300 0.615 0.465 ;
        RECT  0.325 0.695 0.615 0.885 ;
        RECT  0.255 0.185 0.325 0.465 ;
        RECT  0.255 0.695 0.325 1.035 ;
        RECT  1.515 0.545 2.185 0.615 ;
    END
END INVD12BWP

MACRO INVD16BWP
    CLASS CORE ;
    FOREIGN INVD16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8064 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.775 0.695 2.845 1.035 ;
        RECT  2.485 0.300 2.775 0.465 ;
        RECT  2.485 0.695 2.775 0.885 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.695 2.485 1.035 ;
        RECT  2.125 0.300 2.415 0.465 ;
        RECT  2.125 0.695 2.415 0.885 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.695 2.125 1.035 ;
        RECT  1.765 0.300 2.055 0.465 ;
        RECT  1.770 0.695 2.055 0.885 ;
        RECT  1.715 0.695 1.770 1.045 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.695 0.185 1.715 1.045 ;
        RECT  1.385 0.300 1.695 0.885 ;
        RECT  1.365 0.185 1.385 1.045 ;
        RECT  1.315 0.185 1.365 0.465 ;
        RECT  1.315 0.695 1.365 1.045 ;
        RECT  1.025 0.300 1.315 0.465 ;
        RECT  1.025 0.695 1.315 0.885 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.035 ;
        RECT  0.665 0.300 0.955 0.465 ;
        RECT  0.665 0.695 0.955 0.885 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4608 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.255 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.465 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.230 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.230 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.230 ;
        RECT  1.600 -0.115 1.850 0.115 ;
        RECT  1.480 -0.115 1.600 0.230 ;
        RECT  1.230 -0.115 1.480 0.115 ;
        RECT  1.110 -0.115 1.230 0.230 ;
        RECT  0.870 -0.115 1.110 0.115 ;
        RECT  0.750 -0.115 0.870 0.230 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.230 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.680 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 0.955 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 0.955 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 0.955 1.970 1.375 ;
        RECT  1.600 1.145 1.850 1.375 ;
        RECT  1.480 0.955 1.600 1.375 ;
        RECT  1.230 1.145 1.480 1.375 ;
        RECT  1.110 0.955 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 0.955 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.955 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.775 0.695 2.845 1.035 ;
        RECT  2.485 0.300 2.775 0.465 ;
        RECT  2.485 0.695 2.775 0.885 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.695 2.485 1.035 ;
        RECT  2.125 0.300 2.415 0.465 ;
        RECT  2.125 0.695 2.415 0.885 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.695 2.125 1.035 ;
        RECT  1.785 0.300 2.055 0.465 ;
        RECT  1.785 0.695 2.055 0.885 ;
        RECT  1.025 0.300 1.295 0.465 ;
        RECT  1.025 0.695 1.295 0.885 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.035 ;
        RECT  0.665 0.300 0.955 0.465 ;
        RECT  0.665 0.695 0.955 0.885 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        RECT  1.840 0.545 2.880 0.615 ;
    END
END INVD16BWP

MACRO INVD1BWP
    CLASS CORE ;
    FOREIGN INVD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.185 0.385 1.045 ;
        RECT  0.280 0.185 0.315 0.430 ;
        RECT  0.295 0.735 0.315 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.115 0.420 0.115 ;
        RECT  0.115 -0.115 0.185 0.415 ;
        RECT  0.000 -0.115 0.115 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.145 0.420 1.375 ;
        RECT  0.115 0.845 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
END INVD1BWP

MACRO INVD20BWP
    CLASS CORE ;
    FOREIGN INVD20BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.0080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.475 0.695 3.545 1.035 ;
        RECT  3.185 0.300 3.475 0.465 ;
        RECT  3.185 0.695 3.475 0.885 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.695 3.185 1.035 ;
        RECT  2.825 0.300 3.115 0.465 ;
        RECT  2.825 0.695 3.115 0.885 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.755 0.695 2.825 1.035 ;
        RECT  2.465 0.300 2.755 0.465 ;
        RECT  2.465 0.695 2.755 0.885 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.395 0.695 2.465 1.035 ;
        RECT  2.135 0.300 2.395 0.465 ;
        RECT  2.135 0.695 2.395 0.885 ;
        RECT  2.105 0.300 2.135 0.885 ;
        RECT  2.035 0.185 2.105 1.035 ;
        RECT  1.785 0.300 2.035 0.885 ;
        RECT  1.745 0.300 1.785 0.465 ;
        RECT  1.745 0.695 1.785 0.885 ;
        RECT  1.675 0.185 1.745 0.465 ;
        RECT  1.675 0.695 1.745 1.035 ;
        RECT  1.385 0.300 1.675 0.465 ;
        RECT  1.385 0.695 1.675 0.885 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.315 0.695 1.385 1.035 ;
        RECT  1.025 0.300 1.315 0.465 ;
        RECT  1.025 0.695 1.315 0.885 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.035 ;
        RECT  0.665 0.300 0.955 0.465 ;
        RECT  0.665 0.695 0.955 0.885 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.5760 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.675 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.465 ;
        RECT  3.390 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.390 0.230 ;
        RECT  3.030 -0.115 3.270 0.115 ;
        RECT  2.910 -0.115 3.030 0.230 ;
        RECT  2.670 -0.115 2.910 0.115 ;
        RECT  2.550 -0.115 2.670 0.230 ;
        RECT  2.310 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.310 0.230 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.230 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.230 ;
        RECT  1.230 -0.115 1.470 0.115 ;
        RECT  1.110 -0.115 1.230 0.230 ;
        RECT  0.870 -0.115 1.110 0.115 ;
        RECT  0.750 -0.115 0.870 0.230 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.230 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.685 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 0.955 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 0.955 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 0.955 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 0.955 2.310 1.375 ;
        RECT  1.950 1.145 2.190 1.375 ;
        RECT  1.830 0.955 1.950 1.375 ;
        RECT  1.590 1.145 1.830 1.375 ;
        RECT  1.470 0.955 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 0.955 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 0.955 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.955 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.475 0.695 3.545 1.035 ;
        RECT  3.185 0.300 3.475 0.465 ;
        RECT  3.185 0.695 3.475 0.885 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.695 3.185 1.035 ;
        RECT  2.825 0.300 3.115 0.465 ;
        RECT  2.825 0.695 3.115 0.885 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.755 0.695 2.825 1.035 ;
        RECT  2.465 0.300 2.755 0.465 ;
        RECT  2.465 0.695 2.755 0.885 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.395 0.695 2.465 1.035 ;
        RECT  2.205 0.300 2.395 0.465 ;
        RECT  2.205 0.695 2.395 0.885 ;
        RECT  1.675 0.185 1.715 0.465 ;
        RECT  1.675 0.695 1.715 1.035 ;
        RECT  1.385 0.300 1.675 0.465 ;
        RECT  1.385 0.695 1.675 0.885 ;
        RECT  1.315 0.185 1.385 0.465 ;
        RECT  1.315 0.695 1.385 1.035 ;
        RECT  1.025 0.300 1.315 0.465 ;
        RECT  1.025 0.695 1.315 0.885 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.035 ;
        RECT  0.665 0.300 0.955 0.465 ;
        RECT  0.665 0.695 0.955 0.885 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        RECT  2.245 0.545 3.645 0.615 ;
    END
END INVD20BWP

MACRO INVD24BWP
    CLASS CORE ;
    FOREIGN INVD24BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.2096 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.255 0.185 4.325 0.465 ;
        RECT  4.255 0.695 4.325 1.035 ;
        RECT  3.965 0.300 4.255 0.465 ;
        RECT  3.965 0.695 4.255 0.885 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.695 3.965 1.035 ;
        RECT  3.605 0.300 3.895 0.465 ;
        RECT  3.605 0.695 3.895 0.885 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.695 3.605 1.035 ;
        RECT  3.245 0.300 3.535 0.465 ;
        RECT  3.245 0.695 3.535 0.885 ;
        RECT  3.175 0.185 3.245 0.465 ;
        RECT  3.175 0.695 3.245 1.035 ;
        RECT  2.885 0.300 3.175 0.465 ;
        RECT  2.885 0.695 3.175 0.885 ;
        RECT  2.815 0.185 2.885 0.465 ;
        RECT  2.815 0.695 2.885 1.035 ;
        RECT  2.525 0.300 2.815 0.465 ;
        RECT  2.525 0.695 2.815 0.885 ;
        RECT  2.455 0.185 2.525 0.465 ;
        RECT  2.455 0.695 2.525 1.035 ;
        RECT  2.415 0.300 2.455 0.465 ;
        RECT  2.415 0.695 2.455 0.885 ;
        RECT  2.165 0.300 2.415 0.885 ;
        RECT  2.095 0.185 2.165 1.035 ;
        RECT  2.065 0.300 2.095 0.885 ;
        RECT  1.805 0.300 2.065 0.465 ;
        RECT  1.805 0.695 2.065 0.885 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.735 0.695 1.805 1.035 ;
        RECT  1.445 0.300 1.735 0.465 ;
        RECT  1.445 0.695 1.735 0.885 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.695 1.445 1.035 ;
        RECT  1.085 0.300 1.375 0.465 ;
        RECT  1.085 0.695 1.375 0.885 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.695 1.085 1.035 ;
        RECT  0.725 0.300 1.015 0.465 ;
        RECT  0.725 0.695 1.015 0.885 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.695 0.725 1.035 ;
        RECT  0.365 0.300 0.655 0.465 ;
        RECT  0.365 0.695 0.655 0.885 ;
        RECT  0.295 0.185 0.365 0.465 ;
        RECT  0.295 0.695 0.365 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6912 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.965 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.115 4.620 0.115 ;
        RECT  4.420 -0.115 4.520 0.455 ;
        RECT  4.170 -0.115 4.420 0.115 ;
        RECT  4.050 -0.115 4.170 0.230 ;
        RECT  3.810 -0.115 4.050 0.115 ;
        RECT  3.690 -0.115 3.810 0.230 ;
        RECT  3.450 -0.115 3.690 0.115 ;
        RECT  3.330 -0.115 3.450 0.230 ;
        RECT  3.090 -0.115 3.330 0.115 ;
        RECT  2.970 -0.115 3.090 0.230 ;
        RECT  2.730 -0.115 2.970 0.115 ;
        RECT  2.610 -0.115 2.730 0.230 ;
        RECT  2.370 -0.115 2.610 0.115 ;
        RECT  2.250 -0.115 2.370 0.230 ;
        RECT  2.010 -0.115 2.250 0.115 ;
        RECT  1.890 -0.115 2.010 0.230 ;
        RECT  1.650 -0.115 1.890 0.115 ;
        RECT  1.530 -0.115 1.650 0.230 ;
        RECT  1.290 -0.115 1.530 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.930 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.570 -0.115 0.810 0.115 ;
        RECT  0.450 -0.115 0.570 0.230 ;
        RECT  0.200 -0.115 0.450 0.115 ;
        RECT  0.100 -0.115 0.200 0.415 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.145 4.620 1.375 ;
        RECT  4.420 0.695 4.520 1.375 ;
        RECT  4.170 1.145 4.420 1.375 ;
        RECT  4.050 0.955 4.170 1.375 ;
        RECT  3.810 1.145 4.050 1.375 ;
        RECT  3.690 0.955 3.810 1.375 ;
        RECT  3.450 1.145 3.690 1.375 ;
        RECT  3.330 0.955 3.450 1.375 ;
        RECT  3.090 1.145 3.330 1.375 ;
        RECT  2.970 0.955 3.090 1.375 ;
        RECT  2.730 1.145 2.970 1.375 ;
        RECT  2.610 0.955 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 0.955 2.370 1.375 ;
        RECT  2.010 1.145 2.250 1.375 ;
        RECT  1.890 0.955 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 0.955 1.650 1.375 ;
        RECT  1.290 1.145 1.530 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.930 1.145 1.170 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.570 1.145 0.810 1.375 ;
        RECT  0.450 0.955 0.570 1.375 ;
        RECT  0.200 1.145 0.450 1.375 ;
        RECT  0.100 0.845 0.200 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.255 0.185 4.325 0.465 ;
        RECT  4.255 0.695 4.325 1.035 ;
        RECT  3.965 0.300 4.255 0.465 ;
        RECT  3.965 0.695 4.255 0.885 ;
        RECT  3.895 0.185 3.965 0.465 ;
        RECT  3.895 0.695 3.965 1.035 ;
        RECT  3.605 0.300 3.895 0.465 ;
        RECT  3.605 0.695 3.895 0.885 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.695 3.605 1.035 ;
        RECT  3.245 0.300 3.535 0.465 ;
        RECT  3.245 0.695 3.535 0.885 ;
        RECT  3.175 0.185 3.245 0.465 ;
        RECT  3.175 0.695 3.245 1.035 ;
        RECT  2.885 0.300 3.175 0.465 ;
        RECT  2.885 0.695 3.175 0.885 ;
        RECT  2.815 0.185 2.885 0.465 ;
        RECT  2.815 0.695 2.885 1.035 ;
        RECT  2.525 0.300 2.815 0.465 ;
        RECT  2.525 0.695 2.815 0.885 ;
        RECT  2.485 0.185 2.525 0.465 ;
        RECT  2.485 0.695 2.525 1.035 ;
        RECT  1.805 0.300 1.995 0.465 ;
        RECT  1.805 0.695 1.995 0.885 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.735 0.695 1.805 1.035 ;
        RECT  1.445 0.300 1.735 0.465 ;
        RECT  1.445 0.695 1.735 0.885 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.695 1.445 1.035 ;
        RECT  1.085 0.300 1.375 0.465 ;
        RECT  1.085 0.695 1.375 0.885 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.695 1.085 1.035 ;
        RECT  0.725 0.300 1.015 0.465 ;
        RECT  0.725 0.695 1.015 0.885 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.695 0.725 1.035 ;
        RECT  0.365 0.300 0.655 0.465 ;
        RECT  0.365 0.695 0.655 0.885 ;
        RECT  0.295 0.185 0.365 0.465 ;
        RECT  0.295 0.695 0.365 1.035 ;
        RECT  2.515 0.545 4.435 0.615 ;
    END
END INVD24BWP

MACRO INVD2BWP
    CLASS CORE ;
    FOREIGN INVD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.355 0.385 0.815 ;
        RECT  0.315 0.185 0.320 0.815 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.735 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.515 -0.115 0.560 0.115 ;
        RECT  0.405 -0.115 0.515 0.280 ;
        RECT  0.150 -0.115 0.405 0.115 ;
        RECT  0.050 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.145 0.560 1.375 ;
        RECT  0.420 0.910 0.500 1.375 ;
        RECT  0.150 1.145 0.420 1.375 ;
        RECT  0.050 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END INVD2BWP

MACRO INVD3BWP
    CLASS CORE ;
    FOREIGN INVD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1944 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 0.195 0.760 0.455 ;
        RECT  0.685 0.705 0.755 1.035 ;
        RECT  0.595 0.705 0.685 0.820 ;
        RECT  0.595 0.340 0.680 0.455 ;
        RECT  0.385 0.340 0.595 0.820 ;
        RECT  0.340 0.340 0.385 0.455 ;
        RECT  0.335 0.705 0.385 0.820 ;
        RECT  0.260 0.195 0.340 0.455 ;
        RECT  0.265 0.705 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 -0.115 0.840 0.115 ;
        RECT  0.450 -0.115 0.570 0.260 ;
        RECT  0.160 -0.115 0.450 0.115 ;
        RECT  0.080 -0.115 0.160 0.415 ;
        RECT  0.000 -0.115 0.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.145 0.840 1.375 ;
        RECT  0.450 0.890 0.570 1.375 ;
        RECT  0.160 1.145 0.450 1.375 ;
        RECT  0.080 0.845 0.160 1.375 ;
        RECT  0.000 1.145 0.080 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.680 0.195 0.760 0.455 ;
        RECT  0.685 0.705 0.755 1.035 ;
        RECT  0.665 0.705 0.685 0.820 ;
        RECT  0.665 0.340 0.680 0.455 ;
        RECT  0.260 0.195 0.315 0.455 ;
        RECT  0.265 0.705 0.315 1.035 ;
    END
END INVD3BWP

MACRO INVD4BWP
    CLASS CORE ;
    FOREIGN INVD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.185 0.730 0.445 ;
        RECT  0.655 0.705 0.725 1.030 ;
        RECT  0.595 0.705 0.655 0.820 ;
        RECT  0.595 0.310 0.650 0.445 ;
        RECT  0.385 0.310 0.595 0.820 ;
        RECT  0.310 0.310 0.385 0.445 ;
        RECT  0.305 0.705 0.385 0.820 ;
        RECT  0.230 0.185 0.310 0.445 ;
        RECT  0.235 0.705 0.305 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.465 ;
        RECT  0.540 -0.115 0.830 0.115 ;
        RECT  0.420 -0.115 0.540 0.240 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.695 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.890 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.185 0.730 0.445 ;
        RECT  0.665 0.705 0.725 1.030 ;
        RECT  0.310 0.310 0.315 0.445 ;
        RECT  0.305 0.705 0.315 0.820 ;
        RECT  0.230 0.185 0.310 0.445 ;
        RECT  0.235 0.705 0.305 1.030 ;
    END
END INVD4BWP

MACRO INVD6BWP
    CLASS CORE ;
    FOREIGN INVD6BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3024 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.030 ;
        RECT  0.735 0.355 0.955 0.465 ;
        RECT  0.735 0.695 0.955 0.810 ;
        RECT  0.665 0.355 0.735 0.810 ;
        RECT  0.595 0.185 0.665 1.030 ;
        RECT  0.525 0.355 0.595 0.810 ;
        RECT  0.305 0.355 0.525 0.465 ;
        RECT  0.305 0.695 0.525 0.810 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1728 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.445 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.465 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.280 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.280 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.685 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.880 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.880 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.185 1.025 0.465 ;
        RECT  0.955 0.695 1.025 1.030 ;
        RECT  0.805 0.355 0.955 0.465 ;
        RECT  0.805 0.695 0.955 0.810 ;
        RECT  0.305 0.355 0.455 0.465 ;
        RECT  0.305 0.695 0.455 0.810 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.030 ;
        RECT  0.815 0.545 1.150 0.615 ;
    END
END INVD6BWP

MACRO INVD8BWP
    CLASS CORE ;
    FOREIGN INVD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.695 1.445 1.035 ;
        RECT  1.085 0.300 1.375 0.465 ;
        RECT  1.085 0.695 1.375 0.885 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.695 1.085 1.045 ;
        RECT  0.995 0.185 1.015 1.045 ;
        RECT  0.685 0.300 0.995 0.885 ;
        RECT  0.665 0.185 0.685 1.045 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.695 0.665 1.045 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.560 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.465 ;
        RECT  1.280 -0.115 1.550 0.115 ;
        RECT  1.160 -0.115 1.280 0.230 ;
        RECT  0.900 -0.115 1.160 0.115 ;
        RECT  0.780 -0.115 0.900 0.230 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.230 ;
        RECT  0.140 -0.115 0.400 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.695 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.160 0.955 1.280 1.375 ;
        RECT  0.900 1.145 1.160 1.375 ;
        RECT  0.780 0.955 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 0.955 0.520 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.185 1.445 0.465 ;
        RECT  1.375 0.695 1.445 1.035 ;
        RECT  1.085 0.300 1.375 0.465 ;
        RECT  1.085 0.695 1.375 0.885 ;
        RECT  0.305 0.300 0.595 0.465 ;
        RECT  0.305 0.695 0.595 0.885 ;
        RECT  0.235 0.185 0.305 0.465 ;
        RECT  0.235 0.695 0.305 1.035 ;
        RECT  1.105 0.545 1.545 0.615 ;
    END
END INVD8BWP

MACRO IOA21D0BWP
    CLASS CORE ;
    FOREIGN IOA21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0488 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.205 0.945 0.840 ;
        RECT  0.815 0.205 0.875 0.285 ;
        RECT  0.725 0.770 0.875 0.840 ;
        RECT  0.655 0.770 0.725 1.040 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.540 -0.115 0.980 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.920 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.975 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.510 0.345 0.580 0.905 ;
        RECT  0.350 0.345 0.510 0.415 ;
        RECT  0.305 0.835 0.510 0.905 ;
        RECT  0.280 0.215 0.350 0.415 ;
        RECT  0.235 0.835 0.305 1.040 ;
        RECT  0.145 0.215 0.280 0.285 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END IOA21D0BWP

MACRO IOA21D1BWP
    CLASS CORE ;
    FOREIGN IOA21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0977 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.210 0.945 0.790 ;
        RECT  0.810 0.210 0.875 0.285 ;
        RECT  0.725 0.720 0.875 0.790 ;
        RECT  0.655 0.720 0.725 1.025 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.540 -0.115 0.980 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.860 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.995 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.930 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.510 0.345 0.580 0.915 ;
        RECT  0.340 0.345 0.510 0.415 ;
        RECT  0.310 0.845 0.510 0.915 ;
        RECT  0.270 0.215 0.340 0.415 ;
        RECT  0.230 0.845 0.310 1.050 ;
        RECT  0.140 0.215 0.270 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA21D1BWP

MACRO IOA21D2BWP
    CLASS CORE ;
    FOREIGN IOA21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1582 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.845 1.050 0.915 ;
        RECT  0.805 0.355 0.870 0.425 ;
        RECT  0.735 0.355 0.805 0.915 ;
        RECT  0.665 0.845 0.735 0.915 ;
        RECT  0.595 0.845 0.665 0.965 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.140 -0.115 1.210 0.280 ;
        RECT  0.490 -0.115 1.140 0.115 ;
        RECT  0.410 -0.115 0.490 0.285 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.260 1.375 ;
        RECT  1.120 0.710 1.220 1.375 ;
        RECT  0.870 1.145 1.120 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.360 1.130 0.640 ;
        RECT  1.060 0.205 1.070 0.640 ;
        RECT  1.000 0.205 1.060 0.430 ;
        RECT  0.665 0.205 1.000 0.275 ;
        RECT  0.595 0.205 0.665 0.425 ;
        RECT  0.525 0.355 0.595 0.425 ;
        RECT  0.525 0.520 0.550 0.640 ;
        RECT  0.455 0.355 0.525 0.915 ;
        RECT  0.330 0.355 0.455 0.425 ;
        RECT  0.210 0.845 0.455 0.915 ;
        RECT  0.260 0.215 0.330 0.425 ;
        RECT  0.145 0.215 0.260 0.285 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END IOA21D2BWP

MACRO IOA21D4BWP
    CLASS CORE ;
    FOREIGN IOA21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3164 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.915 0.345 1.995 1.045 ;
        RECT  1.785 0.345 1.915 0.810 ;
        RECT  1.530 0.345 1.785 0.415 ;
        RECT  1.630 0.695 1.785 0.810 ;
        RECT  1.560 0.695 1.630 1.045 ;
        RECT  1.270 0.845 1.560 0.915 ;
        RECT  1.190 0.845 1.270 1.075 ;
        RECT  0.930 0.845 1.190 0.915 ;
        RECT  0.810 0.845 0.930 1.075 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 0.495 1.305 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.235 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.115 2.240 0.115 ;
        RECT  1.190 -0.115 1.270 0.285 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.830 -0.115 0.910 0.285 ;
        RECT  0.510 -0.115 0.830 0.115 ;
        RECT  0.430 -0.115 0.510 0.285 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.145 2.240 1.375 ;
        RECT  2.090 0.685 2.170 1.375 ;
        RECT  1.830 1.145 2.090 1.375 ;
        RECT  1.710 0.880 1.830 1.375 ;
        RECT  1.450 1.145 1.710 1.375 ;
        RECT  1.370 0.985 1.450 1.375 ;
        RECT  1.090 1.145 1.370 1.375 ;
        RECT  1.010 0.985 1.090 1.375 ;
        RECT  0.730 1.145 1.010 1.375 ;
        RECT  0.650 0.845 0.730 1.375 ;
        RECT  0.510 1.145 0.650 1.375 ;
        RECT  0.430 0.985 0.510 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.705 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.345 1.715 0.415 ;
        RECT  1.630 0.695 1.715 0.810 ;
        RECT  1.560 0.695 1.630 1.045 ;
        RECT  1.270 0.845 1.560 0.915 ;
        RECT  1.190 0.845 1.270 1.075 ;
        RECT  0.930 0.845 1.190 0.915 ;
        RECT  0.810 0.845 0.930 1.075 ;
        RECT  2.090 0.205 2.165 0.465 ;
        RECT  1.450 0.205 2.090 0.275 ;
        RECT  1.480 0.545 1.705 0.615 ;
        RECT  1.410 0.545 1.480 0.775 ;
        RECT  1.375 0.205 1.450 0.425 ;
        RECT  0.555 0.705 1.410 0.775 ;
        RECT  1.085 0.355 1.375 0.425 ;
        RECT  1.015 0.190 1.085 0.425 ;
        RECT  0.485 0.355 0.555 0.905 ;
        RECT  0.350 0.355 0.485 0.425 ;
        RECT  0.340 0.835 0.485 0.905 ;
        RECT  0.280 0.215 0.350 0.425 ;
        RECT  0.240 0.835 0.340 1.075 ;
        RECT  0.160 0.215 0.280 0.285 ;
        RECT  0.060 0.185 0.160 0.285 ;
        RECT  0.740 0.355 1.015 0.425 ;
        RECT  0.640 0.185 0.740 0.425 ;
    END
END IOA21D4BWP

MACRO IOA22D0BWP
    CLASS CORE ;
    FOREIGN IOA22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0621 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.975 1.220 1.075 ;
        RECT  1.030 0.975 1.120 1.045 ;
        RECT  0.960 0.845 1.030 1.045 ;
        RECT  0.710 0.845 0.960 0.915 ;
        RECT  0.665 0.195 0.710 0.915 ;
        RECT  0.640 0.195 0.665 1.045 ;
        RECT  0.595 0.195 0.640 0.315 ;
        RECT  0.595 0.775 0.640 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.635 1.225 0.905 ;
        RECT  1.040 0.635 1.135 0.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.115 1.260 0.115 ;
        RECT  0.930 -0.115 1.050 0.285 ;
        RECT  0.510 -0.115 0.930 0.115 ;
        RECT  0.390 -0.115 0.510 0.285 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 1.145 1.260 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.975 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.195 1.205 0.425 ;
        RECT  0.850 0.355 1.135 0.425 ;
        RECT  0.780 0.195 0.850 0.425 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.905 ;
        RECT  0.300 0.355 0.455 0.425 ;
        RECT  0.305 0.835 0.455 0.905 ;
        RECT  0.235 0.835 0.305 1.050 ;
        RECT  0.230 0.215 0.300 0.425 ;
        RECT  0.140 0.215 0.230 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA22D0BWP

MACRO IOA22D1BWP
    CLASS CORE ;
    FOREIGN IOA22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1243 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.975 1.225 1.075 ;
        RECT  1.020 0.975 1.120 1.045 ;
        RECT  0.950 0.845 1.020 1.045 ;
        RECT  0.700 0.845 0.950 0.915 ;
        RECT  0.665 0.185 0.700 0.915 ;
        RECT  0.630 0.185 0.665 1.055 ;
        RECT  0.595 0.185 0.630 0.450 ;
        RECT  0.595 0.775 0.630 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.225 0.905 ;
        RECT  1.040 0.545 1.135 0.615 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.115 1.260 0.115 ;
        RECT  0.950 -0.115 1.030 0.285 ;
        RECT  0.490 -0.115 0.950 0.115 ;
        RECT  0.410 -0.115 0.490 0.285 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 1.145 1.260 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.975 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.935 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.120 0.185 1.220 0.425 ;
        RECT  0.850 0.355 1.120 0.425 ;
        RECT  0.770 0.265 0.850 0.425 ;
        RECT  0.525 0.520 0.560 0.640 ;
        RECT  0.455 0.355 0.525 0.905 ;
        RECT  0.300 0.355 0.455 0.425 ;
        RECT  0.310 0.835 0.455 0.905 ;
        RECT  0.230 0.835 0.310 1.055 ;
        RECT  0.230 0.215 0.300 0.425 ;
        RECT  0.145 0.215 0.230 0.285 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END IOA22D1BWP

MACRO IOA22D2BWP
    CLASS CORE ;
    FOREIGN IOA22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.195 1.085 0.800 ;
        RECT  0.930 0.195 1.015 0.275 ;
        RECT  0.930 0.720 1.015 0.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.270 0.645 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.520 1.645 0.905 ;
        RECT  1.490 0.520 1.555 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.310 ;
        RECT  1.235 -0.115 1.550 0.115 ;
        RECT  1.165 -0.115 1.235 0.310 ;
        RECT  0.850 -0.115 1.165 0.115 ;
        RECT  0.770 -0.115 0.850 0.285 ;
        RECT  0.670 -0.115 0.770 0.115 ;
        RECT  0.590 -0.115 0.670 0.285 ;
        RECT  0.140 -0.115 0.590 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.145 1.680 1.375 ;
        RECT  1.150 1.010 1.250 1.375 ;
        RECT  0.865 1.145 1.150 1.375 ;
        RECT  0.755 1.010 0.865 1.375 ;
        RECT  0.310 1.145 0.755 1.375 ;
        RECT  0.230 0.975 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.975 1.640 1.075 ;
        RECT  1.420 0.975 1.540 1.045 ;
        RECT  1.420 0.205 1.470 0.275 ;
        RECT  1.350 0.205 1.420 1.045 ;
        RECT  0.805 0.870 1.350 0.940 ;
        RECT  0.875 0.355 0.945 0.640 ;
        RECT  0.545 0.355 0.875 0.425 ;
        RECT  0.735 0.545 0.805 0.940 ;
        RECT  0.625 0.545 0.735 0.615 ;
        RECT  0.595 0.695 0.665 1.055 ;
        RECT  0.545 0.695 0.595 0.765 ;
        RECT  0.500 0.355 0.545 0.765 ;
        RECT  0.475 0.185 0.500 0.765 ;
        RECT  0.400 0.835 0.500 1.075 ;
        RECT  0.400 0.185 0.475 0.425 ;
        RECT  0.130 0.835 0.400 0.905 ;
        RECT  0.050 0.765 0.130 1.045 ;
    END
END IOA22D2BWP

MACRO IOA22D4BWP
    CLASS CORE ;
    FOREIGN IOA22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 0.465 ;
        RECT  1.855 0.680 1.925 0.800 ;
        RECT  1.645 0.355 1.855 0.800 ;
        RECT  1.575 0.355 1.645 0.465 ;
        RECT  1.480 0.680 1.645 0.800 ;
        RECT  1.495 0.185 1.575 0.465 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.470 2.205 0.790 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.485 0.625 ;
        RECT  2.300 0.545 2.415 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.385 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 -0.115 2.520 0.115 ;
        RECT  2.380 -0.115 2.480 0.275 ;
        RECT  2.130 -0.115 2.380 0.115 ;
        RECT  2.010 -0.115 2.130 0.250 ;
        RECT  1.750 -0.115 2.010 0.115 ;
        RECT  1.670 -0.115 1.750 0.280 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.285 ;
        RECT  1.030 -0.115 1.310 0.115 ;
        RECT  0.950 -0.115 1.030 0.285 ;
        RECT  0.310 -0.115 0.950 0.115 ;
        RECT  0.230 -0.115 0.310 0.285 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.145 2.520 1.375 ;
        RECT  2.010 1.010 2.130 1.375 ;
        RECT  1.770 1.145 2.010 1.375 ;
        RECT  1.650 1.010 1.770 1.375 ;
        RECT  1.410 1.145 1.650 1.375 ;
        RECT  1.290 1.010 1.410 1.375 ;
        RECT  0.670 1.145 1.290 1.375 ;
        RECT  0.590 0.855 0.670 1.375 ;
        RECT  0.310 1.145 0.590 1.375 ;
        RECT  0.230 0.855 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.495 0.185 1.575 0.465 ;
        RECT  1.480 0.680 1.575 0.800 ;
        RECT  2.390 0.745 2.470 1.025 ;
        RECT  2.065 0.870 2.390 0.940 ;
        RECT  2.210 0.185 2.290 0.390 ;
        RECT  2.065 0.320 2.210 0.390 ;
        RECT  1.995 0.320 2.065 0.940 ;
        RECT  1.380 0.870 1.995 0.940 ;
        RECT  1.375 0.540 1.500 0.610 ;
        RECT  1.310 0.690 1.380 0.940 ;
        RECT  1.305 0.355 1.375 0.610 ;
        RECT  1.225 0.690 1.310 0.760 ;
        RECT  1.210 0.355 1.305 0.425 ;
        RECT  1.155 0.510 1.225 0.760 ;
        RECT  1.130 0.190 1.210 0.425 ;
        RECT  1.130 0.830 1.210 1.065 ;
        RECT  1.025 0.355 1.130 0.425 ;
        RECT  0.845 0.995 1.130 1.065 ;
        RECT  0.955 0.355 1.025 0.925 ;
        RECT  0.570 0.355 0.955 0.425 ;
        RECT  0.490 0.205 0.870 0.275 ;
        RECT  0.775 0.705 0.845 1.065 ;
        RECT  0.485 0.705 0.775 0.785 ;
        RECT  0.410 0.205 0.490 0.425 ;
        RECT  0.415 0.705 0.485 1.035 ;
        RECT  0.125 0.705 0.415 0.785 ;
        RECT  0.140 0.355 0.410 0.425 ;
        RECT  0.040 0.185 0.140 0.425 ;
        RECT  0.055 0.705 0.125 1.035 ;
    END
END IOA22D4BWP

MACRO ISOHID1BWP
    CLASS CORE ;
    FOREIGN ISOHID1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.700 0.185 0.735 0.465 ;
        RECT  0.700 0.750 0.735 1.045 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.210 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 -0.115 0.840 0.115 ;
        RECT  0.470 -0.115 0.590 0.275 ;
        RECT  0.160 -0.115 0.470 0.115 ;
        RECT  0.060 -0.115 0.160 0.275 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.460 0.990 0.580 1.375 ;
        RECT  0.000 1.145 0.460 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.650 0.640 ;
        RECT  0.515 0.345 0.585 0.915 ;
        RECT  0.330 0.345 0.515 0.415 ;
        RECT  0.150 0.845 0.515 0.915 ;
        RECT  0.250 0.245 0.330 0.415 ;
        RECT  0.070 0.845 0.150 1.015 ;
    END
END ISOHID1BWP

MACRO ISOHID2BWP
    CLASS CORE ;
    FOREIGN ISOHID2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.745 0.355 0.805 0.820 ;
        RECT  0.735 0.185 0.745 1.045 ;
        RECT  0.675 0.185 0.735 0.465 ;
        RECT  0.675 0.750 0.735 1.045 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.300 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.275 ;
        RECT  0.145 -0.115 0.440 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.910 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.990 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.585 0.520 0.630 0.640 ;
        RECT  0.515 0.345 0.585 0.915 ;
        RECT  0.320 0.345 0.515 0.415 ;
        RECT  0.130 0.845 0.515 0.915 ;
        RECT  0.240 0.245 0.320 0.415 ;
        RECT  0.050 0.845 0.130 1.015 ;
    END
END ISOHID2BWP

MACRO ISOHID4BWP
    CLASS CORE ;
    FOREIGN ISOHID4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.025 0.465 ;
        RECT  1.015 0.755 1.025 1.045 ;
        RECT  0.955 0.185 1.015 1.045 ;
        RECT  0.805 0.355 0.955 0.905 ;
        RECT  0.665 0.355 0.805 0.465 ;
        RECT  0.665 0.755 0.805 0.905 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.755 0.665 1.045 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 0.495 0.385 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.475 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.145 -0.115 0.390 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.675 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.990 0.510 1.375 ;
        RECT  0.000 1.145 0.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.355 0.735 0.465 ;
        RECT  0.665 0.755 0.735 0.905 ;
        RECT  0.595 0.185 0.665 0.465 ;
        RECT  0.595 0.755 0.665 1.045 ;
        RECT  0.525 0.545 0.645 0.615 ;
        RECT  0.455 0.345 0.525 0.915 ;
        RECT  0.310 0.345 0.455 0.415 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.230 0.245 0.310 0.415 ;
        RECT  0.050 0.845 0.130 1.015 ;
    END
END ISOHID4BWP

MACRO ISOHID8BWP
    CLASS CORE ;
    FOREIGN ISOHID8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.725 2.590 0.955 ;
        RECT  2.185 0.320 2.570 0.440 ;
        RECT  2.135 0.185 2.185 0.440 ;
        RECT  2.115 0.185 2.135 0.955 ;
        RECT  1.925 0.320 2.115 0.955 ;
        RECT  1.805 0.320 1.925 0.440 ;
        RECT  1.350 0.725 1.925 0.955 ;
        RECT  1.735 0.185 1.805 0.440 ;
        RECT  1.350 0.320 1.735 0.440 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.495 1.130 0.640 ;
        RECT  1.015 0.495 1.095 0.770 ;
        RECT  0.535 0.700 1.015 0.770 ;
        RECT  0.445 0.495 0.535 0.770 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.545 0.875 0.625 ;
        RECT  0.735 0.350 0.805 0.625 ;
        RECT  0.280 0.350 0.735 0.420 ;
        RECT  0.210 0.350 0.280 0.615 ;
        RECT  0.100 0.545 0.210 0.615 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.465 ;
        RECT  2.400 -0.115 2.670 0.115 ;
        RECT  2.280 -0.115 2.400 0.250 ;
        RECT  2.020 -0.115 2.280 0.115 ;
        RECT  1.900 -0.115 2.020 0.250 ;
        RECT  1.640 -0.115 1.900 0.115 ;
        RECT  1.520 -0.115 1.640 0.250 ;
        RECT  1.270 -0.115 1.520 0.115 ;
        RECT  1.150 -0.115 1.270 0.275 ;
        RECT  0.900 -0.115 1.150 0.115 ;
        RECT  0.780 -0.115 0.900 0.140 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.140 ;
        RECT  0.125 -0.115 0.400 0.115 ;
        RECT  0.055 -0.115 0.125 0.465 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.675 2.750 1.375 ;
        RECT  2.400 1.145 2.670 1.375 ;
        RECT  2.280 1.025 2.400 1.375 ;
        RECT  2.020 1.145 2.280 1.375 ;
        RECT  1.900 1.025 2.020 1.375 ;
        RECT  1.640 1.145 1.900 1.375 ;
        RECT  1.520 1.025 1.640 1.375 ;
        RECT  1.270 1.145 1.520 1.375 ;
        RECT  1.150 0.990 1.270 1.375 ;
        RECT  0.520 1.145 1.150 1.375 ;
        RECT  0.400 0.990 0.520 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.725 2.590 0.955 ;
        RECT  1.350 0.320 1.735 0.440 ;
        RECT  2.235 0.545 2.630 0.615 ;
        RECT  1.270 0.545 1.825 0.615 ;
        RECT  1.200 0.345 1.270 0.910 ;
        RECT  1.065 0.345 1.200 0.415 ;
        RECT  0.880 0.840 1.200 0.910 ;
        RECT  0.995 0.210 1.065 0.415 ;
        RECT  0.210 0.210 0.995 0.280 ;
        RECT  0.800 0.840 0.880 1.075 ;
        RECT  0.125 0.840 0.800 0.910 ;
        RECT  0.055 0.730 0.125 1.030 ;
        RECT  2.205 0.320 2.570 0.440 ;
        RECT  1.805 0.320 1.855 0.440 ;
        RECT  1.350 0.725 1.855 0.955 ;
        RECT  1.735 0.185 1.805 0.440 ;
    END
END ISOHID8BWP

MACRO ISOLOD1BWP
    CLASS CORE ;
    FOREIGN ISOLOD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.195 1.085 1.070 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.530 0.600 0.630 ;
        RECT  0.455 0.355 0.525 0.630 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 1.120 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.340 -0.115 0.790 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.145 1.120 1.375 ;
        RECT  0.810 0.885 0.890 1.375 ;
        RECT  0.710 1.145 0.810 1.375 ;
        RECT  0.630 0.885 0.710 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.845 0.380 0.915 0.805 ;
        RECT  0.720 0.380 0.845 0.450 ;
        RECT  0.525 0.735 0.845 0.805 ;
        RECT  0.620 0.210 0.720 0.450 ;
        RECT  0.455 0.735 0.525 1.045 ;
        RECT  0.305 0.345 0.375 0.915 ;
        RECT  0.130 0.345 0.305 0.415 ;
        RECT  0.130 0.845 0.305 0.915 ;
        RECT  0.050 0.205 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END ISOLOD1BWP

MACRO ISOLOD2BWP
    CLASS CORE ;
    FOREIGN ISOLOD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.355 1.085 0.820 ;
        RECT  1.015 0.185 1.025 1.045 ;
        RECT  0.955 0.185 1.015 0.465 ;
        RECT  0.955 0.750 1.015 1.045 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.530 0.570 0.630 ;
        RECT  0.455 0.355 0.525 0.630 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.280 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.330 -0.115 0.750 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.910 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.885 0.850 1.375 ;
        RECT  0.670 1.145 0.770 1.375 ;
        RECT  0.590 0.885 0.670 1.375 ;
        RECT  0.330 1.145 0.590 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.800 0.380 0.875 0.805 ;
        RECT  0.665 0.380 0.800 0.450 ;
        RECT  0.485 0.735 0.800 0.805 ;
        RECT  0.595 0.190 0.665 0.450 ;
        RECT  0.415 0.735 0.485 1.045 ;
        RECT  0.335 0.520 0.375 0.640 ;
        RECT  0.265 0.345 0.335 0.915 ;
        RECT  0.130 0.345 0.265 0.415 ;
        RECT  0.130 0.845 0.265 0.915 ;
        RECT  0.050 0.205 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END ISOLOD2BWP

MACRO ISOLOD4BWP
    CLASS CORE ;
    FOREIGN ISOLOD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.445 0.465 ;
        RECT  1.435 0.755 1.445 1.045 ;
        RECT  1.375 0.185 1.435 1.045 ;
        RECT  1.225 0.345 1.375 0.905 ;
        RECT  1.085 0.345 1.225 0.465 ;
        RECT  1.085 0.755 1.225 0.905 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.755 1.085 1.045 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.645 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.495 0.665 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.475 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.275 ;
        RECT  0.930 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.930 0.270 ;
        RECT  0.360 -0.115 0.810 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.675 1.630 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.985 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.730 1.145 0.830 1.375 ;
        RECT  0.650 0.980 0.730 1.375 ;
        RECT  0.360 1.145 0.650 1.375 ;
        RECT  0.240 0.985 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.345 1.155 0.465 ;
        RECT  1.085 0.755 1.155 0.905 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.755 1.085 1.045 ;
        RECT  0.870 0.545 1.080 0.615 ;
        RECT  0.800 0.345 0.870 0.905 ;
        RECT  0.630 0.345 0.800 0.415 ;
        RECT  0.545 0.835 0.800 0.905 ;
        RECT  0.475 0.835 0.545 1.045 ;
        RECT  0.380 0.520 0.435 0.640 ;
        RECT  0.310 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.310 0.415 ;
        RECT  0.130 0.845 0.310 0.915 ;
        RECT  0.050 0.205 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END ISOLOD4BWP

MACRO ISOLOD8BWP
    CLASS CORE ;
    FOREIGN ISOLOD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.775 0.690 2.845 0.970 ;
        RECT  2.485 0.345 2.775 0.465 ;
        RECT  2.485 0.690 2.775 0.820 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.690 2.485 0.970 ;
        RECT  2.205 0.345 2.415 0.820 ;
        RECT  2.125 0.345 2.205 0.465 ;
        RECT  2.125 0.690 2.205 0.820 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.690 2.125 0.970 ;
        RECT  1.765 0.345 2.055 0.465 ;
        RECT  1.765 0.690 2.055 0.820 ;
        RECT  1.695 0.185 1.765 0.465 ;
        RECT  1.695 0.690 1.765 0.970 ;
        END
    END Z
    PIN ISO
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END ISO
    PIN I
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.290 0.640 ;
        RECT  1.155 0.495 1.225 0.770 ;
        RECT  0.665 0.700 1.155 0.770 ;
        RECT  0.595 0.495 0.665 0.770 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.475 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.275 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.275 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.275 ;
        RECT  1.590 -0.115 1.850 0.115 ;
        RECT  1.510 -0.115 1.590 0.465 ;
        RECT  1.060 -0.115 1.510 0.115 ;
        RECT  0.940 -0.115 1.060 0.140 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.675 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 0.890 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 0.890 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 0.890 1.970 1.375 ;
        RECT  1.590 1.145 1.850 1.375 ;
        RECT  1.510 0.765 1.590 1.375 ;
        RECT  1.430 1.145 1.510 1.375 ;
        RECT  1.310 0.990 1.430 1.375 ;
        RECT  1.060 1.145 1.310 1.375 ;
        RECT  0.940 0.990 1.060 1.375 ;
        RECT  0.690 1.145 0.940 1.375 ;
        RECT  0.570 0.990 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.775 0.185 2.845 0.465 ;
        RECT  2.775 0.690 2.845 0.970 ;
        RECT  2.485 0.345 2.775 0.465 ;
        RECT  2.485 0.690 2.775 0.820 ;
        RECT  2.125 0.345 2.135 0.465 ;
        RECT  2.125 0.690 2.135 0.820 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  2.055 0.690 2.125 0.970 ;
        RECT  1.765 0.345 2.055 0.465 ;
        RECT  1.765 0.690 2.055 0.820 ;
        RECT  1.695 0.185 1.765 0.465 ;
        RECT  1.695 0.690 1.765 0.970 ;
        RECT  2.515 0.545 2.900 0.615 ;
        RECT  1.440 0.545 2.105 0.615 ;
        RECT  1.370 0.210 1.440 0.910 ;
        RECT  0.570 0.210 1.370 0.280 ;
        RECT  1.230 0.840 1.370 0.910 ;
        RECT  1.150 0.840 1.230 1.075 ;
        RECT  0.850 0.840 1.150 0.910 ;
        RECT  0.945 0.545 1.050 0.615 ;
        RECT  0.865 0.350 0.945 0.615 ;
        RECT  0.515 0.350 0.865 0.420 ;
        RECT  0.770 0.840 0.850 1.075 ;
        RECT  0.490 0.840 0.770 0.910 ;
        RECT  0.445 0.350 0.515 0.615 ;
        RECT  0.410 0.745 0.490 1.045 ;
        RECT  0.330 0.545 0.445 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.130 0.345 0.260 0.415 ;
        RECT  0.130 0.845 0.260 0.915 ;
        RECT  0.050 0.245 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END ISOLOD8BWP

MACRO LHCND1BWP
    CLASS CORE ;
    FOREIGN LHCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.710 2.290 0.780 ;
        RECT  2.205 0.185 2.245 0.465 ;
        RECT  2.135 0.185 2.205 0.780 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.195 2.625 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.115 2.660 0.115 ;
        RECT  2.350 -0.115 2.430 0.440 ;
        RECT  2.065 -0.115 2.350 0.115 ;
        RECT  1.990 -0.115 2.065 0.300 ;
        RECT  1.530 -0.115 1.990 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.145 2.660 1.375 ;
        RECT  2.340 0.990 2.440 1.375 ;
        RECT  2.080 1.145 2.340 1.375 ;
        RECT  1.980 0.990 2.080 1.375 ;
        RECT  1.520 1.145 1.980 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.380 0.520 2.460 0.920 ;
        RECT  1.970 0.850 2.380 0.920 ;
        RECT  1.900 0.380 1.970 0.920 ;
        RECT  1.890 0.380 1.900 0.465 ;
        RECT  1.890 0.720 1.900 0.920 ;
        RECT  1.810 0.185 1.890 0.465 ;
        RECT  1.810 0.720 1.890 1.040 ;
        RECT  1.715 0.545 1.830 0.615 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCND1BWP

MACRO LHCND2BWP
    CLASS CORE ;
    FOREIGN LHCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.710 2.290 0.780 ;
        RECT  2.205 0.185 2.245 0.465 ;
        RECT  2.135 0.185 2.205 0.780 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.355 2.765 0.765 ;
        RECT  2.695 0.185 2.700 1.045 ;
        RECT  2.620 0.185 2.695 0.470 ;
        RECT  2.620 0.695 2.695 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.300 ;
        RECT  2.490 -0.115 2.810 0.115 ;
        RECT  2.390 -0.115 2.490 0.440 ;
        RECT  2.065 -0.115 2.390 0.115 ;
        RECT  1.990 -0.115 2.065 0.300 ;
        RECT  1.530 -0.115 1.990 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.845 2.890 1.375 ;
        RECT  2.490 1.145 2.810 1.375 ;
        RECT  2.390 0.990 2.490 1.375 ;
        RECT  2.080 1.145 2.390 1.375 ;
        RECT  1.980 0.990 2.080 1.375 ;
        RECT  1.520 1.145 1.980 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.460 0.540 2.610 0.620 ;
        RECT  2.380 0.540 2.460 0.920 ;
        RECT  1.970 0.850 2.380 0.920 ;
        RECT  1.900 0.380 1.970 0.920 ;
        RECT  1.890 0.380 1.900 0.465 ;
        RECT  1.890 0.720 1.900 0.920 ;
        RECT  1.810 0.185 1.890 0.465 ;
        RECT  1.810 0.720 1.890 1.040 ;
        RECT  1.715 0.545 1.830 0.615 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCND2BWP

MACRO LHCND4BWP
    CLASS CORE ;
    FOREIGN LHCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.700 2.850 0.800 ;
        RECT  2.755 0.185 2.825 0.485 ;
        RECT  2.695 0.355 2.755 0.485 ;
        RECT  2.485 0.355 2.695 0.800 ;
        RECT  2.465 0.355 2.485 0.485 ;
        RECT  2.370 0.700 2.485 0.800 ;
        RECT  2.395 0.185 2.465 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.545 0.465 ;
        RECT  3.535 0.735 3.545 1.035 ;
        RECT  3.475 0.185 3.535 1.035 ;
        RECT  3.325 0.355 3.475 0.905 ;
        RECT  3.185 0.355 3.325 0.465 ;
        RECT  3.185 0.735 3.325 0.905 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.735 3.185 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.460 ;
        RECT  3.380 -0.115 3.650 0.115 ;
        RECT  3.280 -0.115 3.380 0.275 ;
        RECT  3.010 -0.115 3.280 0.115 ;
        RECT  2.930 -0.115 3.010 0.460 ;
        RECT  2.660 -0.115 2.930 0.115 ;
        RECT  2.560 -0.115 2.660 0.275 ;
        RECT  2.290 -0.115 2.560 0.115 ;
        RECT  2.210 -0.115 2.290 0.320 ;
        RECT  1.900 -0.115 2.210 0.115 ;
        RECT  1.820 -0.115 1.900 0.460 ;
        RECT  1.530 -0.115 1.820 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.665 3.730 1.375 ;
        RECT  3.380 1.145 3.650 1.375 ;
        RECT  3.280 0.985 3.380 1.375 ;
        RECT  3.030 1.145 3.280 1.375 ;
        RECT  2.910 1.010 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.010 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.010 2.310 1.375 ;
        RECT  1.920 1.145 2.190 1.375 ;
        RECT  1.840 0.745 1.920 1.375 ;
        RECT  1.520 1.145 1.840 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.355 3.255 0.465 ;
        RECT  3.185 0.735 3.255 0.905 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.735 3.185 1.035 ;
        RECT  2.765 0.700 2.850 0.800 ;
        RECT  2.765 0.185 2.825 0.485 ;
        RECT  2.395 0.185 2.415 0.485 ;
        RECT  2.370 0.700 2.415 0.800 ;
        RECT  3.000 0.540 3.230 0.620 ;
        RECT  2.930 0.540 3.000 0.940 ;
        RECT  2.170 0.870 2.930 0.940 ;
        RECT  2.110 0.395 2.170 0.940 ;
        RECT  2.100 0.185 2.110 1.065 ;
        RECT  2.030 0.185 2.100 0.465 ;
        RECT  2.030 0.745 2.100 1.065 ;
        RECT  1.730 0.540 2.020 0.620 ;
        RECT  1.725 0.540 1.730 1.060 ;
        RECT  1.650 0.185 1.725 1.060 ;
        RECT  1.630 0.185 1.650 0.465 ;
        RECT  1.370 0.990 1.650 1.060 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCND4BWP

MACRO LHCNDD1BWP
    CLASS CORE ;
    FOREIGN LHCNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.710 2.570 0.780 ;
        RECT  2.485 0.185 2.525 0.465 ;
        RECT  2.415 0.185 2.485 0.780 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.815 0.195 2.905 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.110 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.940 0.115 ;
        RECT  2.630 -0.115 2.710 0.440 ;
        RECT  2.345 -0.115 2.630 0.115 ;
        RECT  2.270 -0.115 2.345 0.300 ;
        RECT  1.810 -0.115 2.270 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 2.940 1.375 ;
        RECT  2.620 0.990 2.720 1.375 ;
        RECT  2.360 1.145 2.620 1.375 ;
        RECT  2.260 0.990 2.360 1.375 ;
        RECT  1.800 1.145 2.260 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.520 2.740 0.920 ;
        RECT  2.250 0.850 2.660 0.920 ;
        RECT  2.180 0.380 2.250 0.920 ;
        RECT  2.170 0.380 2.180 0.465 ;
        RECT  2.170 0.720 2.180 0.920 ;
        RECT  2.090 0.185 2.170 0.465 ;
        RECT  2.090 0.720 2.170 1.040 ;
        RECT  1.995 0.545 2.110 0.615 ;
        RECT  1.925 0.185 1.995 1.060 ;
        RECT  1.915 0.185 1.925 0.465 ;
        RECT  1.915 0.730 1.925 1.060 ;
        RECT  1.650 0.985 1.915 1.060 ;
        RECT  1.830 0.520 1.855 0.640 ;
        RECT  1.760 0.210 1.830 0.915 ;
        RECT  1.110 0.210 1.760 0.280 ;
        RECT  0.590 0.845 1.760 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.440 0.260 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHCNDD1BWP

MACRO LHCNDD2BWP
    CLASS CORE ;
    FOREIGN LHCNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.185 2.490 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.055 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.735 2.835 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.115 3.080 0.115 ;
        RECT  2.955 -0.115 3.025 0.305 ;
        RECT  2.670 -0.115 2.955 0.115 ;
        RECT  2.590 -0.115 2.670 0.465 ;
        RECT  2.310 -0.115 2.590 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.780 -0.115 2.230 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 1.145 3.080 1.375 ;
        RECT  2.955 0.960 3.025 1.375 ;
        RECT  2.690 1.145 2.955 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  0.910 1.145 2.210 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.615 ;
        RECT  2.595 0.545 2.665 0.935 ;
        RECT  2.240 0.865 2.595 0.935 ;
        RECT  2.170 0.385 2.240 0.935 ;
        RECT  2.130 0.385 2.170 0.465 ;
        RECT  2.130 0.735 2.170 0.935 ;
        RECT  2.050 0.185 2.130 0.465 ;
        RECT  2.050 0.735 2.130 1.055 ;
        RECT  1.955 0.545 2.100 0.620 ;
        RECT  1.885 0.185 1.955 1.055 ;
        RECT  1.875 0.185 1.885 0.465 ;
        RECT  1.875 0.775 1.885 1.055 ;
        RECT  1.670 0.985 1.875 1.055 ;
        RECT  1.795 0.520 1.815 0.640 ;
        RECT  1.725 0.205 1.795 0.915 ;
        RECT  1.090 0.205 1.725 0.275 ;
        RECT  0.590 0.845 1.725 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.195 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCNDD2BWP

MACRO LHCNDD4BWP
    CLASS CORE ;
    FOREIGN LHCNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.705 3.130 0.795 ;
        RECT  3.035 0.185 3.105 0.485 ;
        RECT  2.975 0.355 3.035 0.485 ;
        RECT  2.765 0.355 2.975 0.795 ;
        RECT  2.745 0.355 2.765 0.485 ;
        RECT  2.650 0.705 2.765 0.795 ;
        RECT  2.675 0.185 2.745 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.825 0.465 ;
        RECT  3.815 0.775 3.825 1.055 ;
        RECT  3.755 0.185 3.815 1.055 ;
        RECT  3.605 0.355 3.755 0.905 ;
        RECT  3.465 0.355 3.605 0.465 ;
        RECT  3.465 0.775 3.605 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.345 1.660 0.485 ;
        RECT  0.665 0.345 1.580 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.485 ;
        RECT  3.670 -0.115 3.930 0.115 ;
        RECT  3.550 -0.115 3.670 0.275 ;
        RECT  3.290 -0.115 3.550 0.115 ;
        RECT  3.210 -0.115 3.290 0.465 ;
        RECT  2.950 -0.115 3.210 0.115 ;
        RECT  2.830 -0.115 2.950 0.275 ;
        RECT  2.570 -0.115 2.830 0.115 ;
        RECT  2.490 -0.115 2.570 0.305 ;
        RECT  2.200 -0.115 2.490 0.115 ;
        RECT  2.120 -0.115 2.200 0.465 ;
        RECT  1.800 -0.115 2.120 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.680 -0.115 1.680 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.665 4.010 1.375 ;
        RECT  3.670 1.145 3.930 1.375 ;
        RECT  3.550 0.985 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 1.005 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 1.005 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 1.005 2.590 1.375 ;
        RECT  2.200 1.145 2.470 1.375 ;
        RECT  2.120 0.755 2.200 1.375 ;
        RECT  1.800 1.145 2.120 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.355 3.535 0.465 ;
        RECT  3.465 0.775 3.535 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        RECT  3.045 0.705 3.130 0.795 ;
        RECT  3.045 0.185 3.105 0.485 ;
        RECT  2.675 0.185 2.695 0.485 ;
        RECT  2.650 0.705 2.695 0.795 ;
        RECT  3.285 0.540 3.515 0.620 ;
        RECT  3.215 0.540 3.285 0.935 ;
        RECT  2.530 0.865 3.215 0.935 ;
        RECT  2.460 0.385 2.530 0.935 ;
        RECT  2.390 0.385 2.460 0.465 ;
        RECT  2.390 0.735 2.460 0.935 ;
        RECT  2.310 0.185 2.390 0.465 ;
        RECT  2.310 0.735 2.390 1.055 ;
        RECT  2.050 0.545 2.380 0.620 ;
        RECT  1.980 0.280 2.050 1.055 ;
        RECT  1.920 0.280 1.980 0.440 ;
        RECT  1.930 0.775 1.980 1.055 ;
        RECT  1.650 0.985 1.930 1.055 ;
        RECT  1.840 0.520 1.910 0.640 ;
        RECT  1.770 0.205 1.840 0.915 ;
        RECT  1.090 0.205 1.770 0.275 ;
        RECT  0.590 0.845 1.770 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCNDD4BWP

MACRO LHCNDQD1BWP
    CLASS CORE ;
    FOREIGN LHCNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.625 1.055 ;
        RECT  2.535 0.185 2.555 0.465 ;
        RECT  2.535 0.775 2.555 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.110 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.115 2.660 0.115 ;
        RECT  2.320 -0.115 2.400 0.305 ;
        RECT  1.810 -0.115 2.320 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 1.145 2.660 1.375 ;
        RECT  2.320 0.925 2.400 1.375 ;
        RECT  1.800 1.145 2.320 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.465 0.520 2.485 0.640 ;
        RECT  2.395 0.385 2.465 0.805 ;
        RECT  2.185 0.385 2.395 0.465 ;
        RECT  2.190 0.735 2.395 0.805 ;
        RECT  1.990 0.545 2.290 0.615 ;
        RECT  2.110 0.735 2.190 1.055 ;
        RECT  2.115 0.185 2.185 0.465 ;
        RECT  1.915 0.195 1.990 1.060 ;
        RECT  1.650 0.985 1.915 1.060 ;
        RECT  1.775 0.210 1.845 0.915 ;
        RECT  1.110 0.210 1.775 0.280 ;
        RECT  0.590 0.845 1.775 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.440 0.260 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHCNDQD1BWP

MACRO LHCNDQD2BWP
    CLASS CORE ;
    FOREIGN LHCNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.355 2.625 0.905 ;
        RECT  2.565 0.355 2.570 1.055 ;
        RECT  2.555 0.185 2.565 1.055 ;
        RECT  2.490 0.185 2.555 0.465 ;
        RECT  2.490 0.735 2.555 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.345 1.660 0.485 ;
        RECT  0.665 0.345 1.580 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.745 -0.115 2.800 0.115 ;
        RECT  2.675 -0.115 2.745 0.305 ;
        RECT  2.360 -0.115 2.675 0.115 ;
        RECT  2.280 -0.115 2.360 0.305 ;
        RECT  1.800 -0.115 2.280 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.680 -0.115 1.680 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.745 1.145 2.800 1.375 ;
        RECT  2.675 0.960 2.745 1.375 ;
        RECT  2.360 1.145 2.675 1.375 ;
        RECT  2.280 0.915 2.360 1.375 ;
        RECT  1.800 1.145 2.280 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.420 0.520 2.440 0.640 ;
        RECT  2.350 0.385 2.420 0.805 ;
        RECT  2.165 0.385 2.350 0.465 ;
        RECT  2.170 0.735 2.350 0.805 ;
        RECT  1.990 0.545 2.270 0.620 ;
        RECT  2.090 0.735 2.170 1.055 ;
        RECT  2.095 0.185 2.165 0.465 ;
        RECT  1.910 0.195 1.990 1.055 ;
        RECT  1.650 0.985 1.910 1.055 ;
        RECT  1.770 0.205 1.840 0.915 ;
        RECT  1.090 0.205 1.770 0.275 ;
        RECT  0.590 0.845 1.770 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.195 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCNDQD2BWP

MACRO LHCNDQD4BWP
    CLASS CORE ;
    FOREIGN LHCNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.775 3.125 1.055 ;
        RECT  3.055 0.185 3.115 1.055 ;
        RECT  2.905 0.355 3.055 0.905 ;
        RECT  2.765 0.355 2.905 0.465 ;
        RECT  2.765 0.775 2.905 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.345 1.660 0.485 ;
        RECT  0.665 0.345 1.580 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.485 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.275 ;
        RECT  2.560 -0.115 2.850 0.115 ;
        RECT  2.475 -0.115 2.560 0.305 ;
        RECT  2.170 -0.115 2.475 0.115 ;
        RECT  2.090 -0.115 2.170 0.465 ;
        RECT  1.800 -0.115 2.090 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.680 -0.115 1.680 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.665 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.985 2.970 1.375 ;
        RECT  2.560 1.145 2.850 1.375 ;
        RECT  2.480 0.925 2.560 1.375 ;
        RECT  2.170 1.145 2.480 1.375 ;
        RECT  2.090 0.755 2.170 1.375 ;
        RECT  1.800 1.145 2.090 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.465 ;
        RECT  2.765 0.775 2.835 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        RECT  2.625 0.545 2.815 0.620 ;
        RECT  2.555 0.385 2.625 0.845 ;
        RECT  2.360 0.385 2.555 0.465 ;
        RECT  2.360 0.735 2.555 0.845 ;
        RECT  1.990 0.545 2.390 0.620 ;
        RECT  2.280 0.185 2.360 0.465 ;
        RECT  2.280 0.735 2.360 1.055 ;
        RECT  1.910 0.195 1.990 1.055 ;
        RECT  1.650 0.985 1.910 1.055 ;
        RECT  1.770 0.205 1.840 0.915 ;
        RECT  1.090 0.205 1.770 0.275 ;
        RECT  0.590 0.845 1.770 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCNDQD4BWP

MACRO LHCNQD1BWP
    CLASS CORE ;
    FOREIGN LHCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.345 1.045 ;
        RECT  2.250 0.185 2.275 0.465 ;
        RECT  2.250 0.705 2.275 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.040 -0.115 2.120 0.300 ;
        RECT  1.530 -0.115 2.040 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.040 0.880 2.120 1.375 ;
        RECT  1.520 1.145 2.040 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.540 2.205 0.620 ;
        RECT  2.050 0.380 2.120 0.800 ;
        RECT  1.910 0.380 2.050 0.465 ;
        RECT  1.910 0.720 2.050 0.800 ;
        RECT  1.715 0.545 1.980 0.620 ;
        RECT  1.830 0.185 1.910 0.465 ;
        RECT  1.830 0.720 1.910 1.040 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCNQD1BWP

MACRO LHCNQD2BWP
    CLASS CORE ;
    FOREIGN LHCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.355 2.345 0.765 ;
        RECT  2.275 0.185 2.290 1.050 ;
        RECT  2.210 0.185 2.275 0.465 ;
        RECT  2.210 0.695 2.275 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.290 ;
        RECT  2.100 -0.115 2.390 0.115 ;
        RECT  2.020 -0.115 2.100 0.300 ;
        RECT  1.530 -0.115 2.020 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.850 2.480 1.375 ;
        RECT  2.100 1.145 2.380 1.375 ;
        RECT  2.020 0.880 2.100 1.375 ;
        RECT  1.520 1.145 2.020 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.545 2.195 0.615 ;
        RECT  2.050 0.380 2.120 0.800 ;
        RECT  1.910 0.380 2.050 0.465 ;
        RECT  1.910 0.720 2.050 0.800 ;
        RECT  1.710 0.545 1.980 0.615 ;
        RECT  1.830 0.185 1.910 0.465 ;
        RECT  1.830 0.720 1.910 1.040 ;
        RECT  1.635 0.185 1.710 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.485 0.205 1.555 0.920 ;
        RECT  0.830 0.205 1.485 0.275 ;
        RECT  0.370 0.850 1.485 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCNQD2BWP

MACRO LHCNQD4BWP
    CLASS CORE ;
    FOREIGN LHCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.185 2.850 0.485 ;
        RECT  2.770 0.760 2.850 1.040 ;
        RECT  2.695 0.355 2.770 0.485 ;
        RECT  2.695 0.760 2.770 0.905 ;
        RECT  2.485 0.355 2.695 0.905 ;
        RECT  2.455 0.355 2.485 0.485 ;
        RECT  2.450 0.760 2.485 0.905 ;
        RECT  2.370 0.185 2.455 0.485 ;
        RECT  2.370 0.760 2.450 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.465 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.670 0.275 ;
        RECT  2.260 -0.115 2.570 0.115 ;
        RECT  2.180 -0.115 2.260 0.460 ;
        RECT  1.890 -0.115 2.180 0.115 ;
        RECT  1.810 -0.115 1.890 0.460 ;
        RECT  1.530 -0.115 1.810 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.685 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.570 0.985 2.670 1.375 ;
        RECT  2.260 1.145 2.570 1.375 ;
        RECT  2.180 0.750 2.260 1.375 ;
        RECT  1.890 1.145 2.180 1.375 ;
        RECT  1.810 0.750 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.770 0.185 2.850 0.485 ;
        RECT  2.770 0.760 2.850 1.040 ;
        RECT  2.765 0.355 2.770 0.485 ;
        RECT  2.765 0.760 2.770 0.905 ;
        RECT  2.370 0.185 2.415 0.485 ;
        RECT  2.370 0.760 2.415 1.040 ;
        RECT  2.070 0.560 2.380 0.630 ;
        RECT  1.990 0.185 2.070 1.060 ;
        RECT  1.710 0.540 1.910 0.620 ;
        RECT  1.630 0.185 1.710 1.060 ;
        RECT  1.370 0.990 1.630 1.060 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.125 0.990 0.850 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCNQD4BWP

MACRO LHCSND1BWP
    CLASS CORE ;
    FOREIGN LHCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.950 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.720 2.550 0.790 ;
        RECT  2.485 0.185 2.515 0.465 ;
        RECT  2.410 0.185 2.485 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.185 2.905 1.045 ;
        RECT  2.815 0.185 2.835 0.465 ;
        RECT  2.815 0.745 2.835 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.105 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.105 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 -0.115 2.940 0.115 ;
        RECT  2.620 -0.115 2.700 0.375 ;
        RECT  2.170 -0.115 2.620 0.115 ;
        RECT  2.050 -0.115 2.170 0.275 ;
        RECT  1.530 -0.115 2.050 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 2.940 1.375 ;
        RECT  2.600 1.020 2.720 1.375 ;
        RECT  2.110 1.145 2.600 1.375 ;
        RECT  2.010 0.990 2.110 1.375 ;
        RECT  1.520 1.145 2.010 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.705 0.520 2.765 0.640 ;
        RECT  2.635 0.520 2.705 0.940 ;
        RECT  2.330 0.870 2.635 0.940 ;
        RECT  2.250 0.185 2.330 1.045 ;
        RECT  2.090 0.345 2.170 0.910 ;
        RECT  1.810 0.345 2.090 0.415 ;
        RECT  1.890 0.840 2.090 0.910 ;
        RECT  1.810 0.840 1.890 1.060 ;
        RECT  1.370 0.990 1.810 1.060 ;
        RECT  1.505 0.205 1.585 0.920 ;
        RECT  0.830 0.205 1.505 0.275 ;
        RECT  0.370 0.850 1.505 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.840 0.990 1.000 1.075 ;
        RECT  0.125 0.990 0.840 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCSND1BWP

MACRO LHCSND2BWP
    CLASS CORE ;
    FOREIGN LHCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.805 0.495 1.855 0.640 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.400 0.185 2.485 0.820 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.060 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.740 2.835 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 -0.115 3.080 0.115 ;
        RECT  2.940 -0.115 3.040 0.290 ;
        RECT  2.660 -0.115 2.940 0.115 ;
        RECT  2.580 -0.115 2.660 0.465 ;
        RECT  2.300 -0.115 2.580 0.115 ;
        RECT  2.180 -0.115 2.300 0.135 ;
        RECT  1.530 -0.115 2.180 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.985 3.030 1.375 ;
        RECT  2.680 1.145 2.950 1.375 ;
        RECT  2.560 1.040 2.680 1.375 ;
        RECT  2.305 1.145 2.560 1.375 ;
        RECT  2.185 1.040 2.305 1.375 ;
        RECT  1.910 1.145 2.185 1.375 ;
        RECT  1.830 0.960 1.910 1.375 ;
        RECT  1.520 1.145 1.830 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.620 ;
        RECT  2.590 0.545 2.665 0.970 ;
        RECT  2.090 0.900 2.590 0.970 ;
        RECT  2.190 0.205 2.270 0.660 ;
        RECT  1.730 0.205 2.190 0.275 ;
        RECT  2.010 0.345 2.090 0.970 ;
        RECT  1.655 0.205 1.730 1.060 ;
        RECT  1.370 0.990 1.655 1.060 ;
        RECT  1.505 0.205 1.585 0.920 ;
        RECT  0.830 0.205 1.505 0.275 ;
        RECT  0.370 0.850 1.505 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.840 0.990 1.000 1.075 ;
        RECT  0.125 0.990 0.840 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCSND2BWP

MACRO LHCSND4BWP
    CLASS CORE ;
    FOREIGN LHCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.700 3.270 0.800 ;
        RECT  3.175 0.185 3.245 0.485 ;
        RECT  3.115 0.355 3.175 0.485 ;
        RECT  2.905 0.355 3.115 0.800 ;
        RECT  2.885 0.355 2.905 0.485 ;
        RECT  2.790 0.700 2.905 0.800 ;
        RECT  2.815 0.185 2.885 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.465 ;
        RECT  3.955 0.735 3.965 1.035 ;
        RECT  3.895 0.185 3.955 1.035 ;
        RECT  3.745 0.355 3.895 0.905 ;
        RECT  3.605 0.355 3.745 0.465 ;
        RECT  3.605 0.735 3.745 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.735 3.605 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.460 ;
        RECT  3.800 -0.115 4.070 0.115 ;
        RECT  3.700 -0.115 3.800 0.275 ;
        RECT  3.430 -0.115 3.700 0.115 ;
        RECT  3.350 -0.115 3.430 0.460 ;
        RECT  3.080 -0.115 3.350 0.115 ;
        RECT  2.980 -0.115 3.080 0.275 ;
        RECT  2.710 -0.115 2.980 0.115 ;
        RECT  2.630 -0.115 2.710 0.315 ;
        RECT  2.340 -0.115 2.630 0.115 ;
        RECT  2.220 -0.115 2.340 0.265 ;
        RECT  1.520 -0.115 2.220 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.665 4.150 1.375 ;
        RECT  3.800 1.145 4.070 1.375 ;
        RECT  3.700 0.985 3.800 1.375 ;
        RECT  3.450 1.145 3.700 1.375 ;
        RECT  3.330 1.010 3.450 1.375 ;
        RECT  3.090 1.145 3.330 1.375 ;
        RECT  2.970 1.010 3.090 1.375 ;
        RECT  2.730 1.145 2.970 1.375 ;
        RECT  2.610 1.010 2.730 1.375 ;
        RECT  2.340 1.145 2.610 1.375 ;
        RECT  2.220 1.000 2.340 1.375 ;
        RECT  1.920 1.145 2.220 1.375 ;
        RECT  1.800 1.000 1.920 1.375 ;
        RECT  1.520 1.145 1.800 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.355 3.675 0.465 ;
        RECT  3.605 0.735 3.675 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.735 3.605 1.035 ;
        RECT  3.185 0.700 3.270 0.800 ;
        RECT  3.185 0.185 3.245 0.485 ;
        RECT  2.815 0.185 2.835 0.485 ;
        RECT  2.790 0.700 2.835 0.800 ;
        RECT  3.420 0.540 3.650 0.620 ;
        RECT  3.350 0.540 3.420 0.940 ;
        RECT  2.720 0.870 3.350 0.940 ;
        RECT  2.650 0.395 2.720 0.940 ;
        RECT  2.100 0.500 2.180 0.780 ;
        RECT  1.600 0.710 2.100 0.780 ;
        RECT  1.800 0.205 1.920 0.415 ;
        RECT  1.630 0.850 1.710 1.060 ;
        RECT  1.370 0.990 1.630 1.060 ;
        RECT  1.550 0.520 1.600 0.780 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.840 0.990 1.000 1.075 ;
        RECT  0.125 0.990 0.840 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
        RECT  2.525 0.395 2.650 0.465 ;
        RECT  2.530 0.870 2.650 0.940 ;
        RECT  2.380 0.545 2.580 0.625 ;
        RECT  2.450 0.740 2.530 1.060 ;
        RECT  2.455 0.185 2.525 0.465 ;
        RECT  2.310 0.345 2.380 0.920 ;
        RECT  1.920 0.345 2.310 0.415 ;
        RECT  1.710 0.850 2.310 0.920 ;
    END
END LHCSND4BWP

MACRO LHCSNDD1BWP
    CLASS CORE ;
    FOREIGN LHCSNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.230 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.720 2.830 0.790 ;
        RECT  2.765 0.185 2.795 0.465 ;
        RECT  2.690 0.185 2.765 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.185 1.045 ;
        RECT  3.095 0.185 3.115 0.465 ;
        RECT  3.095 0.745 3.115 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.110 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.980 0.375 ;
        RECT  2.450 -0.115 2.900 0.115 ;
        RECT  2.330 -0.115 2.450 0.275 ;
        RECT  1.810 -0.115 2.330 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 1.145 3.220 1.375 ;
        RECT  2.880 1.020 3.000 1.375 ;
        RECT  2.390 1.145 2.880 1.375 ;
        RECT  2.290 0.990 2.390 1.375 ;
        RECT  1.800 1.145 2.290 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.985 0.520 3.045 0.640 ;
        RECT  2.915 0.520 2.985 0.940 ;
        RECT  2.610 0.870 2.915 0.940 ;
        RECT  2.530 0.185 2.610 1.045 ;
        RECT  2.370 0.345 2.450 0.910 ;
        RECT  2.090 0.345 2.370 0.415 ;
        RECT  2.170 0.840 2.370 0.910 ;
        RECT  2.090 0.840 2.170 1.060 ;
        RECT  1.650 0.985 2.090 1.060 ;
        RECT  1.790 0.210 1.870 0.915 ;
        RECT  1.110 0.210 1.790 0.280 ;
        RECT  0.590 0.845 1.790 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.440 0.260 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHCSNDD1BWP

MACRO LHCSNDD2BWP
    CLASS CORE ;
    FOREIGN LHCSNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.105 0.640 ;
        RECT  1.995 0.495 2.065 0.780 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.690 0.185 2.770 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 0.355 3.185 0.905 ;
        RECT  3.115 0.185 3.130 1.055 ;
        RECT  3.050 0.185 3.115 0.465 ;
        RECT  3.050 0.735 3.115 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.110 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.115 3.360 0.115 ;
        RECT  3.235 -0.115 3.305 0.305 ;
        RECT  2.950 -0.115 3.235 0.115 ;
        RECT  2.870 -0.115 2.950 0.465 ;
        RECT  2.590 -0.115 2.870 0.115 ;
        RECT  2.510 -0.115 2.590 0.305 ;
        RECT  1.810 -0.115 2.510 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.145 3.360 1.375 ;
        RECT  3.235 0.960 3.305 1.375 ;
        RECT  2.970 1.145 3.235 1.375 ;
        RECT  2.850 1.005 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.005 2.610 1.375 ;
        RECT  2.240 1.145 2.490 1.375 ;
        RECT  2.140 0.990 2.240 1.375 ;
        RECT  1.800 1.145 2.140 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.545 3.045 0.615 ;
        RECT  2.875 0.545 2.945 0.935 ;
        RECT  2.520 0.865 2.875 0.935 ;
        RECT  2.450 0.385 2.520 0.935 ;
        RECT  2.410 0.385 2.450 0.465 ;
        RECT  2.410 0.735 2.450 0.935 ;
        RECT  2.330 0.185 2.410 0.465 ;
        RECT  2.330 0.735 2.410 1.055 ;
        RECT  2.255 0.545 2.380 0.620 ;
        RECT  2.185 0.275 2.255 0.920 ;
        RECT  2.090 0.275 2.185 0.355 ;
        RECT  2.020 0.850 2.185 0.920 ;
        RECT  1.940 0.850 2.020 1.060 ;
        RECT  1.650 0.985 1.940 1.060 ;
        RECT  1.790 0.210 1.870 0.915 ;
        RECT  1.110 0.210 1.790 0.280 ;
        RECT  0.590 0.845 1.790 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.440 0.260 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHCSNDD2BWP

MACRO LHCSNDD4BWP
    CLASS CORE ;
    FOREIGN LHCSNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.705 3.410 0.795 ;
        RECT  3.315 0.185 3.385 0.485 ;
        RECT  3.255 0.355 3.315 0.485 ;
        RECT  3.045 0.355 3.255 0.795 ;
        RECT  3.025 0.355 3.045 0.485 ;
        RECT  2.930 0.705 3.045 0.795 ;
        RECT  2.955 0.185 3.025 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.105 0.465 ;
        RECT  4.095 0.775 4.105 1.055 ;
        RECT  4.035 0.185 4.095 1.055 ;
        RECT  3.885 0.355 4.035 0.905 ;
        RECT  3.745 0.355 3.885 0.465 ;
        RECT  3.745 0.775 3.885 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.775 3.745 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.485 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.570 -0.115 3.830 0.115 ;
        RECT  3.490 -0.115 3.570 0.465 ;
        RECT  3.230 -0.115 3.490 0.115 ;
        RECT  3.110 -0.115 3.230 0.275 ;
        RECT  2.850 -0.115 3.110 0.115 ;
        RECT  2.770 -0.115 2.850 0.305 ;
        RECT  2.500 -0.115 2.770 0.115 ;
        RECT  2.400 -0.115 2.500 0.275 ;
        RECT  1.780 -0.115 2.400 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.665 4.290 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 0.985 3.950 1.375 ;
        RECT  3.590 1.145 3.830 1.375 ;
        RECT  3.470 1.005 3.590 1.375 ;
        RECT  3.230 1.145 3.470 1.375 ;
        RECT  3.110 1.005 3.230 1.375 ;
        RECT  2.870 1.145 3.110 1.375 ;
        RECT  2.750 1.005 2.870 1.375 ;
        RECT  2.510 1.145 2.750 1.375 ;
        RECT  2.390 0.995 2.510 1.375 ;
        RECT  2.150 1.145 2.390 1.375 ;
        RECT  2.030 0.995 2.150 1.375 ;
        RECT  0.910 1.145 2.030 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.355 3.815 0.465 ;
        RECT  3.745 0.775 3.815 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.775 3.745 1.055 ;
        RECT  3.325 0.705 3.410 0.795 ;
        RECT  3.325 0.185 3.385 0.485 ;
        RECT  2.955 0.185 2.975 0.485 ;
        RECT  2.930 0.705 2.975 0.795 ;
        RECT  3.565 0.540 3.795 0.620 ;
        RECT  3.495 0.540 3.565 0.935 ;
        RECT  2.810 0.865 3.495 0.935 ;
        RECT  2.740 0.385 2.810 0.935 ;
        RECT  2.670 0.385 2.740 0.465 ;
        RECT  2.670 0.735 2.740 0.935 ;
        RECT  2.590 0.185 2.670 0.465 ;
        RECT  2.590 0.735 2.670 1.055 ;
        RECT  2.515 0.545 2.660 0.620 ;
        RECT  2.445 0.345 2.515 0.925 ;
        RECT  2.150 0.345 2.445 0.415 ;
        RECT  1.950 0.855 2.445 0.925 ;
        RECT  2.300 0.500 2.375 0.775 ;
        RECT  1.820 0.705 2.300 0.775 ;
        RECT  2.030 0.205 2.150 0.415 ;
        RECT  1.870 0.855 1.950 1.055 ;
        RECT  1.670 0.985 1.870 1.055 ;
        RECT  1.795 0.520 1.820 0.775 ;
        RECT  1.725 0.205 1.795 0.915 ;
        RECT  1.090 0.205 1.725 0.275 ;
        RECT  0.590 0.845 1.725 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCSNDD4BWP

MACRO LHCSNDQD1BWP
    CLASS CORE ;
    FOREIGN LHCSNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.495 2.065 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 0.355 2.765 0.905 ;
        RECT  2.695 0.185 2.730 1.055 ;
        RECT  2.650 0.185 2.695 0.465 ;
        RECT  2.650 0.735 2.695 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 -0.115 2.800 0.115 ;
        RECT  2.460 -0.115 2.540 0.315 ;
        RECT  1.780 -0.115 2.460 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 1.145 2.800 1.375 ;
        RECT  2.460 0.885 2.540 1.375 ;
        RECT  2.160 1.145 2.460 1.375 ;
        RECT  2.060 0.990 2.160 1.375 ;
        RECT  0.910 1.145 2.060 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.545 2.625 0.620 ;
        RECT  2.480 0.395 2.550 0.805 ;
        RECT  2.350 0.395 2.480 0.465 ;
        RECT  2.350 0.735 2.480 0.805 ;
        RECT  2.205 0.545 2.400 0.620 ;
        RECT  2.275 0.185 2.350 0.465 ;
        RECT  2.275 0.735 2.350 1.055 ;
        RECT  2.135 0.275 2.205 0.910 ;
        RECT  2.030 0.275 2.135 0.355 ;
        RECT  1.985 0.840 2.135 0.910 ;
        RECT  1.905 0.840 1.985 1.055 ;
        RECT  1.670 0.985 1.905 1.055 ;
        RECT  1.750 0.205 1.825 0.915 ;
        RECT  1.090 0.205 1.750 0.275 ;
        RECT  0.590 0.845 1.750 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.195 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCSNDQD1BWP

MACRO LHCSNDQD2BWP
    CLASS CORE ;
    FOREIGN LHCSNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.495 2.065 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.710 0.355 2.765 0.905 ;
        RECT  2.695 0.185 2.710 1.055 ;
        RECT  2.630 0.185 2.695 0.465 ;
        RECT  2.630 0.735 2.695 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.815 -0.115 2.890 0.305 ;
        RECT  2.530 -0.115 2.815 0.115 ;
        RECT  2.450 -0.115 2.530 0.315 ;
        RECT  1.780 -0.115 2.450 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.985 2.900 1.375 ;
        RECT  2.530 1.145 2.800 1.375 ;
        RECT  2.450 0.885 2.530 1.375 ;
        RECT  2.160 1.145 2.450 1.375 ;
        RECT  2.060 0.990 2.160 1.375 ;
        RECT  0.910 1.145 2.060 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.545 2.625 0.620 ;
        RECT  2.480 0.395 2.550 0.805 ;
        RECT  2.350 0.395 2.480 0.465 ;
        RECT  2.350 0.735 2.480 0.805 ;
        RECT  2.205 0.545 2.400 0.620 ;
        RECT  2.275 0.185 2.350 0.465 ;
        RECT  2.275 0.735 2.350 1.055 ;
        RECT  2.170 0.345 2.205 0.910 ;
        RECT  2.135 0.205 2.170 0.910 ;
        RECT  2.050 0.205 2.135 0.415 ;
        RECT  1.985 0.840 2.135 0.910 ;
        RECT  1.905 0.840 1.985 1.055 ;
        RECT  1.670 0.985 1.905 1.055 ;
        RECT  1.750 0.205 1.825 0.915 ;
        RECT  1.090 0.205 1.750 0.275 ;
        RECT  0.590 0.845 1.750 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.195 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCSNDQD2BWP

MACRO LHCSNDQD4BWP
    CLASS CORE ;
    FOREIGN LHCSNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.185 3.265 0.465 ;
        RECT  3.255 0.775 3.265 1.055 ;
        RECT  3.195 0.185 3.255 1.055 ;
        RECT  3.045 0.355 3.195 0.905 ;
        RECT  2.905 0.355 3.045 0.465 ;
        RECT  2.905 0.775 3.045 0.905 ;
        RECT  2.835 0.185 2.905 0.465 ;
        RECT  2.835 0.775 2.905 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.485 ;
        RECT  3.110 -0.115 3.370 0.115 ;
        RECT  2.990 -0.115 3.110 0.275 ;
        RECT  2.730 -0.115 2.990 0.115 ;
        RECT  2.650 -0.115 2.730 0.305 ;
        RECT  2.380 -0.115 2.650 0.115 ;
        RECT  2.280 -0.115 2.380 0.275 ;
        RECT  1.780 -0.115 2.280 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.665 3.450 1.375 ;
        RECT  3.110 1.145 3.370 1.375 ;
        RECT  2.990 0.985 3.110 1.375 ;
        RECT  2.730 1.145 2.990 1.375 ;
        RECT  2.650 0.925 2.730 1.375 ;
        RECT  2.370 1.145 2.650 1.375 ;
        RECT  2.290 0.925 2.370 1.375 ;
        RECT  2.190 1.145 2.290 1.375 ;
        RECT  2.110 0.925 2.190 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.355 2.975 0.465 ;
        RECT  2.905 0.775 2.975 0.905 ;
        RECT  2.835 0.185 2.905 0.465 ;
        RECT  2.835 0.775 2.905 1.055 ;
        RECT  2.750 0.545 2.850 0.615 ;
        RECT  2.680 0.385 2.750 0.805 ;
        RECT  2.550 0.385 2.680 0.465 ;
        RECT  2.550 0.735 2.680 0.805 ;
        RECT  2.345 0.545 2.590 0.620 ;
        RECT  2.470 0.185 2.550 0.465 ;
        RECT  2.470 0.735 2.550 1.055 ;
        RECT  2.275 0.345 2.345 0.845 ;
        RECT  2.070 0.345 2.275 0.415 ;
        RECT  2.000 0.775 2.275 0.845 ;
        RECT  1.920 0.775 2.000 1.055 ;
        RECT  1.650 0.985 1.920 1.055 ;
        RECT  1.820 0.540 1.900 0.620 ;
        RECT  1.740 0.205 1.820 0.915 ;
        RECT  1.090 0.205 1.740 0.275 ;
        RECT  0.590 0.845 1.740 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.370 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.130 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.050 0.860 0.130 1.055 ;
    END
END LHCSNDQD4BWP

MACRO LHCSNQD1BWP
    CLASS CORE ;
    FOREIGN LHCSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.450 1.060 ;
        RECT  2.370 0.185 2.415 0.465 ;
        RECT  2.370 0.740 2.415 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.705 1.230 0.775 ;
        RECT  0.870 0.495 0.945 0.775 ;
        RECT  0.780 0.495 0.870 0.565 ;
        RECT  0.250 0.705 0.870 0.775 ;
        RECT  0.175 0.495 0.250 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 0.490 0.680 0.560 ;
        RECT  0.455 0.355 0.530 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0244 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.395 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.770 0.345 1.015 0.415 ;
        RECT  0.700 0.205 0.770 0.415 ;
        RECT  0.480 0.205 0.700 0.275 ;
        RECT  0.340 0.190 0.480 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.180 -0.115 2.260 0.315 ;
        RECT  1.520 -0.115 2.180 0.115 ;
        RECT  1.400 -0.115 1.520 0.130 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.330 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.180 0.900 2.260 1.375 ;
        RECT  1.890 1.145 2.180 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  0.720 1.145 1.810 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.340 0.620 ;
        RECT  2.200 0.395 2.270 0.785 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.710 2.200 0.785 ;
        RECT  1.925 0.545 2.110 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.710 2.070 1.030 ;
        RECT  1.910 0.345 1.925 0.910 ;
        RECT  1.855 0.205 1.910 0.910 ;
        RECT  1.790 0.205 1.855 0.415 ;
        RECT  1.710 0.840 1.855 0.910 ;
        RECT  1.630 0.840 1.710 1.055 ;
        RECT  1.440 0.985 1.630 1.055 ;
        RECT  1.560 0.520 1.575 0.640 ;
        RECT  1.555 0.520 1.560 0.915 ;
        RECT  1.485 0.205 1.555 0.915 ;
        RECT  0.850 0.205 1.485 0.275 ;
        RECT  0.390 0.845 1.485 0.915 ;
        RECT  1.300 0.985 1.440 1.075 ;
        RECT  0.830 0.985 0.950 1.075 ;
        RECT  0.125 0.985 0.830 1.055 ;
        RECT  0.105 0.915 0.125 1.055 ;
        RECT  0.105 0.310 0.120 0.430 ;
        RECT  0.035 0.310 0.105 1.055 ;
    END
END LHCSNQD1BWP

MACRO LHCSNQD2BWP
    CLASS CORE ;
    FOREIGN LHCSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.060 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.740 2.415 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.705 1.230 0.775 ;
        RECT  0.870 0.495 0.945 0.775 ;
        RECT  0.780 0.495 0.870 0.565 ;
        RECT  0.250 0.705 0.870 0.775 ;
        RECT  0.175 0.495 0.250 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0180 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 0.490 0.680 0.560 ;
        RECT  0.455 0.355 0.530 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0244 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.395 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.770 0.345 1.015 0.415 ;
        RECT  0.700 0.205 0.770 0.415 ;
        RECT  0.480 0.205 0.700 0.275 ;
        RECT  0.340 0.190 0.480 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.290 ;
        RECT  2.250 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.520 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.520 0.130 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.330 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.145 2.660 1.375 ;
        RECT  2.520 0.985 2.620 1.375 ;
        RECT  2.250 1.145 2.520 1.375 ;
        RECT  2.170 0.900 2.250 1.375 ;
        RECT  1.890 1.145 2.170 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  0.720 1.145 1.810 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.340 0.620 ;
        RECT  2.200 0.395 2.270 0.785 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.710 2.200 0.785 ;
        RECT  1.925 0.545 2.110 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.710 2.070 1.030 ;
        RECT  1.855 0.300 1.925 0.910 ;
        RECT  1.770 0.300 1.855 0.380 ;
        RECT  1.710 0.840 1.855 0.910 ;
        RECT  1.630 0.840 1.710 1.055 ;
        RECT  1.440 0.985 1.630 1.055 ;
        RECT  1.560 0.520 1.575 0.640 ;
        RECT  1.555 0.520 1.560 0.915 ;
        RECT  1.485 0.205 1.555 0.915 ;
        RECT  0.850 0.205 1.485 0.275 ;
        RECT  0.390 0.845 1.485 0.915 ;
        RECT  1.280 0.985 1.440 1.075 ;
        RECT  0.830 0.985 0.950 1.075 ;
        RECT  0.125 0.985 0.830 1.055 ;
        RECT  0.105 0.915 0.125 1.055 ;
        RECT  0.105 0.310 0.120 0.430 ;
        RECT  0.035 0.310 0.105 1.055 ;
    END
END LHCSNQD2BWP

MACRO LHCSNQD4BWP
    CLASS CORE ;
    FOREIGN LHCSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.185 2.990 0.485 ;
        RECT  2.910 0.760 2.990 1.040 ;
        RECT  2.835 0.355 2.910 0.485 ;
        RECT  2.835 0.760 2.910 0.905 ;
        RECT  2.630 0.355 2.835 0.905 ;
        RECT  2.625 0.355 2.630 1.040 ;
        RECT  2.540 0.185 2.625 0.480 ;
        RECT  2.540 0.760 2.625 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0448 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.705 1.250 0.780 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.780 ;
        RECT  0.250 0.710 0.735 0.780 ;
        RECT  0.175 0.495 0.250 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.485 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.280 ;
        RECT  2.440 -0.115 2.710 0.115 ;
        RECT  2.360 -0.115 2.440 0.465 ;
        RECT  2.090 -0.115 2.360 0.115 ;
        RECT  1.970 -0.115 2.090 0.275 ;
        RECT  1.530 -0.115 1.970 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.665 3.170 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.005 2.830 1.375 ;
        RECT  2.440 1.145 2.710 1.375 ;
        RECT  2.360 0.740 2.440 1.375 ;
        RECT  2.070 1.145 2.360 1.375 ;
        RECT  1.990 0.980 2.070 1.375 ;
        RECT  1.890 1.145 1.990 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.910 0.185 2.990 0.485 ;
        RECT  2.910 0.760 2.990 1.040 ;
        RECT  2.905 0.355 2.910 0.485 ;
        RECT  2.905 0.760 2.910 0.905 ;
        RECT  2.540 0.185 2.555 0.480 ;
        RECT  2.540 0.760 2.555 1.040 ;
        RECT  2.250 0.550 2.530 0.620 ;
        RECT  2.170 0.185 2.250 1.070 ;
        RECT  2.010 0.355 2.090 0.910 ;
        RECT  1.770 0.355 2.010 0.425 ;
        RECT  1.730 0.840 2.010 0.910 ;
        RECT  1.660 0.840 1.730 1.060 ;
        RECT  1.370 0.990 1.660 1.060 ;
        RECT  1.505 0.205 1.585 0.920 ;
        RECT  0.830 0.205 1.505 0.275 ;
        RECT  0.370 0.850 1.505 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.840 0.990 1.000 1.075 ;
        RECT  0.125 0.990 0.840 1.060 ;
        RECT  0.105 0.880 0.125 1.060 ;
        RECT  0.105 0.290 0.120 0.430 ;
        RECT  0.035 0.290 0.105 1.060 ;
    END
END LHCSNQD4BWP

MACRO LHD1BWP
    CLASS CORE ;
    FOREIGN LHD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.185 2.205 1.045 ;
        RECT  2.110 0.185 2.135 0.465 ;
        RECT  2.110 0.725 2.135 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.350 1.805 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.670 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 -0.115 2.240 0.115 ;
        RECT  1.900 -0.115 2.020 0.140 ;
        RECT  1.440 -0.115 1.900 0.115 ;
        RECT  1.360 -0.115 1.440 0.300 ;
        RECT  0.690 -0.115 1.360 0.115 ;
        RECT  0.570 -0.115 0.690 0.275 ;
        RECT  0.360 -0.115 0.570 0.115 ;
        RECT  0.240 -0.115 0.360 0.150 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 1.145 2.240 1.375 ;
        RECT  1.900 1.120 2.020 1.375 ;
        RECT  1.470 1.145 1.900 1.375 ;
        RECT  1.350 0.860 1.470 1.375 ;
        RECT  0.680 1.145 1.350 1.375 ;
        RECT  0.580 0.845 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.990 0.520 2.060 0.640 ;
        RECT  1.920 0.210 1.990 1.050 ;
        RECT  1.630 0.210 1.920 0.280 ;
        RECT  1.630 0.980 1.920 1.050 ;
        RECT  1.550 0.210 1.630 0.465 ;
        RECT  1.480 0.545 1.630 0.620 ;
        RECT  1.550 0.730 1.630 1.050 ;
        RECT  1.310 0.395 1.550 0.465 ;
        RECT  1.410 0.545 1.480 0.790 ;
        RECT  1.140 0.720 1.410 0.790 ;
        RECT  1.240 0.395 1.310 0.640 ;
        RECT  1.020 0.985 1.180 1.075 ;
        RECT  1.070 0.195 1.140 0.905 ;
        RECT  0.930 0.195 1.070 0.275 ;
        RECT  0.930 0.835 1.070 0.905 ;
        RECT  0.830 0.985 1.020 1.055 ;
        RECT  0.830 0.395 1.000 0.465 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.440 0.345 0.510 1.060 ;
        RECT  0.400 0.345 0.440 0.445 ;
        RECT  0.410 0.900 0.440 1.060 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.260 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.130 0.850 0.260 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHD1BWP

MACRO LHD2BWP
    CLASS CORE ;
    FOREIGN LHD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.355 2.345 0.905 ;
        RECT  2.275 0.185 2.290 1.030 ;
        RECT  2.210 0.185 2.275 0.465 ;
        RECT  2.210 0.730 2.275 1.030 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.195 1.925 0.780 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.670 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.295 ;
        RECT  2.110 -0.115 2.390 0.115 ;
        RECT  2.030 -0.115 2.110 0.460 ;
        RECT  1.750 -0.115 2.030 0.115 ;
        RECT  1.670 -0.115 1.750 0.315 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.315 ;
        RECT  0.670 -0.115 1.310 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.360 -0.115 0.590 0.115 ;
        RECT  0.240 -0.115 0.360 0.150 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.485 1.145 2.520 1.375 ;
        RECT  2.375 0.980 2.485 1.375 ;
        RECT  2.120 1.145 2.375 1.375 ;
        RECT  2.020 0.990 2.120 1.375 ;
        RECT  1.760 1.145 2.020 1.375 ;
        RECT  1.660 0.990 1.760 1.375 ;
        RECT  1.405 1.145 1.660 1.375 ;
        RECT  1.300 0.860 1.405 1.375 ;
        RECT  0.680 1.145 1.300 1.375 ;
        RECT  0.580 0.845 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.090 0.545 2.200 0.620 ;
        RECT  2.020 0.545 2.090 0.920 ;
        RECT  1.730 0.850 2.020 0.920 ;
        RECT  1.660 0.395 1.730 0.920 ;
        RECT  1.570 0.395 1.660 0.465 ;
        RECT  1.570 0.850 1.660 0.920 ;
        RECT  1.420 0.545 1.580 0.615 ;
        RECT  1.490 0.185 1.570 0.465 ;
        RECT  1.490 0.720 1.570 1.040 ;
        RECT  1.280 0.395 1.490 0.465 ;
        RECT  1.350 0.545 1.420 0.790 ;
        RECT  1.120 0.720 1.350 0.790 ;
        RECT  1.200 0.395 1.280 0.640 ;
        RECT  1.000 0.985 1.160 1.075 ;
        RECT  1.050 0.195 1.120 0.915 ;
        RECT  0.910 0.195 1.050 0.275 ;
        RECT  0.910 0.840 1.050 0.915 ;
        RECT  0.830 0.985 1.000 1.055 ;
        RECT  0.830 0.390 0.970 0.470 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.440 0.345 0.510 1.060 ;
        RECT  0.400 0.345 0.440 0.445 ;
        RECT  0.410 0.900 0.440 1.060 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.260 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.130 0.850 0.260 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHD2BWP

MACRO LHD4BWP
    CLASS CORE ;
    FOREIGN LHD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.775 3.125 1.055 ;
        RECT  3.055 0.185 3.115 1.055 ;
        RECT  2.905 0.355 3.055 0.905 ;
        RECT  2.765 0.355 2.905 0.465 ;
        RECT  2.765 0.775 2.905 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.705 2.430 0.795 ;
        RECT  2.335 0.185 2.405 0.485 ;
        RECT  2.275 0.355 2.335 0.485 ;
        RECT  2.065 0.355 2.275 0.795 ;
        RECT  2.045 0.355 2.065 0.485 ;
        RECT  1.950 0.705 2.065 0.795 ;
        RECT  1.975 0.185 2.045 0.485 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.680 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.485 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.275 ;
        RECT  2.590 -0.115 2.850 0.115 ;
        RECT  2.510 -0.115 2.590 0.465 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.275 ;
        RECT  1.865 -0.115 2.130 0.115 ;
        RECT  1.795 -0.115 1.865 0.310 ;
        RECT  1.460 -0.115 1.795 0.115 ;
        RECT  1.380 -0.115 1.460 0.300 ;
        RECT  0.680 -0.115 1.380 0.115 ;
        RECT  0.580 -0.115 0.680 0.265 ;
        RECT  0.330 -0.115 0.580 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.665 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.985 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.005 2.610 1.375 ;
        RECT  2.250 1.145 2.490 1.375 ;
        RECT  2.130 1.005 2.250 1.375 ;
        RECT  1.890 1.145 2.130 1.375 ;
        RECT  1.770 1.005 1.890 1.375 ;
        RECT  1.470 1.145 1.770 1.375 ;
        RECT  1.370 0.850 1.470 1.375 ;
        RECT  0.680 1.145 1.370 1.375 ;
        RECT  0.580 0.850 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.465 ;
        RECT  2.765 0.775 2.835 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        RECT  2.345 0.705 2.430 0.795 ;
        RECT  2.345 0.185 2.405 0.485 ;
        RECT  1.975 0.185 1.995 0.485 ;
        RECT  1.950 0.705 1.995 0.795 ;
        RECT  2.585 0.540 2.815 0.620 ;
        RECT  2.515 0.540 2.585 0.935 ;
        RECT  1.860 0.865 2.515 0.935 ;
        RECT  1.790 0.395 1.860 0.935 ;
        RECT  1.650 0.395 1.790 0.465 ;
        RECT  1.650 0.865 1.790 0.935 ;
        RECT  1.490 0.545 1.710 0.620 ;
        RECT  1.570 0.185 1.650 0.465 ;
        RECT  1.570 0.720 1.650 1.040 ;
        RECT  1.340 0.395 1.570 0.465 ;
        RECT  1.420 0.545 1.490 0.780 ;
        RECT  1.120 0.710 1.420 0.780 ;
        RECT  1.260 0.395 1.340 0.640 ;
        RECT  1.010 0.985 1.170 1.075 ;
        RECT  1.050 0.195 1.120 0.910 ;
        RECT  0.910 0.195 1.050 0.265 ;
        RECT  0.910 0.840 1.050 0.910 ;
        RECT  0.830 0.985 1.010 1.055 ;
        RECT  0.830 0.390 0.970 0.470 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.490 0.345 0.510 0.790 ;
        RECT  0.440 0.185 0.490 1.040 ;
        RECT  0.415 0.185 0.440 0.465 ;
        RECT  0.410 0.720 0.440 1.040 ;
        RECT  0.340 0.520 0.370 0.640 ;
        RECT  0.270 0.320 0.340 0.920 ;
        RECT  0.130 0.320 0.270 0.390 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.230 0.130 0.390 ;
        RECT  0.050 0.850 0.130 1.020 ;
    END
END LHD4BWP

MACRO LHQD1BWP
    CLASS CORE ;
    FOREIGN LHQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.185 2.065 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0210 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.670 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 -0.115 2.100 0.115 ;
        RECT  1.790 -0.115 1.870 0.485 ;
        RECT  1.460 -0.115 1.790 0.115 ;
        RECT  1.380 -0.115 1.460 0.310 ;
        RECT  0.690 -0.115 1.380 0.115 ;
        RECT  0.570 -0.115 0.690 0.275 ;
        RECT  0.360 -0.115 0.570 0.115 ;
        RECT  0.240 -0.115 0.360 0.150 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.145 2.100 1.375 ;
        RECT  1.790 0.685 1.870 1.375 ;
        RECT  1.480 1.145 1.790 1.375 ;
        RECT  1.360 0.860 1.480 1.375 ;
        RECT  0.680 1.145 1.360 1.375 ;
        RECT  0.580 0.845 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.595 0.190 1.670 0.975 ;
        RECT  1.590 0.190 1.595 0.460 ;
        RECT  1.320 0.390 1.590 0.460 ;
        RECT  1.425 0.530 1.525 0.790 ;
        RECT  1.140 0.720 1.425 0.790 ;
        RECT  1.240 0.390 1.320 0.640 ;
        RECT  1.020 0.985 1.180 1.075 ;
        RECT  1.070 0.210 1.140 0.905 ;
        RECT  0.930 0.210 1.070 0.290 ;
        RECT  0.930 0.835 1.070 0.905 ;
        RECT  0.830 0.985 1.020 1.055 ;
        RECT  0.830 0.395 1.000 0.465 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.440 0.345 0.510 1.060 ;
        RECT  0.400 0.345 0.440 0.445 ;
        RECT  0.410 0.900 0.440 1.060 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.260 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.130 0.850 0.260 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD1BWP

MACRO LHQD2BWP
    CLASS CORE ;
    FOREIGN LHQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.195 1.925 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.670 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.115 2.240 0.115 ;
        RECT  2.050 -0.115 2.140 0.460 ;
        RECT  1.750 -0.115 2.050 0.115 ;
        RECT  1.670 -0.115 1.750 0.315 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.315 ;
        RECT  0.670 -0.115 1.310 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.360 -0.115 0.590 0.115 ;
        RECT  0.240 -0.115 0.360 0.150 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.145 2.240 1.375 ;
        RECT  2.050 0.665 2.140 1.375 ;
        RECT  1.400 1.145 2.050 1.375 ;
        RECT  1.300 0.860 1.400 1.375 ;
        RECT  0.680 1.145 1.300 1.375 ;
        RECT  0.580 0.845 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.660 0.395 1.730 0.935 ;
        RECT  1.570 0.395 1.660 0.465 ;
        RECT  1.470 0.865 1.660 0.935 ;
        RECT  1.420 0.545 1.580 0.615 ;
        RECT  1.490 0.185 1.570 0.465 ;
        RECT  1.280 0.395 1.490 0.465 ;
        RECT  1.350 0.545 1.420 0.790 ;
        RECT  1.120 0.720 1.350 0.790 ;
        RECT  1.200 0.395 1.280 0.640 ;
        RECT  1.000 0.985 1.160 1.075 ;
        RECT  1.050 0.195 1.120 0.915 ;
        RECT  0.910 0.195 1.050 0.275 ;
        RECT  0.910 0.840 1.050 0.915 ;
        RECT  0.830 0.985 1.000 1.055 ;
        RECT  0.830 0.390 0.980 0.470 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.440 0.345 0.510 1.060 ;
        RECT  0.400 0.345 0.440 0.445 ;
        RECT  0.410 0.900 0.440 1.060 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.260 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.130 0.850 0.260 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD2BWP

MACRO LHQD4BWP
    CLASS CORE ;
    FOREIGN LHQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.185 2.290 0.485 ;
        RECT  2.210 0.760 2.290 1.040 ;
        RECT  2.135 0.355 2.210 0.485 ;
        RECT  2.135 0.760 2.210 0.905 ;
        RECT  1.930 0.355 2.135 0.905 ;
        RECT  1.925 0.185 1.930 1.045 ;
        RECT  1.855 0.185 1.925 0.485 ;
        RECT  1.855 0.760 1.925 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0212 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.670 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.485 ;
        RECT  2.120 -0.115 2.390 0.115 ;
        RECT  2.020 -0.115 2.120 0.275 ;
        RECT  1.750 -0.115 2.020 0.115 ;
        RECT  1.675 -0.115 1.750 0.485 ;
        RECT  1.390 -0.115 1.675 0.115 ;
        RECT  1.310 -0.115 1.390 0.315 ;
        RECT  0.670 -0.115 1.310 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.330 -0.115 0.590 0.115 ;
        RECT  0.210 -0.115 0.330 0.265 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.665 2.470 1.375 ;
        RECT  2.120 1.145 2.390 1.375 ;
        RECT  2.020 0.985 2.120 1.375 ;
        RECT  1.750 1.145 2.020 1.375 ;
        RECT  1.675 0.685 1.750 1.375 ;
        RECT  1.400 1.145 1.675 1.375 ;
        RECT  1.300 0.860 1.400 1.375 ;
        RECT  0.680 1.145 1.300 1.375 ;
        RECT  0.580 0.845 0.680 1.375 ;
        RECT  0.330 1.145 0.580 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.210 0.185 2.290 0.485 ;
        RECT  2.210 0.760 2.290 1.040 ;
        RECT  2.205 0.355 2.210 0.485 ;
        RECT  2.205 0.760 2.210 0.905 ;
        RECT  1.570 0.395 1.605 0.940 ;
        RECT  1.535 0.185 1.570 0.940 ;
        RECT  1.490 0.185 1.535 0.465 ;
        RECT  1.470 0.860 1.535 0.940 ;
        RECT  1.280 0.395 1.490 0.465 ;
        RECT  1.380 0.545 1.460 0.770 ;
        RECT  1.120 0.700 1.380 0.770 ;
        RECT  1.200 0.395 1.280 0.620 ;
        RECT  1.000 0.985 1.160 1.075 ;
        RECT  1.050 0.195 1.120 0.915 ;
        RECT  0.910 0.195 1.050 0.275 ;
        RECT  0.910 0.840 1.050 0.915 ;
        RECT  0.830 0.985 1.000 1.055 ;
        RECT  0.830 0.390 0.980 0.470 ;
        RECT  0.760 0.345 0.830 1.055 ;
        RECT  0.510 0.345 0.760 0.415 ;
        RECT  0.500 0.345 0.510 1.060 ;
        RECT  0.440 0.185 0.500 1.060 ;
        RECT  0.400 0.185 0.440 0.445 ;
        RECT  0.410 0.740 0.440 1.060 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.345 0.330 0.920 ;
        RECT  0.130 0.345 0.260 0.415 ;
        RECT  0.130 0.850 0.260 0.920 ;
        RECT  0.050 0.255 0.130 0.415 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD4BWP

MACRO LHSND1BWP
    CLASS CORE ;
    FOREIGN LHSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.390 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.720 1.990 0.790 ;
        RECT  1.925 0.185 1.955 0.465 ;
        RECT  1.850 0.185 1.925 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.345 1.045 ;
        RECT  2.255 0.185 2.275 0.465 ;
        RECT  2.255 0.745 2.275 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0252 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.115 2.380 0.115 ;
        RECT  2.060 -0.115 2.140 0.375 ;
        RECT  1.610 -0.115 2.060 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  1.050 -0.115 1.490 0.115 ;
        RECT  0.970 -0.115 1.050 0.440 ;
        RECT  0.340 -0.115 0.970 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.145 2.380 1.375 ;
        RECT  2.040 1.020 2.160 1.375 ;
        RECT  1.550 1.145 2.040 1.375 ;
        RECT  1.450 0.990 1.550 1.375 ;
        RECT  0.350 1.145 1.450 1.375 ;
        RECT  0.230 1.130 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.145 0.520 2.205 0.640 ;
        RECT  2.075 0.520 2.145 0.940 ;
        RECT  1.770 0.870 2.075 0.940 ;
        RECT  1.690 0.185 1.770 1.045 ;
        RECT  1.530 0.345 1.610 0.910 ;
        RECT  1.290 0.345 1.530 0.415 ;
        RECT  1.310 0.840 1.530 0.910 ;
        RECT  1.230 0.840 1.310 1.055 ;
        RECT  0.840 0.985 1.230 1.055 ;
        RECT  1.080 0.515 1.160 0.640 ;
        RECT  0.975 0.515 1.080 0.585 ;
        RECT  0.905 0.515 0.975 0.915 ;
        RECT  0.865 0.515 0.905 0.585 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.585 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.120 0.960 0.450 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.105 0.890 0.120 1.030 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSND1BWP

MACRO LHSND2BWP
    CLASS CORE ;
    FOREIGN LHSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.365 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.065 0.800 ;
        RECT  1.960 0.185 1.995 0.465 ;
        RECT  1.925 0.730 1.995 0.800 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.050 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.730 2.415 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0252 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.290 ;
        RECT  2.240 -0.115 2.520 0.115 ;
        RECT  2.160 -0.115 2.240 0.465 ;
        RECT  1.845 -0.115 2.160 0.115 ;
        RECT  1.770 -0.115 1.845 0.465 ;
        RECT  1.050 -0.115 1.770 0.115 ;
        RECT  0.970 -0.115 1.050 0.440 ;
        RECT  0.340 -0.115 0.970 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.145 2.660 1.375 ;
        RECT  2.520 0.985 2.620 1.375 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.140 1.025 2.260 1.375 ;
        RECT  1.870 1.145 2.140 1.375 ;
        RECT  1.750 1.020 1.870 1.375 ;
        RECT  1.500 1.145 1.750 1.375 ;
        RECT  1.380 1.000 1.500 1.375 ;
        RECT  0.340 1.145 1.380 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.265 0.545 2.345 0.620 ;
        RECT  2.185 0.545 2.265 0.940 ;
        RECT  1.700 0.870 2.185 0.940 ;
        RECT  1.670 0.205 1.700 0.940 ;
        RECT  1.630 0.205 1.670 1.020 ;
        RECT  1.530 0.205 1.630 0.275 ;
        RECT  1.590 0.700 1.630 1.020 ;
        RECT  1.520 0.520 1.550 0.640 ;
        RECT  1.450 0.345 1.520 0.915 ;
        RECT  1.350 0.345 1.450 0.415 ;
        RECT  1.290 0.845 1.450 0.915 ;
        RECT  1.210 0.845 1.290 1.055 ;
        RECT  0.840 0.985 1.210 1.055 ;
        RECT  0.975 0.545 1.200 0.615 ;
        RECT  0.905 0.545 0.975 0.915 ;
        RECT  0.865 0.545 0.905 0.615 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.615 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.130 0.960 0.450 1.030 ;
        RECT  0.105 0.890 0.130 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSND2BWP

MACRO LHSND4BWP
    CLASS CORE ;
    FOREIGN LHSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.705 2.710 0.795 ;
        RECT  2.615 0.185 2.685 0.485 ;
        RECT  2.555 0.355 2.615 0.485 ;
        RECT  2.345 0.355 2.555 0.795 ;
        RECT  2.325 0.355 2.345 0.485 ;
        RECT  2.230 0.705 2.345 0.795 ;
        RECT  2.255 0.185 2.325 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.185 3.405 0.465 ;
        RECT  3.395 0.775 3.405 1.055 ;
        RECT  3.335 0.185 3.395 1.055 ;
        RECT  3.185 0.355 3.335 0.905 ;
        RECT  3.045 0.355 3.185 0.465 ;
        RECT  3.045 0.775 3.185 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0396 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.640 0.115 ;
        RECT  3.510 -0.115 3.590 0.485 ;
        RECT  3.250 -0.115 3.510 0.115 ;
        RECT  3.130 -0.115 3.250 0.275 ;
        RECT  2.870 -0.115 3.130 0.115 ;
        RECT  2.790 -0.115 2.870 0.465 ;
        RECT  2.530 -0.115 2.790 0.115 ;
        RECT  2.410 -0.115 2.530 0.275 ;
        RECT  2.150 -0.115 2.410 0.115 ;
        RECT  2.070 -0.115 2.150 0.315 ;
        RECT  1.810 -0.115 2.070 0.115 ;
        RECT  1.690 -0.115 1.810 0.265 ;
        RECT  1.070 -0.115 1.690 0.115 ;
        RECT  0.990 -0.115 1.070 0.320 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.665 3.590 1.375 ;
        RECT  3.250 1.145 3.510 1.375 ;
        RECT  3.130 0.985 3.250 1.375 ;
        RECT  2.890 1.145 3.130 1.375 ;
        RECT  2.770 1.005 2.890 1.375 ;
        RECT  2.530 1.145 2.770 1.375 ;
        RECT  2.410 1.005 2.530 1.375 ;
        RECT  2.170 1.145 2.410 1.375 ;
        RECT  2.050 1.005 2.170 1.375 ;
        RECT  1.810 1.145 2.050 1.375 ;
        RECT  1.690 1.010 1.810 1.375 ;
        RECT  1.450 1.145 1.690 1.375 ;
        RECT  1.330 1.010 1.450 1.375 ;
        RECT  0.340 1.145 1.330 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.355 3.115 0.465 ;
        RECT  3.045 0.775 3.115 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        RECT  2.625 0.705 2.710 0.795 ;
        RECT  2.625 0.185 2.685 0.485 ;
        RECT  2.255 0.185 2.275 0.485 ;
        RECT  2.230 0.705 2.275 0.795 ;
        RECT  2.865 0.540 3.095 0.620 ;
        RECT  2.795 0.540 2.865 0.935 ;
        RECT  2.160 0.865 2.795 0.935 ;
        RECT  2.090 0.395 2.160 0.935 ;
        RECT  1.970 0.395 2.090 0.465 ;
        RECT  1.970 0.865 2.090 0.935 ;
        RECT  1.820 0.545 2.010 0.620 ;
        RECT  1.890 0.185 1.970 0.465 ;
        RECT  1.890 0.740 1.970 1.060 ;
        RECT  1.750 0.345 1.820 0.940 ;
        RECT  1.450 0.345 1.750 0.415 ;
        RECT  1.250 0.870 1.750 0.940 ;
        RECT  1.600 0.500 1.680 0.800 ;
        RECT  1.180 0.730 1.600 0.800 ;
        RECT  1.330 0.205 1.450 0.415 ;
        RECT  1.170 0.870 1.250 1.055 ;
        RECT  1.100 0.500 1.180 0.800 ;
        RECT  0.830 0.985 1.170 1.055 ;
        RECT  0.975 0.500 1.100 0.570 ;
        RECT  0.905 0.500 0.975 0.915 ;
        RECT  0.865 0.500 0.905 0.570 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.570 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.130 0.960 0.450 1.030 ;
        RECT  0.105 0.890 0.130 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSND4BWP

MACRO LHSNDD1BWP
    CLASS CORE ;
    FOREIGN LHSNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.720 2.410 0.790 ;
        RECT  2.345 0.185 2.375 0.465 ;
        RECT  2.270 0.185 2.345 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.765 1.045 ;
        RECT  2.675 0.185 2.695 0.465 ;
        RECT  2.675 0.745 2.695 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 -0.115 2.800 0.115 ;
        RECT  2.480 -0.115 2.560 0.375 ;
        RECT  2.030 -0.115 2.480 0.115 ;
        RECT  1.910 -0.115 2.030 0.275 ;
        RECT  1.480 -0.115 1.910 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  0.700 -0.115 1.360 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.145 2.800 1.375 ;
        RECT  2.460 1.020 2.580 1.375 ;
        RECT  1.970 1.145 2.460 1.375 ;
        RECT  1.870 0.990 1.970 1.375 ;
        RECT  0.730 1.145 1.870 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.565 0.520 2.625 0.640 ;
        RECT  2.495 0.520 2.565 0.940 ;
        RECT  2.190 0.870 2.495 0.940 ;
        RECT  2.110 0.185 2.190 1.045 ;
        RECT  1.950 0.345 2.030 0.910 ;
        RECT  1.710 0.345 1.950 0.415 ;
        RECT  1.730 0.840 1.950 0.910 ;
        RECT  1.650 0.840 1.730 1.055 ;
        RECT  1.420 0.985 1.650 1.055 ;
        RECT  1.500 0.205 1.580 0.915 ;
        RECT  0.960 0.205 1.500 0.275 ;
        RECT  0.960 0.845 1.500 0.915 ;
        RECT  1.280 0.985 1.420 1.075 ;
        RECT  1.020 0.700 1.260 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.850 0.985 0.970 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.370 0.985 0.850 1.055 ;
        RECT  0.440 0.240 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.125 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.055 0.260 0.125 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDD1BWP

MACRO LHSNDD2BWP
    CLASS CORE ;
    FOREIGN LHSNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 1.835 0.640 ;
        RECT  1.715 0.495 1.785 0.780 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.055 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.735 2.835 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.115 3.080 0.115 ;
        RECT  2.955 -0.115 3.025 0.305 ;
        RECT  2.670 -0.115 2.955 0.115 ;
        RECT  2.590 -0.115 2.670 0.465 ;
        RECT  2.310 -0.115 2.590 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.520 -0.115 2.230 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.145 3.080 1.375 ;
        RECT  2.940 0.985 3.040 1.375 ;
        RECT  2.690 1.145 2.940 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  1.960 1.145 2.210 1.375 ;
        RECT  1.860 0.990 1.960 1.375 ;
        RECT  0.730 1.145 1.860 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.620 ;
        RECT  2.595 0.545 2.665 0.935 ;
        RECT  2.335 0.865 2.595 0.935 ;
        RECT  2.265 0.385 2.335 0.935 ;
        RECT  2.130 0.385 2.265 0.465 ;
        RECT  2.130 0.865 2.265 0.935 ;
        RECT  1.975 0.545 2.185 0.620 ;
        RECT  2.055 0.185 2.130 0.465 ;
        RECT  2.050 0.735 2.130 1.055 ;
        RECT  1.905 0.205 1.975 0.920 ;
        RECT  1.850 0.205 1.905 0.415 ;
        RECT  1.760 0.850 1.905 0.920 ;
        RECT  1.680 0.850 1.760 1.055 ;
        RECT  1.420 0.985 1.680 1.055 ;
        RECT  1.520 0.205 1.600 0.915 ;
        RECT  0.960 0.205 1.520 0.275 ;
        RECT  0.930 0.845 1.520 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.370 0.985 0.820 1.055 ;
        RECT  0.440 0.240 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDD2BWP

MACRO LHSNDD4BWP
    CLASS CORE ;
    FOREIGN LHSNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.705 3.130 0.795 ;
        RECT  3.035 0.185 3.105 0.485 ;
        RECT  2.975 0.355 3.035 0.485 ;
        RECT  2.765 0.355 2.975 0.795 ;
        RECT  2.745 0.355 2.765 0.485 ;
        RECT  2.650 0.705 2.765 0.795 ;
        RECT  2.675 0.185 2.745 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.825 0.465 ;
        RECT  3.815 0.775 3.825 1.055 ;
        RECT  3.755 0.185 3.815 1.055 ;
        RECT  3.605 0.355 3.755 0.905 ;
        RECT  3.465 0.355 3.605 0.465 ;
        RECT  3.465 0.775 3.605 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.485 ;
        RECT  3.670 -0.115 3.930 0.115 ;
        RECT  3.550 -0.115 3.670 0.275 ;
        RECT  3.290 -0.115 3.550 0.115 ;
        RECT  3.210 -0.115 3.290 0.465 ;
        RECT  2.950 -0.115 3.210 0.115 ;
        RECT  2.830 -0.115 2.950 0.275 ;
        RECT  2.570 -0.115 2.830 0.115 ;
        RECT  2.490 -0.115 2.570 0.305 ;
        RECT  2.220 -0.115 2.490 0.115 ;
        RECT  2.120 -0.115 2.220 0.275 ;
        RECT  1.480 -0.115 2.120 0.115 ;
        RECT  1.400 -0.115 1.480 0.420 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.665 4.010 1.375 ;
        RECT  3.670 1.145 3.930 1.375 ;
        RECT  3.550 0.985 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 1.005 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 1.005 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 1.005 2.590 1.375 ;
        RECT  2.230 1.145 2.470 1.375 ;
        RECT  2.110 0.995 2.230 1.375 ;
        RECT  1.870 1.145 2.110 1.375 ;
        RECT  1.750 0.995 1.870 1.375 ;
        RECT  0.730 1.145 1.750 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.355 3.535 0.465 ;
        RECT  3.465 0.775 3.535 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        RECT  3.045 0.705 3.130 0.795 ;
        RECT  3.045 0.185 3.105 0.485 ;
        RECT  2.675 0.185 2.695 0.485 ;
        RECT  2.650 0.705 2.695 0.795 ;
        RECT  3.285 0.540 3.515 0.620 ;
        RECT  3.215 0.540 3.285 0.935 ;
        RECT  2.570 0.865 3.215 0.935 ;
        RECT  2.500 0.385 2.570 0.935 ;
        RECT  2.390 0.385 2.500 0.465 ;
        RECT  2.390 0.865 2.500 0.935 ;
        RECT  2.240 0.545 2.420 0.620 ;
        RECT  2.310 0.185 2.390 0.465 ;
        RECT  2.310 0.735 2.390 1.055 ;
        RECT  2.170 0.345 2.240 0.925 ;
        RECT  1.870 0.345 2.170 0.415 ;
        RECT  1.670 0.855 2.170 0.925 ;
        RECT  2.020 0.500 2.100 0.775 ;
        RECT  1.600 0.705 2.020 0.775 ;
        RECT  1.750 0.205 1.870 0.415 ;
        RECT  1.590 0.855 1.670 1.055 ;
        RECT  1.520 0.540 1.600 0.775 ;
        RECT  1.410 0.985 1.590 1.055 ;
        RECT  1.380 0.540 1.520 0.620 ;
        RECT  1.260 0.985 1.410 1.075 ;
        RECT  1.310 0.540 1.380 0.915 ;
        RECT  1.270 0.540 1.310 0.620 ;
        RECT  0.930 0.845 1.310 0.915 ;
        RECT  1.200 0.205 1.270 0.620 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.960 0.205 1.200 0.275 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.370 0.985 0.820 1.055 ;
        RECT  0.440 0.190 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDD4BWP

MACRO LHSNDQD1BWP
    CLASS CORE ;
    FOREIGN LHSNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.450 1.055 ;
        RECT  2.370 0.185 2.415 0.465 ;
        RECT  2.370 0.735 2.415 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.520 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.145 2.520 1.375 ;
        RECT  2.170 0.885 2.250 1.375 ;
        RECT  1.900 1.145 2.170 1.375 ;
        RECT  1.800 0.990 1.900 1.375 ;
        RECT  0.730 1.145 1.800 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.345 0.620 ;
        RECT  2.200 0.395 2.270 0.805 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.735 2.200 0.805 ;
        RECT  1.925 0.545 2.120 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.735 2.070 1.055 ;
        RECT  1.855 0.275 1.925 0.915 ;
        RECT  1.770 0.275 1.855 0.355 ;
        RECT  1.710 0.845 1.855 0.915 ;
        RECT  1.630 0.845 1.710 1.055 ;
        RECT  1.420 0.985 1.630 1.055 ;
        RECT  1.425 0.540 1.620 0.620 ;
        RECT  1.345 0.205 1.425 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  0.960 0.205 1.345 0.275 ;
        RECT  0.930 0.845 1.345 0.915 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.370 0.985 0.820 1.055 ;
        RECT  0.440 0.240 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDQD1BWP

MACRO LHSNDQD2BWP
    CLASS CORE ;
    FOREIGN LHSNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.055 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.735 2.415 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.535 -0.115 2.610 0.305 ;
        RECT  2.250 -0.115 2.535 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.520 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.975 2.610 1.375 ;
        RECT  2.250 1.145 2.530 1.375 ;
        RECT  2.170 0.885 2.250 1.375 ;
        RECT  1.900 1.145 2.170 1.375 ;
        RECT  1.800 0.990 1.900 1.375 ;
        RECT  0.730 1.145 1.800 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.345 0.620 ;
        RECT  2.200 0.395 2.270 0.805 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.735 2.200 0.805 ;
        RECT  1.925 0.545 2.120 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.735 2.070 1.055 ;
        RECT  1.855 0.275 1.925 0.915 ;
        RECT  1.770 0.275 1.855 0.355 ;
        RECT  1.710 0.845 1.855 0.915 ;
        RECT  1.630 0.845 1.710 1.055 ;
        RECT  1.420 0.985 1.630 1.055 ;
        RECT  1.425 0.540 1.620 0.620 ;
        RECT  1.345 0.205 1.425 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  0.960 0.205 1.345 0.275 ;
        RECT  0.930 0.845 1.345 0.915 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.370 0.985 0.820 1.055 ;
        RECT  0.440 0.240 0.510 0.905 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.050 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDQD2BWP

MACRO LHSNDQD4BWP
    CLASS CORE ;
    FOREIGN LHSNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.185 2.845 0.465 ;
        RECT  2.835 0.775 2.845 1.055 ;
        RECT  2.775 0.185 2.835 1.055 ;
        RECT  2.625 0.355 2.775 0.905 ;
        RECT  2.485 0.355 2.625 0.465 ;
        RECT  2.485 0.775 2.625 0.905 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.775 2.485 1.055 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.485 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.275 ;
        RECT  2.310 -0.115 2.570 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.960 -0.115 2.230 0.115 ;
        RECT  1.860 -0.115 1.960 0.275 ;
        RECT  1.445 -0.115 1.860 0.115 ;
        RECT  1.300 -0.115 1.445 0.280 ;
        RECT  0.680 -0.115 1.300 0.115 ;
        RECT  0.585 -0.115 0.680 0.265 ;
        RECT  0.310 -0.115 0.585 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.665 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 0.985 2.690 1.375 ;
        RECT  2.300 1.145 2.570 1.375 ;
        RECT  2.220 0.925 2.300 1.375 ;
        RECT  1.925 1.145 2.220 1.375 ;
        RECT  1.790 0.990 1.925 1.375 ;
        RECT  0.730 1.145 1.790 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.355 2.555 0.465 ;
        RECT  2.485 0.775 2.555 0.905 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.775 2.485 1.055 ;
        RECT  2.345 0.545 2.535 0.620 ;
        RECT  2.275 0.385 2.345 0.805 ;
        RECT  2.130 0.385 2.275 0.465 ;
        RECT  2.110 0.735 2.275 0.805 ;
        RECT  1.935 0.545 2.195 0.620 ;
        RECT  2.050 0.185 2.130 0.465 ;
        RECT  2.035 0.735 2.110 1.055 ;
        RECT  1.865 0.345 1.935 0.905 ;
        RECT  1.650 0.345 1.865 0.415 ;
        RECT  1.660 0.835 1.865 0.905 ;
        RECT  1.580 0.835 1.660 1.055 ;
        RECT  1.370 0.985 1.580 1.055 ;
        RECT  1.435 0.355 1.510 0.915 ;
        RECT  1.205 0.355 1.435 0.425 ;
        RECT  0.930 0.845 1.435 0.915 ;
        RECT  1.200 0.985 1.370 1.070 ;
        RECT  0.960 0.690 1.210 0.775 ;
        RECT  1.135 0.195 1.205 0.425 ;
        RECT  0.910 0.195 1.135 0.270 ;
        RECT  0.885 0.340 0.960 0.775 ;
        RECT  0.840 0.985 0.960 1.075 ;
        RECT  0.515 0.695 0.885 0.775 ;
        RECT  0.370 0.985 0.840 1.055 ;
        RECT  0.510 0.200 0.515 0.775 ;
        RECT  0.440 0.200 0.510 0.905 ;
        RECT  0.390 0.200 0.440 0.270 ;
        RECT  0.300 0.350 0.370 1.055 ;
        RECT  0.130 0.350 0.300 0.420 ;
        RECT  0.125 0.985 0.300 1.055 ;
        RECT  0.055 0.260 0.130 0.420 ;
        RECT  0.055 0.860 0.125 1.055 ;
    END
END LHSNDQD4BWP

MACRO LHSNQD1BWP
    CLASS CORE ;
    FOREIGN LHSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.375 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.355 2.065 0.905 ;
        RECT  1.995 0.185 2.030 1.060 ;
        RECT  1.950 0.185 1.995 0.465 ;
        RECT  1.950 0.740 1.995 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0170 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.115 2.100 0.115 ;
        RECT  1.760 -0.115 1.840 0.290 ;
        RECT  1.070 -0.115 1.760 0.115 ;
        RECT  0.990 -0.115 1.070 0.440 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.145 2.100 1.375 ;
        RECT  1.770 0.800 1.850 1.375 ;
        RECT  1.470 1.145 1.770 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.545 1.920 0.620 ;
        RECT  1.620 0.205 1.690 1.050 ;
        RECT  1.530 0.205 1.620 0.275 ;
        RECT  1.550 0.980 1.620 1.050 ;
        RECT  1.460 0.345 1.540 0.910 ;
        RECT  1.330 0.345 1.460 0.415 ;
        RECT  1.290 0.840 1.460 0.910 ;
        RECT  1.210 0.840 1.290 1.055 ;
        RECT  0.840 0.985 1.210 1.055 ;
        RECT  0.975 0.545 1.200 0.615 ;
        RECT  0.905 0.545 0.975 0.915 ;
        RECT  0.865 0.545 0.905 0.615 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.615 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.130 0.960 0.450 1.030 ;
        RECT  0.105 0.890 0.130 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSNQD1BWP

MACRO LHSNQD2BWP
    CLASS CORE ;
    FOREIGN LHSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.375 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.355 2.065 0.905 ;
        RECT  1.995 0.185 2.010 1.060 ;
        RECT  1.930 0.185 1.995 0.465 ;
        RECT  1.930 0.740 1.995 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0170 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 -0.115 2.240 0.115 ;
        RECT  2.100 -0.115 2.200 0.290 ;
        RECT  1.830 -0.115 2.100 0.115 ;
        RECT  1.760 -0.115 1.830 0.450 ;
        RECT  1.070 -0.115 1.760 0.115 ;
        RECT  0.990 -0.115 1.070 0.440 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.145 2.240 1.375 ;
        RECT  2.100 0.985 2.200 1.375 ;
        RECT  1.830 1.145 2.100 1.375 ;
        RECT  1.760 0.800 1.830 1.375 ;
        RECT  1.470 1.145 1.760 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.545 1.910 0.620 ;
        RECT  1.620 0.205 1.690 1.050 ;
        RECT  1.510 0.205 1.620 0.275 ;
        RECT  1.550 0.980 1.620 1.050 ;
        RECT  1.460 0.345 1.540 0.910 ;
        RECT  1.330 0.345 1.460 0.415 ;
        RECT  1.290 0.840 1.460 0.910 ;
        RECT  1.210 0.840 1.290 1.055 ;
        RECT  0.840 0.985 1.210 1.055 ;
        RECT  0.975 0.545 1.200 0.615 ;
        RECT  0.905 0.545 0.975 0.915 ;
        RECT  0.865 0.545 0.905 0.615 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.615 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.130 0.960 0.450 1.030 ;
        RECT  0.105 0.890 0.130 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSNQD2BWP

MACRO LHSNQD4BWP
    CLASS CORE ;
    FOREIGN LHSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.375 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.275 0.355 2.350 0.485 ;
        RECT  2.275 0.760 2.350 0.905 ;
        RECT  2.070 0.355 2.275 0.905 ;
        RECT  2.065 0.355 2.070 1.040 ;
        RECT  1.980 0.185 2.065 0.475 ;
        RECT  1.980 0.760 2.065 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0392 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.685 0.830 0.775 ;
        RECT  0.590 0.355 0.665 0.775 ;
        RECT  0.500 0.355 0.590 0.440 ;
        RECT  0.245 0.705 0.590 0.775 ;
        RECT  0.175 0.495 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0170 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.540 0.480 0.625 ;
        RECT  0.315 0.355 0.390 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.485 ;
        RECT  2.270 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.270 0.280 ;
        RECT  1.860 -0.115 2.150 0.115 ;
        RECT  1.780 -0.115 1.860 0.465 ;
        RECT  1.050 -0.115 1.780 0.115 ;
        RECT  0.970 -0.115 1.050 0.440 ;
        RECT  0.340 -0.115 0.970 0.115 ;
        RECT  0.240 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.665 2.610 1.375 ;
        RECT  2.270 1.145 2.530 1.375 ;
        RECT  2.150 1.005 2.270 1.375 ;
        RECT  1.860 1.145 2.150 1.375 ;
        RECT  1.780 0.800 1.860 1.375 ;
        RECT  1.470 1.145 1.780 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.345 0.355 2.350 0.485 ;
        RECT  2.345 0.760 2.350 0.905 ;
        RECT  1.980 0.185 1.995 0.475 ;
        RECT  1.980 0.760 1.995 1.040 ;
        RECT  1.710 0.545 1.970 0.615 ;
        RECT  1.640 0.205 1.710 1.050 ;
        RECT  1.550 0.205 1.640 0.275 ;
        RECT  1.550 0.980 1.640 1.050 ;
        RECT  1.490 0.345 1.570 0.910 ;
        RECT  1.350 0.345 1.490 0.415 ;
        RECT  1.290 0.840 1.490 0.910 ;
        RECT  1.210 0.840 1.290 1.055 ;
        RECT  0.840 0.985 1.210 1.055 ;
        RECT  0.975 0.545 1.200 0.615 ;
        RECT  0.905 0.545 0.975 0.915 ;
        RECT  0.865 0.545 0.905 0.615 ;
        RECT  0.590 0.845 0.905 0.915 ;
        RECT  0.795 0.195 0.865 0.615 ;
        RECT  0.570 0.195 0.795 0.265 ;
        RECT  0.520 1.005 0.630 1.075 ;
        RECT  0.450 0.960 0.520 1.075 ;
        RECT  0.130 0.960 0.450 1.030 ;
        RECT  0.105 0.890 0.130 1.030 ;
        RECT  0.105 0.220 0.125 0.380 ;
        RECT  0.035 0.220 0.105 1.030 ;
    END
END LHSNQD4BWP

MACRO LNCND1BWP
    CLASS CORE ;
    FOREIGN LNCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.710 2.290 0.780 ;
        RECT  2.205 0.185 2.245 0.465 ;
        RECT  2.135 0.185 2.205 0.780 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.195 2.625 1.070 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.390 0.485 ;
        RECT  1.090 0.345 1.295 0.415 ;
        RECT  1.015 0.345 1.090 0.625 ;
        RECT  0.750 0.345 1.015 0.415 ;
        RECT  0.680 0.205 0.750 0.415 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.115 2.660 0.115 ;
        RECT  2.350 -0.115 2.430 0.440 ;
        RECT  2.065 -0.115 2.350 0.115 ;
        RECT  1.990 -0.115 2.065 0.300 ;
        RECT  1.530 -0.115 1.990 0.115 ;
        RECT  1.400 -0.115 1.530 0.135 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.145 2.660 1.375 ;
        RECT  2.340 0.990 2.440 1.375 ;
        RECT  2.080 1.145 2.340 1.375 ;
        RECT  1.980 0.990 2.080 1.375 ;
        RECT  1.520 1.145 1.980 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.380 0.520 2.460 0.920 ;
        RECT  2.030 0.850 2.380 0.920 ;
        RECT  1.960 0.380 2.030 0.920 ;
        RECT  1.890 0.380 1.960 0.465 ;
        RECT  1.890 0.720 1.960 0.920 ;
        RECT  1.810 0.185 1.890 0.465 ;
        RECT  1.810 0.720 1.890 1.040 ;
        RECT  1.715 0.545 1.880 0.615 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.205 1.550 0.920 ;
        RECT  0.830 0.205 1.480 0.275 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.805 0.705 1.250 0.775 ;
        RECT  0.805 0.490 0.945 0.580 ;
        RECT  0.735 0.490 0.805 0.775 ;
        RECT  0.385 0.705 0.735 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCND1BWP

MACRO LNCND2BWP
    CLASS CORE ;
    FOREIGN LNCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.345 0.780 ;
        RECT  2.270 0.355 2.275 0.465 ;
        RECT  2.190 0.660 2.275 0.780 ;
        RECT  2.190 0.185 2.270 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.355 2.765 0.765 ;
        RECT  2.695 0.185 2.700 1.045 ;
        RECT  2.620 0.185 2.695 0.470 ;
        RECT  2.620 0.695 2.695 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.300 ;
        RECT  2.495 -0.115 2.810 0.115 ;
        RECT  2.415 -0.115 2.495 0.440 ;
        RECT  2.070 -0.115 2.415 0.115 ;
        RECT  1.990 -0.115 2.070 0.300 ;
        RECT  1.530 -0.115 1.990 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.850 2.900 1.375 ;
        RECT  2.490 1.145 2.800 1.375 ;
        RECT  2.390 0.990 2.490 1.375 ;
        RECT  2.080 1.145 2.390 1.375 ;
        RECT  1.980 0.990 2.080 1.375 ;
        RECT  1.520 1.145 1.980 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.505 0.540 2.610 0.620 ;
        RECT  2.425 0.540 2.505 0.920 ;
        RECT  2.120 0.850 2.425 0.920 ;
        RECT  2.050 0.380 2.120 0.920 ;
        RECT  1.890 0.380 2.050 0.465 ;
        RECT  1.890 0.850 2.050 0.920 ;
        RECT  1.715 0.545 1.980 0.620 ;
        RECT  1.810 0.185 1.890 0.465 ;
        RECT  1.810 0.720 1.890 1.040 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCND2BWP

MACRO LNCND4BWP
    CLASS CORE ;
    FOREIGN LNCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.700 2.850 0.800 ;
        RECT  2.755 0.185 2.825 0.485 ;
        RECT  2.695 0.355 2.755 0.485 ;
        RECT  2.485 0.355 2.695 0.800 ;
        RECT  2.465 0.355 2.485 0.485 ;
        RECT  2.370 0.700 2.485 0.800 ;
        RECT  2.395 0.185 2.465 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.185 3.545 0.465 ;
        RECT  3.535 0.735 3.545 1.035 ;
        RECT  3.475 0.185 3.535 1.035 ;
        RECT  3.325 0.355 3.475 0.905 ;
        RECT  3.185 0.355 3.325 0.465 ;
        RECT  3.185 0.735 3.325 0.905 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.735 3.185 1.035 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0374 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.460 ;
        RECT  3.380 -0.115 3.650 0.115 ;
        RECT  3.280 -0.115 3.380 0.275 ;
        RECT  3.010 -0.115 3.280 0.115 ;
        RECT  2.930 -0.115 3.010 0.460 ;
        RECT  2.660 -0.115 2.930 0.115 ;
        RECT  2.560 -0.115 2.660 0.275 ;
        RECT  2.290 -0.115 2.560 0.115 ;
        RECT  2.210 -0.115 2.290 0.320 ;
        RECT  1.900 -0.115 2.210 0.115 ;
        RECT  1.820 -0.115 1.900 0.460 ;
        RECT  1.530 -0.115 1.820 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.665 3.730 1.375 ;
        RECT  3.380 1.145 3.650 1.375 ;
        RECT  3.280 0.985 3.380 1.375 ;
        RECT  3.030 1.145 3.280 1.375 ;
        RECT  2.910 1.010 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 1.010 2.670 1.375 ;
        RECT  2.310 1.145 2.550 1.375 ;
        RECT  2.190 1.010 2.310 1.375 ;
        RECT  1.920 1.145 2.190 1.375 ;
        RECT  1.840 0.745 1.920 1.375 ;
        RECT  1.520 1.145 1.840 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.355 3.255 0.465 ;
        RECT  3.185 0.735 3.255 0.905 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.735 3.185 1.035 ;
        RECT  2.765 0.700 2.850 0.800 ;
        RECT  2.765 0.185 2.825 0.485 ;
        RECT  2.395 0.185 2.415 0.485 ;
        RECT  2.370 0.700 2.415 0.800 ;
        RECT  3.000 0.540 3.230 0.620 ;
        RECT  2.930 0.540 3.000 0.940 ;
        RECT  2.170 0.870 2.930 0.940 ;
        RECT  2.110 0.395 2.170 0.940 ;
        RECT  2.100 0.185 2.110 1.065 ;
        RECT  2.030 0.185 2.100 0.465 ;
        RECT  2.030 0.745 2.100 1.065 ;
        RECT  1.730 0.540 2.020 0.620 ;
        RECT  1.725 0.540 1.730 1.060 ;
        RECT  1.650 0.185 1.725 1.060 ;
        RECT  1.630 0.185 1.650 0.465 ;
        RECT  1.370 0.990 1.650 1.060 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.200 0.120 0.555 ;
        RECT  0.035 0.200 0.105 1.075 ;
    END
END LNCND4BWP

MACRO LNCNDD1BWP
    CLASS CORE ;
    FOREIGN LNCNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.710 2.570 0.780 ;
        RECT  2.485 0.185 2.525 0.465 ;
        RECT  2.415 0.185 2.485 0.780 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.815 0.195 2.905 1.070 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.940 0.115 ;
        RECT  2.630 -0.115 2.710 0.440 ;
        RECT  2.345 -0.115 2.630 0.115 ;
        RECT  2.270 -0.115 2.345 0.300 ;
        RECT  1.810 -0.115 2.270 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 2.940 1.375 ;
        RECT  2.620 0.990 2.720 1.375 ;
        RECT  2.360 1.145 2.620 1.375 ;
        RECT  2.260 0.990 2.360 1.375 ;
        RECT  1.800 1.145 2.260 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.520 2.740 0.920 ;
        RECT  2.280 0.850 2.660 0.920 ;
        RECT  2.210 0.380 2.280 0.920 ;
        RECT  2.170 0.380 2.210 0.465 ;
        RECT  2.170 0.720 2.210 0.920 ;
        RECT  2.090 0.185 2.170 0.465 ;
        RECT  2.090 0.720 2.170 1.040 ;
        RECT  1.995 0.545 2.140 0.615 ;
        RECT  1.925 0.185 1.995 1.060 ;
        RECT  1.915 0.185 1.925 0.465 ;
        RECT  1.915 0.730 1.925 1.060 ;
        RECT  1.650 0.985 1.915 1.060 ;
        RECT  1.830 0.520 1.855 0.640 ;
        RECT  1.760 0.210 1.830 0.915 ;
        RECT  1.110 0.210 1.760 0.280 ;
        RECT  0.590 0.845 1.760 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDD1BWP

MACRO LNCNDD2BWP
    CLASS CORE ;
    FOREIGN LNCNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.185 2.490 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.055 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.735 2.835 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.115 3.080 0.115 ;
        RECT  2.955 -0.115 3.025 0.305 ;
        RECT  2.670 -0.115 2.955 0.115 ;
        RECT  2.590 -0.115 2.670 0.465 ;
        RECT  2.310 -0.115 2.590 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.780 -0.115 2.230 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 1.145 3.080 1.375 ;
        RECT  2.955 0.960 3.025 1.375 ;
        RECT  2.690 1.145 2.955 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  0.910 1.145 2.210 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.615 ;
        RECT  2.595 0.545 2.665 0.935 ;
        RECT  2.240 0.865 2.595 0.935 ;
        RECT  2.170 0.385 2.240 0.935 ;
        RECT  2.130 0.385 2.170 0.465 ;
        RECT  2.130 0.735 2.170 0.935 ;
        RECT  2.050 0.185 2.130 0.465 ;
        RECT  2.050 0.735 2.130 1.055 ;
        RECT  1.955 0.545 2.100 0.620 ;
        RECT  1.885 0.185 1.955 1.055 ;
        RECT  1.875 0.185 1.885 0.465 ;
        RECT  1.875 0.775 1.885 1.055 ;
        RECT  1.670 0.985 1.875 1.055 ;
        RECT  1.795 0.520 1.815 0.640 ;
        RECT  1.725 0.205 1.795 0.915 ;
        RECT  1.090 0.205 1.725 0.275 ;
        RECT  0.590 0.845 1.725 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.410 0.195 0.490 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.245 0.350 0.410 0.420 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDD2BWP

MACRO LNCNDD4BWP
    CLASS CORE ;
    FOREIGN LNCNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.705 3.130 0.795 ;
        RECT  3.035 0.185 3.105 0.485 ;
        RECT  2.975 0.355 3.035 0.485 ;
        RECT  2.765 0.355 2.975 0.795 ;
        RECT  2.745 0.355 2.765 0.485 ;
        RECT  2.650 0.705 2.765 0.795 ;
        RECT  2.675 0.185 2.745 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.825 0.465 ;
        RECT  3.815 0.775 3.825 1.055 ;
        RECT  3.755 0.185 3.815 1.055 ;
        RECT  3.605 0.355 3.755 0.905 ;
        RECT  3.465 0.355 3.605 0.465 ;
        RECT  3.465 0.775 3.605 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 0.345 1.680 0.485 ;
        RECT  0.665 0.345 1.600 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.485 ;
        RECT  3.670 -0.115 3.930 0.115 ;
        RECT  3.550 -0.115 3.670 0.275 ;
        RECT  3.290 -0.115 3.550 0.115 ;
        RECT  3.210 -0.115 3.290 0.465 ;
        RECT  2.950 -0.115 3.210 0.115 ;
        RECT  2.830 -0.115 2.950 0.275 ;
        RECT  2.570 -0.115 2.830 0.115 ;
        RECT  2.490 -0.115 2.570 0.305 ;
        RECT  2.200 -0.115 2.490 0.115 ;
        RECT  2.120 -0.115 2.200 0.465 ;
        RECT  1.820 -0.115 2.120 0.115 ;
        RECT  1.700 -0.115 1.820 0.135 ;
        RECT  0.700 -0.115 1.700 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.665 4.010 1.375 ;
        RECT  3.670 1.145 3.930 1.375 ;
        RECT  3.550 0.985 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 1.005 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 1.005 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 1.005 2.590 1.375 ;
        RECT  2.200 1.145 2.470 1.375 ;
        RECT  2.120 0.755 2.200 1.375 ;
        RECT  1.800 1.145 2.120 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.355 3.535 0.465 ;
        RECT  3.465 0.775 3.535 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        RECT  3.045 0.705 3.130 0.795 ;
        RECT  3.045 0.185 3.105 0.485 ;
        RECT  2.675 0.185 2.695 0.485 ;
        RECT  2.650 0.705 2.695 0.795 ;
        RECT  3.285 0.540 3.515 0.620 ;
        RECT  3.215 0.540 3.285 0.935 ;
        RECT  2.530 0.865 3.215 0.935 ;
        RECT  2.460 0.385 2.530 0.935 ;
        RECT  2.390 0.385 2.460 0.465 ;
        RECT  2.390 0.735 2.460 0.935 ;
        RECT  2.310 0.185 2.390 0.465 ;
        RECT  2.310 0.735 2.390 1.055 ;
        RECT  2.050 0.545 2.380 0.620 ;
        RECT  1.980 0.280 2.050 1.055 ;
        RECT  1.930 0.280 1.980 0.440 ;
        RECT  1.930 0.775 1.980 1.055 ;
        RECT  1.650 0.985 1.930 1.055 ;
        RECT  1.840 0.520 1.910 0.640 ;
        RECT  1.770 0.205 1.840 0.915 ;
        RECT  1.110 0.205 1.770 0.275 ;
        RECT  0.590 0.845 1.770 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.200 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDD4BWP

MACRO LNCNDQD1BWP
    CLASS CORE ;
    FOREIGN LNCNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.625 1.045 ;
        RECT  2.535 0.185 2.555 0.465 ;
        RECT  2.535 0.725 2.555 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.420 -0.115 2.660 0.115 ;
        RECT  2.340 -0.115 2.420 0.305 ;
        RECT  1.810 -0.115 2.340 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.420 1.145 2.660 1.375 ;
        RECT  2.340 0.925 2.420 1.375 ;
        RECT  1.800 1.145 2.340 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.465 0.520 2.485 0.640 ;
        RECT  2.395 0.385 2.465 0.805 ;
        RECT  2.230 0.385 2.395 0.465 ;
        RECT  2.230 0.735 2.395 0.805 ;
        RECT  1.990 0.545 2.310 0.615 ;
        RECT  2.150 0.185 2.230 0.465 ;
        RECT  2.150 0.735 2.230 1.055 ;
        RECT  1.920 0.195 1.990 1.060 ;
        RECT  1.650 0.985 1.920 1.060 ;
        RECT  1.830 0.520 1.850 0.640 ;
        RECT  1.760 0.210 1.830 0.915 ;
        RECT  1.110 0.210 1.760 0.280 ;
        RECT  0.590 0.845 1.760 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDQD1BWP

MACRO LNCNDQD2BWP
    CLASS CORE ;
    FOREIGN LNCNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.355 2.625 0.905 ;
        RECT  2.565 0.355 2.570 1.055 ;
        RECT  2.555 0.185 2.565 1.055 ;
        RECT  2.490 0.185 2.555 0.465 ;
        RECT  2.490 0.735 2.555 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.745 -0.115 2.800 0.115 ;
        RECT  2.675 -0.115 2.745 0.305 ;
        RECT  2.360 -0.115 2.675 0.115 ;
        RECT  2.280 -0.115 2.360 0.305 ;
        RECT  1.780 -0.115 2.280 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.745 1.145 2.800 1.375 ;
        RECT  2.675 0.960 2.745 1.375 ;
        RECT  2.360 1.145 2.675 1.375 ;
        RECT  2.280 0.915 2.360 1.375 ;
        RECT  0.910 1.145 2.280 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.420 0.520 2.440 0.640 ;
        RECT  2.350 0.385 2.420 0.805 ;
        RECT  2.165 0.385 2.350 0.465 ;
        RECT  2.170 0.735 2.350 0.805 ;
        RECT  1.970 0.545 2.200 0.620 ;
        RECT  2.090 0.735 2.170 1.055 ;
        RECT  2.095 0.185 2.165 0.465 ;
        RECT  1.890 0.195 1.970 1.055 ;
        RECT  1.670 0.985 1.890 1.055 ;
        RECT  1.740 0.205 1.815 0.915 ;
        RECT  1.090 0.205 1.740 0.275 ;
        RECT  0.590 0.845 1.740 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.410 0.195 0.490 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.245 0.350 0.410 0.420 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDQD2BWP

MACRO LNCNDQD4BWP
    CLASS CORE ;
    FOREIGN LNCNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.775 3.125 1.055 ;
        RECT  3.055 0.185 3.115 1.055 ;
        RECT  2.905 0.355 3.055 0.905 ;
        RECT  2.765 0.355 2.905 0.465 ;
        RECT  2.765 0.775 2.905 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.345 1.670 0.485 ;
        RECT  0.665 0.345 1.590 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.485 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.275 ;
        RECT  2.560 -0.115 2.850 0.115 ;
        RECT  2.475 -0.115 2.560 0.305 ;
        RECT  2.170 -0.115 2.475 0.115 ;
        RECT  2.090 -0.115 2.170 0.465 ;
        RECT  1.800 -0.115 2.090 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.665 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.985 2.970 1.375 ;
        RECT  2.560 1.145 2.850 1.375 ;
        RECT  2.480 0.925 2.560 1.375 ;
        RECT  2.170 1.145 2.480 1.375 ;
        RECT  2.090 0.755 2.170 1.375 ;
        RECT  1.800 1.145 2.090 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.465 ;
        RECT  2.765 0.775 2.835 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        RECT  2.625 0.545 2.815 0.620 ;
        RECT  2.555 0.385 2.625 0.845 ;
        RECT  2.360 0.385 2.555 0.465 ;
        RECT  2.360 0.735 2.555 0.845 ;
        RECT  1.990 0.545 2.390 0.620 ;
        RECT  2.280 0.185 2.360 0.465 ;
        RECT  2.280 0.735 2.360 1.055 ;
        RECT  1.910 0.195 1.990 1.055 ;
        RECT  1.650 0.985 1.910 1.055 ;
        RECT  1.760 0.205 1.840 0.915 ;
        RECT  1.110 0.205 1.760 0.275 ;
        RECT  0.590 0.845 1.760 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.200 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCNDQD4BWP

MACRO LNCNQD1BWP
    CLASS CORE ;
    FOREIGN LNCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.345 1.045 ;
        RECT  2.250 0.185 2.275 0.465 ;
        RECT  2.250 0.705 2.275 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.040 -0.115 2.120 0.325 ;
        RECT  1.530 -0.115 2.040 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.040 0.780 2.120 1.375 ;
        RECT  1.520 1.145 2.040 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 0.540 2.205 0.620 ;
        RECT  1.900 0.205 1.970 1.065 ;
        RECT  1.810 0.205 1.900 0.285 ;
        RECT  1.810 0.985 1.900 1.065 ;
        RECT  1.715 0.545 1.830 0.620 ;
        RECT  1.645 0.185 1.715 1.060 ;
        RECT  1.635 0.185 1.645 0.465 ;
        RECT  1.635 0.730 1.645 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCNQD1BWP

MACRO LNCNQD2BWP
    CLASS CORE ;
    FOREIGN LNCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.355 2.345 0.765 ;
        RECT  2.275 0.185 2.290 1.050 ;
        RECT  2.210 0.185 2.275 0.465 ;
        RECT  2.210 0.695 2.275 1.050 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.290 ;
        RECT  2.100 -0.115 2.390 0.115 ;
        RECT  2.020 -0.115 2.100 0.300 ;
        RECT  1.530 -0.115 2.020 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.850 2.480 1.375 ;
        RECT  2.100 1.145 2.380 1.375 ;
        RECT  2.020 0.880 2.100 1.375 ;
        RECT  1.520 1.145 2.020 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.130 0.545 2.195 0.615 ;
        RECT  2.060 0.380 2.130 0.800 ;
        RECT  1.910 0.380 2.060 0.465 ;
        RECT  1.910 0.720 2.060 0.800 ;
        RECT  1.710 0.545 1.980 0.615 ;
        RECT  1.830 0.185 1.910 0.465 ;
        RECT  1.830 0.720 1.910 1.040 ;
        RECT  1.635 0.185 1.710 1.060 ;
        RECT  1.370 0.990 1.635 1.060 ;
        RECT  1.485 0.210 1.555 0.920 ;
        RECT  0.830 0.210 1.485 0.280 ;
        RECT  0.370 0.850 1.485 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCNQD2BWP

MACRO LNCNQD4BWP
    CLASS CORE ;
    FOREIGN LNCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.185 2.850 0.485 ;
        RECT  2.770 0.760 2.850 1.040 ;
        RECT  2.695 0.355 2.770 0.485 ;
        RECT  2.695 0.760 2.770 0.905 ;
        RECT  2.485 0.355 2.695 0.905 ;
        RECT  2.455 0.355 2.485 0.485 ;
        RECT  2.450 0.760 2.485 0.905 ;
        RECT  2.370 0.185 2.455 0.485 ;
        RECT  2.370 0.760 2.450 1.040 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0374 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.465 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.670 0.275 ;
        RECT  2.260 -0.115 2.570 0.115 ;
        RECT  2.180 -0.115 2.260 0.460 ;
        RECT  1.890 -0.115 2.180 0.115 ;
        RECT  1.810 -0.115 1.890 0.460 ;
        RECT  1.530 -0.115 1.810 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.685 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.570 0.985 2.670 1.375 ;
        RECT  2.260 1.145 2.570 1.375 ;
        RECT  2.180 0.750 2.260 1.375 ;
        RECT  1.890 1.145 2.180 1.375 ;
        RECT  1.810 0.750 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.770 0.185 2.850 0.485 ;
        RECT  2.770 0.760 2.850 1.040 ;
        RECT  2.765 0.355 2.770 0.485 ;
        RECT  2.765 0.760 2.770 0.905 ;
        RECT  2.370 0.185 2.415 0.485 ;
        RECT  2.370 0.760 2.415 1.040 ;
        RECT  2.070 0.560 2.380 0.630 ;
        RECT  1.990 0.185 2.070 1.060 ;
        RECT  1.710 0.540 1.910 0.620 ;
        RECT  1.630 0.185 1.710 1.060 ;
        RECT  1.370 0.990 1.630 1.060 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.200 0.120 0.555 ;
        RECT  0.035 0.200 0.105 1.075 ;
    END
END LNCNQD4BWP

MACRO LNCSND1BWP
    CLASS CORE ;
    FOREIGN LNCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.950 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.720 2.550 0.790 ;
        RECT  2.485 0.185 2.515 0.465 ;
        RECT  2.410 0.185 2.485 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.185 2.905 1.045 ;
        RECT  2.815 0.185 2.835 0.465 ;
        RECT  2.815 0.745 2.835 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 -0.115 2.940 0.115 ;
        RECT  2.620 -0.115 2.700 0.375 ;
        RECT  2.170 -0.115 2.620 0.115 ;
        RECT  2.050 -0.115 2.170 0.275 ;
        RECT  1.530 -0.115 2.050 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.145 2.940 1.375 ;
        RECT  2.600 1.020 2.720 1.375 ;
        RECT  2.110 1.145 2.600 1.375 ;
        RECT  2.010 0.990 2.110 1.375 ;
        RECT  1.520 1.145 2.010 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.705 0.520 2.765 0.640 ;
        RECT  2.635 0.520 2.705 0.940 ;
        RECT  2.330 0.870 2.635 0.940 ;
        RECT  2.250 0.185 2.330 1.045 ;
        RECT  2.090 0.345 2.170 0.910 ;
        RECT  1.810 0.345 2.090 0.415 ;
        RECT  1.890 0.840 2.090 0.910 ;
        RECT  1.810 0.840 1.890 1.060 ;
        RECT  1.370 0.990 1.810 1.060 ;
        RECT  1.520 0.210 1.600 0.920 ;
        RECT  0.830 0.210 1.520 0.280 ;
        RECT  0.370 0.850 1.520 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCSND1BWP

MACRO LNCSND2BWP
    CLASS CORE ;
    FOREIGN LNCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.805 0.495 1.855 0.640 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.400 0.185 2.485 0.820 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.060 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.740 2.835 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 -0.115 3.080 0.115 ;
        RECT  2.940 -0.115 3.040 0.290 ;
        RECT  2.660 -0.115 2.940 0.115 ;
        RECT  2.580 -0.115 2.660 0.465 ;
        RECT  2.300 -0.115 2.580 0.115 ;
        RECT  2.180 -0.115 2.300 0.135 ;
        RECT  1.530 -0.115 2.180 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.985 3.030 1.375 ;
        RECT  2.680 1.145 2.950 1.375 ;
        RECT  2.560 1.040 2.680 1.375 ;
        RECT  2.305 1.145 2.560 1.375 ;
        RECT  2.185 1.040 2.305 1.375 ;
        RECT  1.910 1.145 2.185 1.375 ;
        RECT  1.830 0.960 1.910 1.375 ;
        RECT  1.520 1.145 1.830 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.620 ;
        RECT  2.590 0.545 2.665 0.970 ;
        RECT  2.090 0.900 2.590 0.970 ;
        RECT  2.190 0.205 2.270 0.660 ;
        RECT  1.730 0.205 2.190 0.275 ;
        RECT  2.010 0.345 2.090 0.970 ;
        RECT  1.655 0.205 1.730 1.060 ;
        RECT  1.370 0.990 1.655 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCSND2BWP

MACRO LNCSND4BWP
    CLASS CORE ;
    FOREIGN LNCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.700 3.270 0.800 ;
        RECT  3.175 0.185 3.245 0.485 ;
        RECT  3.115 0.355 3.175 0.485 ;
        RECT  2.905 0.355 3.115 0.800 ;
        RECT  2.885 0.355 2.905 0.485 ;
        RECT  2.790 0.700 2.905 0.800 ;
        RECT  2.815 0.185 2.885 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.465 ;
        RECT  3.955 0.735 3.965 1.035 ;
        RECT  3.895 0.185 3.955 1.035 ;
        RECT  3.745 0.355 3.895 0.905 ;
        RECT  3.605 0.355 3.745 0.465 ;
        RECT  3.605 0.735 3.745 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.735 3.605 1.035 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0374 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.460 ;
        RECT  3.800 -0.115 4.070 0.115 ;
        RECT  3.700 -0.115 3.800 0.275 ;
        RECT  3.430 -0.115 3.700 0.115 ;
        RECT  3.350 -0.115 3.430 0.460 ;
        RECT  3.080 -0.115 3.350 0.115 ;
        RECT  2.980 -0.115 3.080 0.275 ;
        RECT  2.710 -0.115 2.980 0.115 ;
        RECT  2.630 -0.115 2.710 0.315 ;
        RECT  2.340 -0.115 2.630 0.115 ;
        RECT  2.220 -0.115 2.340 0.265 ;
        RECT  1.520 -0.115 2.220 0.115 ;
        RECT  1.400 -0.115 1.520 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.070 0.665 4.150 1.375 ;
        RECT  3.800 1.145 4.070 1.375 ;
        RECT  3.700 0.985 3.800 1.375 ;
        RECT  3.450 1.145 3.700 1.375 ;
        RECT  3.330 1.010 3.450 1.375 ;
        RECT  3.090 1.145 3.330 1.375 ;
        RECT  2.970 1.010 3.090 1.375 ;
        RECT  2.730 1.145 2.970 1.375 ;
        RECT  2.610 1.010 2.730 1.375 ;
        RECT  2.340 1.145 2.610 1.375 ;
        RECT  2.220 1.000 2.340 1.375 ;
        RECT  1.920 1.145 2.220 1.375 ;
        RECT  1.800 1.000 1.920 1.375 ;
        RECT  1.520 1.145 1.800 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.355 3.675 0.465 ;
        RECT  3.605 0.735 3.675 0.905 ;
        RECT  3.535 0.185 3.605 0.465 ;
        RECT  3.535 0.735 3.605 1.035 ;
        RECT  3.185 0.700 3.270 0.800 ;
        RECT  3.185 0.185 3.245 0.485 ;
        RECT  2.815 0.185 2.835 0.485 ;
        RECT  2.790 0.700 2.835 0.800 ;
        RECT  3.420 0.540 3.650 0.620 ;
        RECT  3.350 0.540 3.420 0.940 ;
        RECT  2.720 0.870 3.350 0.940 ;
        RECT  2.650 0.395 2.720 0.940 ;
        RECT  2.525 0.395 2.650 0.465 ;
        RECT  2.530 0.870 2.650 0.940 ;
        RECT  2.380 0.545 2.580 0.625 ;
        RECT  2.450 0.740 2.530 1.060 ;
        RECT  2.455 0.185 2.525 0.465 ;
        RECT  2.310 0.345 2.380 0.920 ;
        RECT  1.920 0.345 2.310 0.415 ;
        RECT  1.710 0.850 2.310 0.920 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.200 0.120 0.555 ;
        RECT  0.035 0.200 0.105 1.075 ;
        RECT  2.100 0.500 2.180 0.780 ;
        RECT  1.600 0.710 2.100 0.780 ;
        RECT  1.800 0.205 1.920 0.415 ;
        RECT  1.630 0.850 1.710 1.060 ;
        RECT  1.370 0.990 1.630 1.060 ;
        RECT  1.550 0.520 1.600 0.780 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
    END
END LNCSND4BWP

MACRO LNCSNDD1BWP
    CLASS CORE ;
    FOREIGN LNCSNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.230 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.720 2.830 0.790 ;
        RECT  2.765 0.185 2.795 0.465 ;
        RECT  2.690 0.185 2.765 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.185 1.045 ;
        RECT  3.095 0.185 3.115 0.465 ;
        RECT  3.095 0.745 3.115 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.980 0.375 ;
        RECT  2.450 -0.115 2.900 0.115 ;
        RECT  2.330 -0.115 2.450 0.275 ;
        RECT  1.810 -0.115 2.330 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 1.145 3.220 1.375 ;
        RECT  2.880 1.020 3.000 1.375 ;
        RECT  2.390 1.145 2.880 1.375 ;
        RECT  2.290 0.990 2.390 1.375 ;
        RECT  1.800 1.145 2.290 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.985 0.520 3.045 0.640 ;
        RECT  2.915 0.520 2.985 0.940 ;
        RECT  2.610 0.870 2.915 0.940 ;
        RECT  2.530 0.185 2.610 1.070 ;
        RECT  2.370 0.345 2.450 0.910 ;
        RECT  2.230 0.345 2.370 0.415 ;
        RECT  2.170 0.840 2.370 0.910 ;
        RECT  2.110 0.205 2.230 0.415 ;
        RECT  2.090 0.840 2.170 1.060 ;
        RECT  1.650 0.985 2.090 1.060 ;
        RECT  1.790 0.210 1.870 0.915 ;
        RECT  1.110 0.210 1.790 0.280 ;
        RECT  0.590 0.845 1.790 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDD1BWP

MACRO LNCSNDD2BWP
    CLASS CORE ;
    FOREIGN LNCSNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.105 0.640 ;
        RECT  1.995 0.495 2.065 0.780 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.690 0.185 2.770 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 0.355 3.185 0.905 ;
        RECT  3.115 0.185 3.130 1.055 ;
        RECT  3.050 0.185 3.115 0.465 ;
        RECT  3.050 0.735 3.115 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.960 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.350 1.670 0.485 ;
        RECT  0.665 0.350 1.590 0.420 ;
        RECT  0.595 0.350 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.115 3.360 0.115 ;
        RECT  3.235 -0.115 3.305 0.305 ;
        RECT  2.950 -0.115 3.235 0.115 ;
        RECT  2.870 -0.115 2.950 0.465 ;
        RECT  2.590 -0.115 2.870 0.115 ;
        RECT  2.510 -0.115 2.590 0.305 ;
        RECT  1.810 -0.115 2.510 0.115 ;
        RECT  1.680 -0.115 1.810 0.140 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.145 3.360 1.375 ;
        RECT  3.235 0.960 3.305 1.375 ;
        RECT  2.970 1.145 3.235 1.375 ;
        RECT  2.850 1.005 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.005 2.610 1.375 ;
        RECT  2.240 1.145 2.490 1.375 ;
        RECT  2.140 0.990 2.240 1.375 ;
        RECT  1.800 1.145 2.140 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.920 1.145 1.680 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.545 3.045 0.615 ;
        RECT  2.875 0.545 2.945 0.935 ;
        RECT  2.520 0.865 2.875 0.935 ;
        RECT  2.450 0.385 2.520 0.935 ;
        RECT  2.410 0.385 2.450 0.465 ;
        RECT  2.410 0.735 2.450 0.935 ;
        RECT  2.330 0.185 2.410 0.465 ;
        RECT  2.330 0.735 2.410 1.055 ;
        RECT  2.255 0.545 2.380 0.620 ;
        RECT  2.185 0.275 2.255 0.920 ;
        RECT  2.090 0.275 2.185 0.355 ;
        RECT  2.020 0.850 2.185 0.920 ;
        RECT  1.940 0.850 2.020 1.060 ;
        RECT  1.650 0.985 1.940 1.060 ;
        RECT  1.790 0.210 1.870 0.915 ;
        RECT  1.110 0.210 1.790 0.280 ;
        RECT  0.590 0.845 1.790 0.915 ;
        RECT  1.510 0.985 1.650 1.075 ;
        RECT  1.100 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.270 1.075 ;
        RECT  1.100 0.490 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.030 0.490 1.100 0.775 ;
        RECT  0.510 0.705 1.030 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDD2BWP

MACRO LNCSNDD4BWP
    CLASS CORE ;
    FOREIGN LNCSNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.705 3.410 0.795 ;
        RECT  3.315 0.185 3.385 0.485 ;
        RECT  3.255 0.355 3.315 0.485 ;
        RECT  3.045 0.355 3.255 0.795 ;
        RECT  3.025 0.355 3.045 0.485 ;
        RECT  2.930 0.705 3.045 0.795 ;
        RECT  2.955 0.185 3.025 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.105 0.465 ;
        RECT  4.095 0.775 4.105 1.055 ;
        RECT  4.035 0.185 4.095 1.055 ;
        RECT  3.885 0.355 4.035 0.905 ;
        RECT  3.745 0.355 3.885 0.465 ;
        RECT  3.745 0.775 3.885 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.775 3.745 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0250 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.645 0.485 ;
        RECT  0.665 0.345 1.575 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.485 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.570 -0.115 3.830 0.115 ;
        RECT  3.490 -0.115 3.570 0.465 ;
        RECT  3.230 -0.115 3.490 0.115 ;
        RECT  3.110 -0.115 3.230 0.275 ;
        RECT  2.850 -0.115 3.110 0.115 ;
        RECT  2.770 -0.115 2.850 0.305 ;
        RECT  2.500 -0.115 2.770 0.115 ;
        RECT  2.400 -0.115 2.500 0.275 ;
        RECT  1.780 -0.115 2.400 0.115 ;
        RECT  1.660 -0.115 1.780 0.135 ;
        RECT  0.680 -0.115 1.660 0.115 ;
        RECT  0.580 -0.115 0.680 0.270 ;
        RECT  0.310 -0.115 0.580 0.115 ;
        RECT  0.230 -0.115 0.310 0.280 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.665 4.290 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 0.985 3.950 1.375 ;
        RECT  3.590 1.145 3.830 1.375 ;
        RECT  3.470 1.005 3.590 1.375 ;
        RECT  3.230 1.145 3.470 1.375 ;
        RECT  3.110 1.005 3.230 1.375 ;
        RECT  2.870 1.145 3.110 1.375 ;
        RECT  2.750 1.005 2.870 1.375 ;
        RECT  2.510 1.145 2.750 1.375 ;
        RECT  2.390 0.995 2.510 1.375 ;
        RECT  2.150 1.145 2.390 1.375 ;
        RECT  2.030 0.995 2.150 1.375 ;
        RECT  0.910 1.145 2.030 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.355 3.815 0.465 ;
        RECT  3.745 0.775 3.815 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.775 3.745 1.055 ;
        RECT  3.325 0.705 3.410 0.795 ;
        RECT  3.325 0.185 3.385 0.485 ;
        RECT  2.955 0.185 2.975 0.485 ;
        RECT  2.930 0.705 2.975 0.795 ;
        RECT  3.565 0.540 3.795 0.620 ;
        RECT  3.495 0.540 3.565 0.935 ;
        RECT  2.850 0.865 3.495 0.935 ;
        RECT  2.780 0.385 2.850 0.935 ;
        RECT  2.670 0.385 2.780 0.465 ;
        RECT  2.665 0.865 2.780 0.935 ;
        RECT  2.590 0.185 2.670 0.465 ;
        RECT  2.595 0.735 2.665 1.055 ;
        RECT  2.515 0.545 2.660 0.615 ;
        RECT  2.445 0.345 2.515 0.925 ;
        RECT  2.150 0.345 2.445 0.415 ;
        RECT  1.950 0.855 2.445 0.925 ;
        RECT  2.300 0.500 2.375 0.775 ;
        RECT  1.820 0.705 2.300 0.775 ;
        RECT  2.030 0.205 2.150 0.415 ;
        RECT  1.870 0.855 1.950 1.055 ;
        RECT  1.670 0.985 1.870 1.055 ;
        RECT  1.795 0.520 1.820 0.775 ;
        RECT  1.725 0.205 1.795 0.915 ;
        RECT  1.090 0.205 1.725 0.275 ;
        RECT  0.590 0.845 1.725 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.510 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.180 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.410 0.260 0.490 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.245 0.350 0.410 0.420 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDD4BWP

MACRO LNCSNDQD1BWP
    CLASS CORE ;
    FOREIGN LNCSNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.495 2.065 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 0.355 2.765 0.905 ;
        RECT  2.695 0.185 2.730 1.055 ;
        RECT  2.650 0.185 2.695 0.465 ;
        RECT  2.650 0.735 2.695 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.345 1.660 0.485 ;
        RECT  0.665 0.345 1.580 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 -0.115 2.800 0.115 ;
        RECT  2.460 -0.115 2.540 0.315 ;
        RECT  1.800 -0.115 2.460 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 1.145 2.800 1.375 ;
        RECT  2.460 0.885 2.540 1.375 ;
        RECT  2.160 1.145 2.460 1.375 ;
        RECT  2.060 0.990 2.160 1.375 ;
        RECT  0.910 1.145 2.060 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.545 2.625 0.620 ;
        RECT  2.480 0.395 2.550 0.805 ;
        RECT  2.350 0.395 2.480 0.465 ;
        RECT  2.350 0.735 2.480 0.805 ;
        RECT  2.205 0.545 2.400 0.620 ;
        RECT  2.275 0.185 2.350 0.465 ;
        RECT  2.275 0.735 2.350 1.055 ;
        RECT  2.135 0.275 2.205 0.910 ;
        RECT  2.030 0.275 2.135 0.355 ;
        RECT  1.985 0.840 2.135 0.910 ;
        RECT  1.905 0.840 1.985 1.055 ;
        RECT  1.670 0.985 1.905 1.055 ;
        RECT  1.750 0.205 1.825 0.915 ;
        RECT  1.110 0.205 1.750 0.275 ;
        RECT  0.590 0.845 1.750 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.200 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDQD1BWP

MACRO LNCSNDQD2BWP
    CLASS CORE ;
    FOREIGN LNCSNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.495 2.065 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.710 0.355 2.765 0.905 ;
        RECT  2.695 0.185 2.710 1.055 ;
        RECT  2.630 0.185 2.695 0.465 ;
        RECT  2.630 0.735 2.695 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.345 1.660 0.485 ;
        RECT  0.665 0.345 1.580 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.815 -0.115 2.890 0.305 ;
        RECT  2.530 -0.115 2.815 0.115 ;
        RECT  2.450 -0.115 2.530 0.315 ;
        RECT  1.800 -0.115 2.450 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.985 2.900 1.375 ;
        RECT  2.530 1.145 2.800 1.375 ;
        RECT  2.450 0.885 2.530 1.375 ;
        RECT  2.160 1.145 2.450 1.375 ;
        RECT  2.060 0.990 2.160 1.375 ;
        RECT  0.910 1.145 2.060 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.550 0.545 2.625 0.620 ;
        RECT  2.480 0.395 2.550 0.805 ;
        RECT  2.350 0.395 2.480 0.465 ;
        RECT  2.350 0.735 2.480 0.805 ;
        RECT  2.205 0.545 2.400 0.620 ;
        RECT  2.275 0.185 2.350 0.465 ;
        RECT  2.275 0.735 2.350 1.055 ;
        RECT  2.170 0.335 2.205 0.910 ;
        RECT  2.135 0.200 2.170 0.910 ;
        RECT  2.050 0.200 2.135 0.415 ;
        RECT  1.985 0.840 2.135 0.910 ;
        RECT  1.905 0.840 1.985 1.055 ;
        RECT  1.670 0.985 1.905 1.055 ;
        RECT  1.750 0.205 1.825 0.915 ;
        RECT  1.110 0.205 1.750 0.275 ;
        RECT  0.590 0.845 1.750 0.915 ;
        RECT  1.540 0.985 1.670 1.075 ;
        RECT  1.085 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.200 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDQD2BWP

MACRO LNCSNDQD4BWP
    CLASS CORE ;
    FOREIGN LNCSNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.185 3.265 0.465 ;
        RECT  3.255 0.775 3.265 1.055 ;
        RECT  3.195 0.185 3.255 1.055 ;
        RECT  3.045 0.355 3.195 0.905 ;
        RECT  2.905 0.355 3.045 0.465 ;
        RECT  2.905 0.775 3.045 0.905 ;
        RECT  2.835 0.185 2.905 0.465 ;
        RECT  2.835 0.775 2.905 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0248 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0296 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.345 1.670 0.485 ;
        RECT  0.665 0.345 1.590 0.415 ;
        RECT  0.595 0.345 0.665 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.485 ;
        RECT  3.110 -0.115 3.370 0.115 ;
        RECT  2.990 -0.115 3.110 0.275 ;
        RECT  2.730 -0.115 2.990 0.115 ;
        RECT  2.650 -0.115 2.730 0.305 ;
        RECT  2.380 -0.115 2.650 0.115 ;
        RECT  2.280 -0.115 2.380 0.275 ;
        RECT  1.800 -0.115 2.280 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  0.700 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.700 0.270 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.665 3.450 1.375 ;
        RECT  3.110 1.145 3.370 1.375 ;
        RECT  2.990 0.985 3.110 1.375 ;
        RECT  2.730 1.145 2.990 1.375 ;
        RECT  2.650 0.925 2.730 1.375 ;
        RECT  2.370 1.145 2.650 1.375 ;
        RECT  2.290 0.925 2.370 1.375 ;
        RECT  2.190 1.145 2.290 1.375 ;
        RECT  2.110 0.925 2.190 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.140 1.800 1.375 ;
        RECT  0.910 1.145 1.680 1.375 ;
        RECT  0.780 1.125 0.910 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.355 2.975 0.465 ;
        RECT  2.905 0.775 2.975 0.905 ;
        RECT  2.835 0.185 2.905 0.465 ;
        RECT  2.835 0.775 2.905 1.055 ;
        RECT  2.750 0.545 2.850 0.615 ;
        RECT  2.680 0.385 2.750 0.805 ;
        RECT  2.550 0.385 2.680 0.465 ;
        RECT  2.550 0.735 2.680 0.805 ;
        RECT  2.345 0.545 2.590 0.620 ;
        RECT  2.470 0.185 2.550 0.465 ;
        RECT  2.470 0.735 2.550 1.055 ;
        RECT  2.275 0.345 2.345 0.845 ;
        RECT  2.190 0.345 2.275 0.415 ;
        RECT  2.000 0.775 2.275 0.845 ;
        RECT  2.070 0.205 2.190 0.415 ;
        RECT  1.920 0.775 2.000 1.055 ;
        RECT  1.650 0.985 1.920 1.055 ;
        RECT  1.760 0.205 1.840 0.915 ;
        RECT  1.110 0.205 1.760 0.275 ;
        RECT  0.590 0.845 1.760 0.915 ;
        RECT  1.530 0.985 1.650 1.075 ;
        RECT  1.085 0.705 1.530 0.775 ;
        RECT  1.110 0.985 1.230 1.075 ;
        RECT  1.085 0.495 1.200 0.570 ;
        RECT  0.125 0.985 1.110 1.055 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.510 0.705 1.015 0.775 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNCSNDQD4BWP

MACRO LNCSNQD1BWP
    CLASS CORE ;
    FOREIGN LNCSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.450 1.060 ;
        RECT  2.370 0.185 2.415 0.465 ;
        RECT  2.370 0.740 2.415 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.180 -0.115 2.260 0.315 ;
        RECT  1.530 -0.115 2.180 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.180 0.900 2.260 1.375 ;
        RECT  1.890 1.145 2.180 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.340 0.620 ;
        RECT  2.200 0.395 2.270 0.785 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.710 2.200 0.785 ;
        RECT  1.925 0.545 2.110 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.710 2.070 1.030 ;
        RECT  1.910 0.345 1.925 0.910 ;
        RECT  1.855 0.205 1.910 0.910 ;
        RECT  1.790 0.205 1.855 0.415 ;
        RECT  1.710 0.840 1.855 0.910 ;
        RECT  1.630 0.840 1.710 1.060 ;
        RECT  1.370 0.990 1.630 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.370 1.075 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCSNQD1BWP

MACRO LNCSNQD2BWP
    CLASS CORE ;
    FOREIGN LNCSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.060 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.740 2.415 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0270 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.290 ;
        RECT  2.250 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.530 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.145 2.660 1.375 ;
        RECT  2.520 0.985 2.620 1.375 ;
        RECT  2.250 1.145 2.520 1.375 ;
        RECT  2.170 0.900 2.250 1.375 ;
        RECT  1.890 1.145 2.170 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.340 0.620 ;
        RECT  2.200 0.395 2.270 0.785 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.710 2.200 0.785 ;
        RECT  1.925 0.545 2.120 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.710 2.070 1.030 ;
        RECT  1.910 0.345 1.925 0.910 ;
        RECT  1.855 0.200 1.910 0.910 ;
        RECT  1.790 0.200 1.855 0.415 ;
        RECT  1.710 0.840 1.855 0.910 ;
        RECT  1.630 0.840 1.710 1.060 ;
        RECT  1.390 0.990 1.630 1.060 ;
        RECT  1.550 0.520 1.575 0.640 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.390 1.070 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.290 0.120 0.555 ;
        RECT  0.035 0.290 0.105 1.075 ;
    END
END LNCSNQD2BWP

MACRO LNCSNQD4BWP
    CLASS CORE ;
    FOREIGN LNCSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.185 2.990 0.485 ;
        RECT  2.910 0.760 2.990 1.040 ;
        RECT  2.835 0.355 2.910 0.485 ;
        RECT  2.835 0.760 2.910 0.905 ;
        RECT  2.630 0.355 2.835 0.905 ;
        RECT  2.625 0.355 2.630 1.040 ;
        RECT  2.540 0.185 2.625 0.480 ;
        RECT  2.540 0.760 2.625 1.040 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0374 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.990 1.010 1.075 ;
        RECT  0.285 0.990 0.850 1.060 ;
        RECT  0.245 0.840 0.285 1.060 ;
        RECT  0.215 0.635 0.245 1.060 ;
        RECT  0.175 0.635 0.215 0.910 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.525 0.665 0.595 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.390 0.485 ;
        RECT  1.090 0.350 1.295 0.420 ;
        RECT  1.015 0.350 1.090 0.625 ;
        RECT  0.750 0.350 1.015 0.420 ;
        RECT  0.680 0.205 0.750 0.420 ;
        RECT  0.460 0.205 0.680 0.275 ;
        RECT  0.340 0.185 0.460 0.275 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.485 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.280 ;
        RECT  2.440 -0.115 2.710 0.115 ;
        RECT  2.360 -0.115 2.440 0.465 ;
        RECT  2.090 -0.115 2.360 0.115 ;
        RECT  1.970 -0.115 2.090 0.275 ;
        RECT  1.530 -0.115 1.970 0.115 ;
        RECT  1.400 -0.115 1.530 0.140 ;
        RECT  0.260 -0.115 1.400 0.115 ;
        RECT  0.260 0.345 0.375 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.665 3.170 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.005 2.830 1.375 ;
        RECT  2.440 1.145 2.710 1.375 ;
        RECT  2.360 0.740 2.440 1.375 ;
        RECT  2.070 1.145 2.360 1.375 ;
        RECT  1.990 0.980 2.070 1.375 ;
        RECT  1.890 1.145 1.990 1.375 ;
        RECT  1.810 0.980 1.890 1.375 ;
        RECT  1.520 1.145 1.810 1.375 ;
        RECT  1.400 1.140 1.520 1.375 ;
        RECT  0.720 1.145 1.400 1.375 ;
        RECT  0.600 1.130 0.720 1.375 ;
        RECT  0.360 1.145 0.600 1.375 ;
        RECT  0.240 1.130 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.910 0.185 2.990 0.485 ;
        RECT  2.910 0.760 2.990 1.040 ;
        RECT  2.905 0.355 2.910 0.485 ;
        RECT  2.905 0.760 2.910 0.905 ;
        RECT  2.540 0.185 2.555 0.480 ;
        RECT  2.540 0.760 2.555 1.040 ;
        RECT  2.250 0.550 2.530 0.620 ;
        RECT  2.170 0.185 2.250 1.045 ;
        RECT  2.010 0.355 2.090 0.910 ;
        RECT  1.770 0.355 2.010 0.425 ;
        RECT  1.730 0.840 2.010 0.910 ;
        RECT  1.660 0.840 1.730 1.060 ;
        RECT  1.390 0.990 1.660 1.060 ;
        RECT  1.480 0.210 1.550 0.920 ;
        RECT  0.830 0.210 1.480 0.280 ;
        RECT  0.370 0.850 1.480 0.920 ;
        RECT  1.230 0.990 1.390 1.070 ;
        RECT  0.815 0.705 1.250 0.775 ;
        RECT  0.815 0.490 0.945 0.580 ;
        RECT  0.745 0.490 0.815 0.775 ;
        RECT  0.385 0.705 0.745 0.775 ;
        RECT  0.315 0.485 0.385 0.775 ;
        RECT  0.120 0.485 0.315 0.555 ;
        RECT  0.105 0.975 0.145 1.075 ;
        RECT  0.105 0.200 0.120 0.555 ;
        RECT  0.035 0.200 0.105 1.075 ;
    END
END LNCSNQD4BWP

MACRO LND1BWP
    CLASS CORE ;
    FOREIGN LND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.185 2.205 1.045 ;
        RECT  2.110 0.185 2.135 0.465 ;
        RECT  2.110 0.725 2.135 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.350 1.805 0.905 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.355 0.670 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 -0.115 2.240 0.115 ;
        RECT  1.900 -0.115 2.020 0.135 ;
        RECT  1.440 -0.115 1.900 0.115 ;
        RECT  1.360 -0.115 1.440 0.300 ;
        RECT  0.360 -0.115 1.360 0.115 ;
        RECT  0.240 -0.115 0.360 0.135 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 1.145 2.240 1.375 ;
        RECT  1.900 1.120 2.020 1.375 ;
        RECT  1.470 1.145 1.900 1.375 ;
        RECT  1.350 0.860 1.470 1.375 ;
        RECT  0.700 1.145 1.350 1.375 ;
        RECT  0.630 0.750 0.700 1.375 ;
        RECT  0.590 0.750 0.630 0.870 ;
        RECT  0.360 1.145 0.630 1.375 ;
        RECT  0.240 1.110 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.990 0.520 2.060 0.640 ;
        RECT  1.920 0.205 1.990 1.050 ;
        RECT  1.630 0.205 1.920 0.275 ;
        RECT  1.630 0.980 1.920 1.050 ;
        RECT  1.550 0.205 1.630 0.465 ;
        RECT  1.480 0.545 1.630 0.620 ;
        RECT  1.550 0.730 1.630 1.050 ;
        RECT  1.310 0.395 1.550 0.465 ;
        RECT  1.410 0.545 1.480 0.790 ;
        RECT  1.140 0.720 1.410 0.790 ;
        RECT  1.240 0.395 1.310 0.640 ;
        RECT  1.020 0.985 1.180 1.075 ;
        RECT  1.070 0.195 1.140 0.905 ;
        RECT  0.930 0.195 1.070 0.275 ;
        RECT  0.930 0.835 1.070 0.905 ;
        RECT  0.850 0.985 1.020 1.055 ;
        RECT  0.850 0.395 1.000 0.465 ;
        RECT  0.780 0.205 0.850 1.055 ;
        RECT  0.330 0.205 0.780 0.275 ;
        RECT  0.510 0.950 0.555 1.070 ;
        RECT  0.440 0.350 0.510 1.070 ;
        RECT  0.400 0.350 0.440 0.450 ;
        RECT  0.400 0.735 0.440 0.845 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.205 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.125 0.850 0.260 0.920 ;
        RECT  0.055 0.850 0.125 1.020 ;
    END
END LND1BWP

MACRO LND2BWP
    CLASS CORE ;
    FOREIGN LND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.355 2.345 0.905 ;
        RECT  2.275 0.185 2.290 1.030 ;
        RECT  2.210 0.185 2.275 0.465 ;
        RECT  2.210 0.730 2.275 1.030 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.195 1.925 0.780 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0164 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.355 0.670 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.295 ;
        RECT  2.110 -0.115 2.390 0.115 ;
        RECT  2.030 -0.115 2.110 0.460 ;
        RECT  1.750 -0.115 2.030 0.115 ;
        RECT  1.670 -0.115 1.750 0.315 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.315 ;
        RECT  0.360 -0.115 1.310 0.115 ;
        RECT  0.240 -0.115 0.360 0.135 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.975 2.470 1.375 ;
        RECT  2.120 1.145 2.390 1.375 ;
        RECT  2.020 0.990 2.120 1.375 ;
        RECT  1.765 1.145 2.020 1.375 ;
        RECT  1.655 0.990 1.765 1.375 ;
        RECT  1.405 1.145 1.655 1.375 ;
        RECT  1.300 0.860 1.405 1.375 ;
        RECT  0.700 1.145 1.300 1.375 ;
        RECT  0.630 0.750 0.700 1.375 ;
        RECT  0.590 0.750 0.630 0.870 ;
        RECT  0.360 1.145 0.630 1.375 ;
        RECT  0.240 1.110 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.090 0.545 2.200 0.620 ;
        RECT  2.020 0.545 2.090 0.920 ;
        RECT  1.730 0.850 2.020 0.920 ;
        RECT  1.660 0.395 1.730 0.920 ;
        RECT  1.570 0.395 1.660 0.465 ;
        RECT  1.570 0.850 1.660 0.920 ;
        RECT  1.420 0.545 1.580 0.615 ;
        RECT  1.490 0.185 1.570 0.465 ;
        RECT  1.490 0.720 1.570 1.040 ;
        RECT  1.280 0.395 1.490 0.465 ;
        RECT  1.350 0.545 1.420 0.790 ;
        RECT  1.120 0.720 1.350 0.790 ;
        RECT  1.200 0.395 1.280 0.640 ;
        RECT  1.000 0.985 1.160 1.075 ;
        RECT  1.050 0.195 1.120 0.915 ;
        RECT  0.910 0.195 1.050 0.275 ;
        RECT  0.930 0.835 1.050 0.915 ;
        RECT  0.840 0.985 1.000 1.055 ;
        RECT  0.840 0.380 0.980 0.460 ;
        RECT  0.770 0.205 0.840 1.055 ;
        RECT  0.330 0.205 0.770 0.275 ;
        RECT  0.510 0.950 0.555 1.070 ;
        RECT  0.440 0.350 0.510 1.070 ;
        RECT  0.400 0.350 0.440 0.450 ;
        RECT  0.400 0.735 0.440 0.845 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.205 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.125 0.850 0.260 0.920 ;
        RECT  0.055 0.850 0.125 1.020 ;
    END
END LND2BWP

MACRO LND4BWP
    CLASS CORE ;
    FOREIGN LND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.775 3.125 1.055 ;
        RECT  3.055 0.185 3.115 1.055 ;
        RECT  2.905 0.355 3.055 0.905 ;
        RECT  2.765 0.355 2.905 0.465 ;
        RECT  2.765 0.775 2.905 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.705 2.430 0.795 ;
        RECT  2.335 0.185 2.405 0.485 ;
        RECT  2.275 0.355 2.335 0.485 ;
        RECT  2.065 0.355 2.275 0.795 ;
        RECT  2.045 0.355 2.065 0.485 ;
        RECT  1.950 0.705 2.065 0.795 ;
        RECT  1.975 0.185 2.045 0.485 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0156 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.680 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.485 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.275 ;
        RECT  2.590 -0.115 2.850 0.115 ;
        RECT  2.510 -0.115 2.590 0.465 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.275 ;
        RECT  1.865 -0.115 2.130 0.115 ;
        RECT  1.795 -0.115 1.865 0.310 ;
        RECT  1.460 -0.115 1.795 0.115 ;
        RECT  1.380 -0.115 1.460 0.300 ;
        RECT  0.720 -0.115 1.380 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.140 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.665 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.985 2.970 1.375 ;
        RECT  2.610 1.145 2.850 1.375 ;
        RECT  2.490 1.005 2.610 1.375 ;
        RECT  2.250 1.145 2.490 1.375 ;
        RECT  2.130 1.005 2.250 1.375 ;
        RECT  1.890 1.145 2.130 1.375 ;
        RECT  1.770 1.005 1.890 1.375 ;
        RECT  1.470 1.145 1.770 1.375 ;
        RECT  1.370 0.850 1.470 1.375 ;
        RECT  0.730 1.145 1.370 1.375 ;
        RECT  0.660 0.740 0.730 1.375 ;
        RECT  0.630 0.740 0.660 0.860 ;
        RECT  0.330 1.145 0.660 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.465 ;
        RECT  2.765 0.775 2.835 0.905 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.775 2.765 1.055 ;
        RECT  2.345 0.705 2.430 0.795 ;
        RECT  2.345 0.185 2.405 0.485 ;
        RECT  1.975 0.185 1.995 0.485 ;
        RECT  1.950 0.705 1.995 0.795 ;
        RECT  2.585 0.540 2.815 0.620 ;
        RECT  2.515 0.540 2.585 0.935 ;
        RECT  1.860 0.865 2.515 0.935 ;
        RECT  1.790 0.395 1.860 0.935 ;
        RECT  1.650 0.395 1.790 0.465 ;
        RECT  1.650 0.865 1.790 0.935 ;
        RECT  1.490 0.545 1.710 0.620 ;
        RECT  1.570 0.185 1.650 0.465 ;
        RECT  1.570 0.720 1.650 1.040 ;
        RECT  1.340 0.395 1.570 0.465 ;
        RECT  1.420 0.545 1.490 0.780 ;
        RECT  1.170 0.710 1.420 0.780 ;
        RECT  1.260 0.395 1.340 0.640 ;
        RECT  1.040 0.995 1.200 1.075 ;
        RECT  1.100 0.195 1.170 0.915 ;
        RECT  0.950 0.195 1.100 0.275 ;
        RECT  0.950 0.835 1.100 0.915 ;
        RECT  0.870 0.995 1.040 1.065 ;
        RECT  0.870 0.360 1.020 0.440 ;
        RECT  0.800 0.210 0.870 1.065 ;
        RECT  0.340 0.210 0.800 0.280 ;
        RECT  0.520 0.955 0.590 1.075 ;
        RECT  0.450 0.350 0.520 1.075 ;
        RECT  0.420 0.350 0.450 0.450 ;
        RECT  0.410 0.710 0.450 0.850 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.210 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.020 ;
    END
END LND4BWP

MACRO LNQD1BWP
    CLASS CORE ;
    FOREIGN LNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.185 2.065 1.070 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.355 0.670 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 -0.115 2.100 0.115 ;
        RECT  1.790 -0.115 1.870 0.485 ;
        RECT  1.460 -0.115 1.790 0.115 ;
        RECT  1.380 -0.115 1.460 0.310 ;
        RECT  0.360 -0.115 1.380 0.115 ;
        RECT  0.240 -0.115 0.360 0.135 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.145 2.100 1.375 ;
        RECT  1.790 0.665 1.870 1.375 ;
        RECT  1.480 1.145 1.790 1.375 ;
        RECT  1.360 0.860 1.480 1.375 ;
        RECT  0.700 1.145 1.360 1.375 ;
        RECT  0.630 0.750 0.700 1.375 ;
        RECT  0.590 0.750 0.630 0.870 ;
        RECT  0.360 1.145 0.630 1.375 ;
        RECT  0.240 1.110 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.595 0.190 1.670 0.975 ;
        RECT  1.590 0.190 1.595 0.460 ;
        RECT  1.320 0.390 1.590 0.460 ;
        RECT  1.425 0.530 1.525 0.790 ;
        RECT  1.140 0.720 1.425 0.790 ;
        RECT  1.240 0.390 1.320 0.640 ;
        RECT  1.020 0.985 1.180 1.075 ;
        RECT  1.070 0.195 1.140 0.905 ;
        RECT  0.930 0.195 1.070 0.275 ;
        RECT  0.930 0.835 1.070 0.905 ;
        RECT  0.850 0.985 1.020 1.055 ;
        RECT  0.850 0.395 1.000 0.465 ;
        RECT  0.780 0.205 0.850 1.055 ;
        RECT  0.330 0.205 0.780 0.275 ;
        RECT  0.510 0.950 0.555 1.070 ;
        RECT  0.440 0.350 0.510 1.070 ;
        RECT  0.400 0.350 0.440 0.450 ;
        RECT  0.400 0.735 0.440 0.845 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.205 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.125 0.850 0.260 0.920 ;
        RECT  0.055 0.850 0.125 1.020 ;
    END
END LNQD1BWP

MACRO LNQD2BWP
    CLASS CORE ;
    FOREIGN LNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.195 1.925 1.070 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.355 0.670 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.115 2.240 0.115 ;
        RECT  2.050 -0.115 2.140 0.460 ;
        RECT  1.750 -0.115 2.050 0.115 ;
        RECT  1.670 -0.115 1.750 0.315 ;
        RECT  1.390 -0.115 1.670 0.115 ;
        RECT  1.310 -0.115 1.390 0.315 ;
        RECT  0.360 -0.115 1.310 0.115 ;
        RECT  0.240 -0.115 0.360 0.135 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.145 2.240 1.375 ;
        RECT  2.050 0.665 2.140 1.375 ;
        RECT  1.760 1.145 2.050 1.375 ;
        RECT  1.660 0.990 1.760 1.375 ;
        RECT  1.400 1.145 1.660 1.375 ;
        RECT  1.300 0.860 1.400 1.375 ;
        RECT  0.700 1.145 1.300 1.375 ;
        RECT  0.630 0.750 0.700 1.375 ;
        RECT  0.590 0.750 0.630 0.870 ;
        RECT  0.360 1.145 0.630 1.375 ;
        RECT  0.240 1.110 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.660 0.395 1.730 0.920 ;
        RECT  1.570 0.395 1.660 0.465 ;
        RECT  1.470 0.850 1.660 0.920 ;
        RECT  1.420 0.545 1.580 0.615 ;
        RECT  1.490 0.185 1.570 0.465 ;
        RECT  1.280 0.395 1.490 0.465 ;
        RECT  1.350 0.545 1.420 0.790 ;
        RECT  1.120 0.720 1.350 0.790 ;
        RECT  1.200 0.395 1.280 0.640 ;
        RECT  1.000 0.985 1.160 1.075 ;
        RECT  1.050 0.205 1.120 0.915 ;
        RECT  0.910 0.205 1.050 0.285 ;
        RECT  0.930 0.835 1.050 0.915 ;
        RECT  0.840 0.985 1.000 1.055 ;
        RECT  0.840 0.380 0.980 0.460 ;
        RECT  0.770 0.205 0.840 1.055 ;
        RECT  0.330 0.205 0.770 0.275 ;
        RECT  0.510 0.950 0.555 1.070 ;
        RECT  0.440 0.350 0.510 1.070 ;
        RECT  0.400 0.350 0.440 0.450 ;
        RECT  0.400 0.735 0.440 0.845 ;
        RECT  0.330 0.520 0.370 0.640 ;
        RECT  0.260 0.205 0.330 0.920 ;
        RECT  0.055 0.260 0.260 0.380 ;
        RECT  0.125 0.850 0.260 0.920 ;
        RECT  0.055 0.850 0.125 1.020 ;
    END
END LNQD2BWP

MACRO LNQD4BWP
    CLASS CORE ;
    FOREIGN LNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.275 0.355 2.350 0.485 ;
        RECT  2.275 0.760 2.350 0.905 ;
        RECT  2.070 0.355 2.275 0.905 ;
        RECT  2.065 0.185 2.070 1.045 ;
        RECT  1.995 0.185 2.065 0.485 ;
        RECT  1.995 0.760 2.065 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.355 0.680 0.660 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.485 ;
        RECT  2.260 -0.115 2.530 0.115 ;
        RECT  2.160 -0.115 2.260 0.275 ;
        RECT  1.890 -0.115 2.160 0.115 ;
        RECT  1.815 -0.115 1.890 0.485 ;
        RECT  1.480 -0.115 1.815 0.115 ;
        RECT  1.400 -0.115 1.480 0.315 ;
        RECT  0.720 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.140 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.665 2.610 1.375 ;
        RECT  2.260 1.145 2.530 1.375 ;
        RECT  2.160 0.985 2.260 1.375 ;
        RECT  1.890 1.145 2.160 1.375 ;
        RECT  1.815 0.685 1.890 1.375 ;
        RECT  1.490 1.145 1.815 1.375 ;
        RECT  1.390 0.850 1.490 1.375 ;
        RECT  0.730 1.145 1.390 1.375 ;
        RECT  0.660 0.740 0.730 1.375 ;
        RECT  0.630 0.740 0.660 0.860 ;
        RECT  0.330 1.145 0.660 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.345 0.355 2.350 0.485 ;
        RECT  2.345 0.760 2.350 0.905 ;
        RECT  1.690 0.395 1.745 0.930 ;
        RECT  1.675 0.185 1.690 0.930 ;
        RECT  1.610 0.185 1.675 0.465 ;
        RECT  1.570 0.850 1.675 0.930 ;
        RECT  1.340 0.395 1.610 0.465 ;
        RECT  1.500 0.545 1.580 0.780 ;
        RECT  1.170 0.710 1.500 0.780 ;
        RECT  1.260 0.395 1.340 0.640 ;
        RECT  1.040 0.995 1.200 1.075 ;
        RECT  1.100 0.195 1.170 0.915 ;
        RECT  0.950 0.195 1.100 0.275 ;
        RECT  0.950 0.835 1.100 0.915 ;
        RECT  0.870 0.995 1.040 1.065 ;
        RECT  0.870 0.360 1.020 0.440 ;
        RECT  0.800 0.210 0.870 1.065 ;
        RECT  0.340 0.210 0.800 0.280 ;
        RECT  0.520 0.955 0.590 1.075 ;
        RECT  0.450 0.350 0.520 1.075 ;
        RECT  0.420 0.350 0.450 0.450 ;
        RECT  0.410 0.710 0.450 0.850 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.210 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.020 ;
    END
END LNQD4BWP

MACRO LNSND1BWP
    CLASS CORE ;
    FOREIGN LNSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.390 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.720 1.990 0.790 ;
        RECT  1.925 0.185 1.955 0.465 ;
        RECT  1.850 0.185 1.925 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.345 1.045 ;
        RECT  2.255 0.185 2.275 0.465 ;
        RECT  2.255 0.745 2.275 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 0.985 0.600 1.075 ;
        RECT  0.275 0.985 0.470 1.055 ;
        RECT  0.245 0.825 0.275 1.055 ;
        RECT  0.205 0.495 0.245 1.055 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.115 2.380 0.115 ;
        RECT  2.060 -0.115 2.140 0.375 ;
        RECT  1.610 -0.115 2.060 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  1.050 -0.115 1.490 0.115 ;
        RECT  0.970 -0.115 1.050 0.430 ;
        RECT  0.315 -0.115 0.970 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.145 2.380 1.375 ;
        RECT  2.040 1.020 2.160 1.375 ;
        RECT  1.550 1.145 2.040 1.375 ;
        RECT  1.450 0.990 1.550 1.375 ;
        RECT  0.340 1.145 1.450 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.145 0.520 2.205 0.640 ;
        RECT  2.075 0.520 2.145 0.940 ;
        RECT  1.770 0.870 2.075 0.940 ;
        RECT  1.690 0.185 1.770 1.045 ;
        RECT  1.530 0.345 1.610 0.910 ;
        RECT  1.290 0.345 1.530 0.415 ;
        RECT  1.300 0.840 1.530 0.910 ;
        RECT  1.220 0.840 1.300 1.060 ;
        RECT  0.850 0.985 1.220 1.060 ;
        RECT  1.000 0.520 1.160 0.640 ;
        RECT  0.930 0.520 1.000 0.910 ;
        RECT  0.815 0.520 0.930 0.590 ;
        RECT  0.710 0.840 0.930 0.910 ;
        RECT  0.665 0.695 0.850 0.765 ;
        RECT  0.745 0.195 0.815 0.590 ;
        RECT  0.730 0.195 0.745 0.265 ;
        RECT  0.570 0.185 0.730 0.265 ;
        RECT  0.570 0.840 0.710 0.915 ;
        RECT  0.595 0.345 0.665 0.765 ;
        RECT  0.130 0.345 0.595 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSND1BWP

MACRO LNSND2BWP
    CLASS CORE ;
    FOREIGN LNSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.365 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.065 0.800 ;
        RECT  1.960 0.185 1.995 0.465 ;
        RECT  1.925 0.730 1.995 0.800 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.050 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.730 2.415 1.050 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.980 0.610 1.075 ;
        RECT  0.275 0.980 0.480 1.050 ;
        RECT  0.245 0.825 0.275 1.050 ;
        RECT  0.205 0.495 0.245 1.050 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.290 ;
        RECT  2.240 -0.115 2.520 0.115 ;
        RECT  2.160 -0.115 2.240 0.465 ;
        RECT  1.845 -0.115 2.160 0.115 ;
        RECT  1.770 -0.115 1.845 0.465 ;
        RECT  1.090 -0.115 1.770 0.115 ;
        RECT  1.010 -0.115 1.090 0.420 ;
        RECT  0.315 -0.115 1.010 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.145 2.660 1.375 ;
        RECT  2.520 0.985 2.620 1.375 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.140 1.025 2.260 1.375 ;
        RECT  1.870 1.145 2.140 1.375 ;
        RECT  1.750 1.020 1.870 1.375 ;
        RECT  1.500 1.145 1.750 1.375 ;
        RECT  1.380 1.000 1.500 1.375 ;
        RECT  0.340 1.145 1.380 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.265 0.545 2.345 0.620 ;
        RECT  2.185 0.545 2.265 0.940 ;
        RECT  1.700 0.870 2.185 0.940 ;
        RECT  1.670 0.205 1.700 0.940 ;
        RECT  1.630 0.205 1.670 1.020 ;
        RECT  1.530 0.205 1.630 0.275 ;
        RECT  1.590 0.700 1.630 1.020 ;
        RECT  1.520 0.520 1.550 0.640 ;
        RECT  1.450 0.345 1.520 0.915 ;
        RECT  1.350 0.345 1.450 0.415 ;
        RECT  1.280 0.845 1.450 0.915 ;
        RECT  1.200 0.845 1.280 1.055 ;
        RECT  1.000 0.540 1.200 0.620 ;
        RECT  0.850 0.980 1.200 1.055 ;
        RECT  0.930 0.540 1.000 0.900 ;
        RECT  0.815 0.540 0.930 0.610 ;
        RECT  0.570 0.830 0.930 0.900 ;
        RECT  0.665 0.680 0.850 0.755 ;
        RECT  0.745 0.185 0.815 0.610 ;
        RECT  0.600 0.185 0.745 0.265 ;
        RECT  0.595 0.345 0.665 0.755 ;
        RECT  0.130 0.345 0.595 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSND2BWP

MACRO LNSND4BWP
    CLASS CORE ;
    FOREIGN LNSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.630 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.705 2.710 0.795 ;
        RECT  2.615 0.185 2.685 0.485 ;
        RECT  2.555 0.355 2.615 0.485 ;
        RECT  2.345 0.355 2.555 0.795 ;
        RECT  2.325 0.355 2.345 0.485 ;
        RECT  2.230 0.705 2.345 0.795 ;
        RECT  2.255 0.185 2.325 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.185 3.405 0.465 ;
        RECT  3.395 0.775 3.405 1.055 ;
        RECT  3.335 0.185 3.395 1.055 ;
        RECT  3.185 0.355 3.335 0.905 ;
        RECT  3.045 0.355 3.185 0.465 ;
        RECT  3.045 0.775 3.185 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.980 0.610 1.075 ;
        RECT  0.275 0.980 0.480 1.050 ;
        RECT  0.245 0.825 0.275 1.050 ;
        RECT  0.205 0.495 0.245 1.050 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.640 0.115 ;
        RECT  3.510 -0.115 3.590 0.485 ;
        RECT  3.250 -0.115 3.510 0.115 ;
        RECT  3.130 -0.115 3.250 0.275 ;
        RECT  2.870 -0.115 3.130 0.115 ;
        RECT  2.790 -0.115 2.870 0.465 ;
        RECT  2.530 -0.115 2.790 0.115 ;
        RECT  2.410 -0.115 2.530 0.275 ;
        RECT  2.150 -0.115 2.410 0.115 ;
        RECT  2.070 -0.115 2.150 0.315 ;
        RECT  1.810 -0.115 2.070 0.115 ;
        RECT  1.690 -0.115 1.810 0.265 ;
        RECT  1.070 -0.115 1.690 0.115 ;
        RECT  0.990 -0.115 1.070 0.430 ;
        RECT  0.315 -0.115 0.990 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.665 3.590 1.375 ;
        RECT  3.250 1.145 3.510 1.375 ;
        RECT  3.130 0.985 3.250 1.375 ;
        RECT  2.890 1.145 3.130 1.375 ;
        RECT  2.770 1.005 2.890 1.375 ;
        RECT  2.530 1.145 2.770 1.375 ;
        RECT  2.410 1.005 2.530 1.375 ;
        RECT  2.170 1.145 2.410 1.375 ;
        RECT  2.050 1.005 2.170 1.375 ;
        RECT  1.810 1.145 2.050 1.375 ;
        RECT  1.690 1.010 1.810 1.375 ;
        RECT  1.450 1.145 1.690 1.375 ;
        RECT  1.330 1.010 1.450 1.375 ;
        RECT  0.340 1.145 1.330 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.355 3.115 0.465 ;
        RECT  3.045 0.775 3.115 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        RECT  2.625 0.705 2.710 0.795 ;
        RECT  2.625 0.185 2.685 0.485 ;
        RECT  2.255 0.185 2.275 0.485 ;
        RECT  2.230 0.705 2.275 0.795 ;
        RECT  2.865 0.540 3.095 0.620 ;
        RECT  2.795 0.540 2.865 0.935 ;
        RECT  2.160 0.865 2.795 0.935 ;
        RECT  2.090 0.395 2.160 0.935 ;
        RECT  1.970 0.395 2.090 0.465 ;
        RECT  1.970 0.865 2.090 0.935 ;
        RECT  1.820 0.545 2.010 0.620 ;
        RECT  1.890 0.185 1.970 0.465 ;
        RECT  1.890 0.740 1.970 1.060 ;
        RECT  1.750 0.345 1.820 0.940 ;
        RECT  1.450 0.345 1.750 0.415 ;
        RECT  1.250 0.870 1.750 0.940 ;
        RECT  1.600 0.500 1.680 0.800 ;
        RECT  1.180 0.730 1.600 0.800 ;
        RECT  1.330 0.205 1.450 0.415 ;
        RECT  1.170 0.870 1.250 1.055 ;
        RECT  1.100 0.500 1.180 0.800 ;
        RECT  0.830 0.980 1.170 1.055 ;
        RECT  0.815 0.500 1.100 0.570 ;
        RECT  1.000 0.730 1.100 0.800 ;
        RECT  0.930 0.730 1.000 0.900 ;
        RECT  0.570 0.830 0.930 0.900 ;
        RECT  0.665 0.675 0.850 0.755 ;
        RECT  0.745 0.185 0.815 0.570 ;
        RECT  0.590 0.185 0.745 0.265 ;
        RECT  0.595 0.345 0.665 0.755 ;
        RECT  0.130 0.345 0.595 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSND4BWP

MACRO LNSNDD1BWP
    CLASS CORE ;
    FOREIGN LNSNDD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.720 2.410 0.790 ;
        RECT  2.345 0.185 2.375 0.465 ;
        RECT  2.270 0.185 2.345 0.790 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.765 1.045 ;
        RECT  2.675 0.185 2.695 0.465 ;
        RECT  2.675 0.745 2.695 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 -0.115 2.800 0.115 ;
        RECT  2.480 -0.115 2.560 0.375 ;
        RECT  2.030 -0.115 2.480 0.115 ;
        RECT  1.910 -0.115 2.030 0.275 ;
        RECT  1.480 -0.115 1.910 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  0.700 -0.115 1.360 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.145 2.800 1.375 ;
        RECT  2.460 1.020 2.580 1.375 ;
        RECT  1.970 1.145 2.460 1.375 ;
        RECT  1.870 0.990 1.970 1.375 ;
        RECT  0.730 1.145 1.870 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.565 0.520 2.625 0.640 ;
        RECT  2.495 0.520 2.565 0.940 ;
        RECT  2.190 0.870 2.495 0.940 ;
        RECT  2.110 0.185 2.190 1.070 ;
        RECT  1.950 0.345 2.030 0.910 ;
        RECT  1.710 0.345 1.950 0.415 ;
        RECT  1.730 0.840 1.950 0.910 ;
        RECT  1.650 0.840 1.730 1.055 ;
        RECT  1.420 0.985 1.650 1.055 ;
        RECT  1.500 0.205 1.580 0.915 ;
        RECT  0.960 0.205 1.500 0.275 ;
        RECT  0.960 0.845 1.500 0.915 ;
        RECT  1.280 0.985 1.420 1.075 ;
        RECT  1.020 0.700 1.260 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.850 0.985 0.970 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.125 0.985 0.850 1.055 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDD1BWP

MACRO LNSNDD2BWP
    CLASS CORE ;
    FOREIGN LNSNDD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 1.835 0.640 ;
        RECT  1.715 0.495 1.785 0.780 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 0.795 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.355 2.905 0.905 ;
        RECT  2.835 0.185 2.850 1.055 ;
        RECT  2.770 0.185 2.835 0.465 ;
        RECT  2.770 0.735 2.835 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.115 3.080 0.115 ;
        RECT  2.955 -0.115 3.025 0.305 ;
        RECT  2.670 -0.115 2.955 0.115 ;
        RECT  2.590 -0.115 2.670 0.465 ;
        RECT  2.310 -0.115 2.590 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.520 -0.115 2.230 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.145 3.080 1.375 ;
        RECT  2.940 0.985 3.040 1.375 ;
        RECT  2.690 1.145 2.940 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  1.960 1.145 2.210 1.375 ;
        RECT  1.860 0.990 1.960 1.375 ;
        RECT  0.730 1.145 1.860 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.665 0.545 2.765 0.620 ;
        RECT  2.595 0.545 2.665 0.935 ;
        RECT  2.335 0.865 2.595 0.935 ;
        RECT  2.265 0.385 2.335 0.935 ;
        RECT  2.130 0.385 2.265 0.465 ;
        RECT  2.130 0.865 2.265 0.935 ;
        RECT  1.975 0.545 2.185 0.620 ;
        RECT  2.055 0.185 2.130 0.465 ;
        RECT  2.050 0.735 2.130 1.055 ;
        RECT  1.905 0.245 1.975 0.920 ;
        RECT  1.850 0.245 1.905 0.315 ;
        RECT  1.760 0.850 1.905 0.920 ;
        RECT  1.680 0.850 1.760 1.055 ;
        RECT  1.420 0.985 1.680 1.055 ;
        RECT  1.520 0.205 1.600 0.915 ;
        RECT  0.960 0.205 1.520 0.275 ;
        RECT  0.930 0.845 1.520 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.125 0.985 0.820 1.055 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDD2BWP

MACRO LNSNDD4BWP
    CLASS CORE ;
    FOREIGN LNSNDD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.545 1.870 0.625 ;
        RECT  1.715 0.355 1.785 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.705 3.130 0.795 ;
        RECT  3.035 0.185 3.105 0.485 ;
        RECT  2.975 0.355 3.035 0.485 ;
        RECT  2.765 0.355 2.975 0.795 ;
        RECT  2.745 0.355 2.765 0.485 ;
        RECT  2.650 0.705 2.765 0.795 ;
        RECT  2.675 0.185 2.745 0.485 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.825 0.465 ;
        RECT  3.815 0.775 3.825 1.055 ;
        RECT  3.755 0.185 3.815 1.055 ;
        RECT  3.605 0.355 3.755 0.905 ;
        RECT  3.465 0.355 3.605 0.465 ;
        RECT  3.465 0.775 3.605 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.485 ;
        RECT  3.670 -0.115 3.930 0.115 ;
        RECT  3.550 -0.115 3.670 0.275 ;
        RECT  3.290 -0.115 3.550 0.115 ;
        RECT  3.210 -0.115 3.290 0.465 ;
        RECT  2.950 -0.115 3.210 0.115 ;
        RECT  2.830 -0.115 2.950 0.275 ;
        RECT  2.570 -0.115 2.830 0.115 ;
        RECT  2.490 -0.115 2.570 0.305 ;
        RECT  2.220 -0.115 2.490 0.115 ;
        RECT  2.120 -0.115 2.220 0.275 ;
        RECT  1.480 -0.115 2.120 0.115 ;
        RECT  1.400 -0.115 1.480 0.280 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.665 4.010 1.375 ;
        RECT  3.670 1.145 3.930 1.375 ;
        RECT  3.550 0.985 3.670 1.375 ;
        RECT  3.310 1.145 3.550 1.375 ;
        RECT  3.190 1.005 3.310 1.375 ;
        RECT  2.950 1.145 3.190 1.375 ;
        RECT  2.830 1.005 2.950 1.375 ;
        RECT  2.590 1.145 2.830 1.375 ;
        RECT  2.470 1.005 2.590 1.375 ;
        RECT  2.230 1.145 2.470 1.375 ;
        RECT  2.110 0.995 2.230 1.375 ;
        RECT  1.870 1.145 2.110 1.375 ;
        RECT  1.750 0.995 1.870 1.375 ;
        RECT  0.730 1.145 1.750 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.355 3.535 0.465 ;
        RECT  3.465 0.775 3.535 0.905 ;
        RECT  3.395 0.185 3.465 0.465 ;
        RECT  3.395 0.775 3.465 1.055 ;
        RECT  3.045 0.705 3.130 0.795 ;
        RECT  3.045 0.185 3.105 0.485 ;
        RECT  2.675 0.185 2.695 0.485 ;
        RECT  2.650 0.705 2.695 0.795 ;
        RECT  3.285 0.540 3.515 0.620 ;
        RECT  3.215 0.540 3.285 0.935 ;
        RECT  2.570 0.865 3.215 0.935 ;
        RECT  2.500 0.385 2.570 0.935 ;
        RECT  2.390 0.385 2.500 0.465 ;
        RECT  2.390 0.865 2.500 0.935 ;
        RECT  2.240 0.545 2.420 0.620 ;
        RECT  2.310 0.185 2.390 0.465 ;
        RECT  2.310 0.735 2.390 1.055 ;
        RECT  2.170 0.345 2.240 0.925 ;
        RECT  1.985 0.345 2.170 0.415 ;
        RECT  1.670 0.855 2.170 0.925 ;
        RECT  2.020 0.500 2.100 0.775 ;
        RECT  1.600 0.705 2.020 0.775 ;
        RECT  1.915 0.205 1.985 0.415 ;
        RECT  1.730 0.205 1.915 0.275 ;
        RECT  1.590 0.855 1.670 1.055 ;
        RECT  1.520 0.540 1.600 0.775 ;
        RECT  1.410 0.985 1.590 1.055 ;
        RECT  1.380 0.540 1.520 0.620 ;
        RECT  1.260 0.985 1.410 1.075 ;
        RECT  1.310 0.540 1.380 0.915 ;
        RECT  1.270 0.540 1.310 0.620 ;
        RECT  0.930 0.845 1.310 0.915 ;
        RECT  1.200 0.205 1.270 0.620 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.960 0.205 1.200 0.275 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.125 0.985 0.820 1.055 ;
        RECT  0.245 0.350 0.530 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDD4BWP

MACRO LNSNDQD1BWP
    CLASS CORE ;
    FOREIGN LNSNDQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.450 1.055 ;
        RECT  2.370 0.185 2.415 0.465 ;
        RECT  2.370 0.735 2.415 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.520 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.145 2.520 1.375 ;
        RECT  2.170 0.885 2.250 1.375 ;
        RECT  1.900 1.145 2.170 1.375 ;
        RECT  1.800 0.990 1.900 1.375 ;
        RECT  0.730 1.145 1.800 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.345 0.620 ;
        RECT  2.200 0.395 2.270 0.805 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.735 2.200 0.805 ;
        RECT  1.925 0.545 2.120 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.735 2.070 1.055 ;
        RECT  1.855 0.275 1.925 0.915 ;
        RECT  1.770 0.275 1.855 0.355 ;
        RECT  1.710 0.845 1.855 0.915 ;
        RECT  1.630 0.845 1.710 1.055 ;
        RECT  1.420 0.985 1.630 1.055 ;
        RECT  1.425 0.540 1.620 0.620 ;
        RECT  1.345 0.205 1.425 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  0.960 0.205 1.345 0.275 ;
        RECT  0.930 0.845 1.345 0.915 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.125 0.985 0.820 1.055 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDQD1BWP

MACRO LNSNDQD2BWP
    CLASS CORE ;
    FOREIGN LNSNDQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.355 2.485 0.905 ;
        RECT  2.415 0.185 2.430 1.055 ;
        RECT  2.350 0.185 2.415 0.465 ;
        RECT  2.350 0.735 2.415 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.535 -0.115 2.610 0.305 ;
        RECT  2.250 -0.115 2.535 0.115 ;
        RECT  2.170 -0.115 2.250 0.315 ;
        RECT  1.520 -0.115 2.170 0.115 ;
        RECT  1.400 -0.115 1.520 0.135 ;
        RECT  0.700 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.320 0.270 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.975 2.610 1.375 ;
        RECT  2.250 1.145 2.530 1.375 ;
        RECT  2.170 0.885 2.250 1.375 ;
        RECT  1.900 1.145 2.170 1.375 ;
        RECT  1.800 0.990 1.900 1.375 ;
        RECT  0.730 1.145 1.800 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.545 2.345 0.620 ;
        RECT  2.200 0.395 2.270 0.805 ;
        RECT  2.070 0.395 2.200 0.465 ;
        RECT  2.070 0.735 2.200 0.805 ;
        RECT  1.925 0.545 2.120 0.620 ;
        RECT  1.995 0.185 2.070 0.465 ;
        RECT  1.995 0.735 2.070 1.055 ;
        RECT  1.855 0.275 1.925 0.915 ;
        RECT  1.770 0.275 1.855 0.355 ;
        RECT  1.710 0.845 1.855 0.915 ;
        RECT  1.630 0.845 1.710 1.055 ;
        RECT  1.420 0.985 1.630 1.055 ;
        RECT  1.425 0.540 1.620 0.620 ;
        RECT  1.345 0.205 1.425 0.915 ;
        RECT  1.270 0.985 1.420 1.075 ;
        RECT  0.960 0.205 1.345 0.275 ;
        RECT  0.930 0.845 1.345 0.915 ;
        RECT  1.020 0.700 1.230 0.775 ;
        RECT  0.930 0.350 1.020 0.775 ;
        RECT  0.820 0.985 0.980 1.075 ;
        RECT  0.510 0.705 0.930 0.775 ;
        RECT  0.125 0.985 0.820 1.055 ;
        RECT  0.430 0.195 0.510 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.350 0.430 0.420 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDQD2BWP

MACRO LNSNDQD4BWP
    CLASS CORE ;
    FOREIGN LNSNDQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.545 1.740 0.615 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.185 2.845 0.465 ;
        RECT  2.835 0.775 2.845 1.055 ;
        RECT  2.775 0.185 2.835 1.055 ;
        RECT  2.625 0.355 2.775 0.905 ;
        RECT  2.485 0.355 2.625 0.465 ;
        RECT  2.485 0.775 2.625 0.905 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.775 2.485 1.055 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0234 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.685 0.495 0.735 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.485 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.275 ;
        RECT  2.310 -0.115 2.570 0.115 ;
        RECT  2.230 -0.115 2.310 0.305 ;
        RECT  1.960 -0.115 2.230 0.115 ;
        RECT  1.860 -0.115 1.960 0.275 ;
        RECT  1.410 -0.115 1.860 0.115 ;
        RECT  1.330 -0.115 1.410 0.420 ;
        RECT  0.700 -0.115 1.330 0.115 ;
        RECT  0.600 -0.115 0.700 0.260 ;
        RECT  0.310 -0.115 0.600 0.115 ;
        RECT  0.230 -0.115 0.310 0.270 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.665 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 0.985 2.690 1.375 ;
        RECT  2.300 1.145 2.570 1.375 ;
        RECT  2.220 0.925 2.300 1.375 ;
        RECT  1.890 1.145 2.220 1.375 ;
        RECT  1.770 0.995 1.890 1.375 ;
        RECT  0.730 1.145 1.770 1.375 ;
        RECT  0.610 1.130 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.125 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.355 2.555 0.465 ;
        RECT  2.485 0.775 2.555 0.905 ;
        RECT  2.415 0.185 2.485 0.465 ;
        RECT  2.415 0.775 2.485 1.055 ;
        RECT  2.345 0.545 2.535 0.620 ;
        RECT  2.275 0.385 2.345 0.805 ;
        RECT  2.130 0.385 2.275 0.465 ;
        RECT  2.090 0.735 2.275 0.805 ;
        RECT  1.935 0.545 2.195 0.620 ;
        RECT  2.050 0.185 2.130 0.465 ;
        RECT  2.015 0.735 2.090 1.055 ;
        RECT  1.865 0.345 1.935 0.915 ;
        RECT  1.650 0.345 1.865 0.415 ;
        RECT  1.660 0.845 1.865 0.915 ;
        RECT  1.580 0.845 1.660 1.055 ;
        RECT  1.320 0.985 1.580 1.055 ;
        RECT  1.420 0.495 1.495 0.915 ;
        RECT  1.130 0.495 1.420 0.565 ;
        RECT  0.930 0.845 1.420 0.915 ;
        RECT  1.200 0.985 1.320 1.075 ;
        RECT  0.980 0.700 1.210 0.775 ;
        RECT  1.060 0.195 1.130 0.565 ;
        RECT  0.930 0.195 1.060 0.265 ;
        RECT  0.905 0.335 0.980 0.775 ;
        RECT  0.840 0.985 0.960 1.075 ;
        RECT  0.510 0.705 0.905 0.775 ;
        RECT  0.125 0.985 0.840 1.055 ;
        RECT  0.245 0.350 0.530 0.420 ;
        RECT  0.430 0.705 0.510 0.905 ;
        RECT  0.245 0.705 0.430 0.775 ;
        RECT  0.175 0.350 0.245 0.775 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.860 0.125 1.055 ;
        RECT  0.035 0.185 0.105 1.055 ;
    END
END LNSNDQD4BWP

MACRO LNSNQD1BWP
    CLASS CORE ;
    FOREIGN LNSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.375 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.355 2.065 0.905 ;
        RECT  1.995 0.185 2.030 1.060 ;
        RECT  1.950 0.185 1.995 0.465 ;
        RECT  1.950 0.740 1.995 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.980 0.610 1.075 ;
        RECT  0.275 0.980 0.480 1.050 ;
        RECT  0.245 0.825 0.275 1.050 ;
        RECT  0.205 0.495 0.245 1.050 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.115 2.100 0.115 ;
        RECT  1.760 -0.115 1.840 0.430 ;
        RECT  1.090 -0.115 1.760 0.115 ;
        RECT  1.010 -0.115 1.090 0.290 ;
        RECT  0.315 -0.115 1.010 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.145 2.100 1.375 ;
        RECT  1.770 0.800 1.850 1.375 ;
        RECT  1.470 1.145 1.770 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.545 1.920 0.620 ;
        RECT  1.620 0.205 1.690 1.050 ;
        RECT  1.530 0.205 1.620 0.275 ;
        RECT  1.550 0.980 1.620 1.050 ;
        RECT  1.460 0.345 1.540 0.910 ;
        RECT  1.330 0.345 1.460 0.415 ;
        RECT  1.290 0.840 1.460 0.910 ;
        RECT  1.210 0.840 1.290 1.055 ;
        RECT  0.850 0.980 1.210 1.055 ;
        RECT  1.000 0.540 1.200 0.620 ;
        RECT  0.930 0.520 1.000 0.900 ;
        RECT  0.860 0.520 0.930 0.590 ;
        RECT  0.570 0.830 0.930 0.900 ;
        RECT  0.790 0.185 0.860 0.590 ;
        RECT  0.710 0.675 0.850 0.755 ;
        RECT  0.615 0.185 0.790 0.265 ;
        RECT  0.640 0.345 0.710 0.755 ;
        RECT  0.130 0.345 0.640 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSNQD1BWP

MACRO LNSNQD2BWP
    CLASS CORE ;
    FOREIGN LNSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.495 1.375 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.355 2.065 0.905 ;
        RECT  1.995 0.185 2.010 1.060 ;
        RECT  1.930 0.185 1.995 0.465 ;
        RECT  1.930 0.740 1.995 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0290 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.980 0.610 1.075 ;
        RECT  0.275 0.980 0.480 1.050 ;
        RECT  0.245 0.825 0.275 1.050 ;
        RECT  0.205 0.495 0.245 1.050 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 -0.115 2.240 0.115 ;
        RECT  2.100 -0.115 2.200 0.290 ;
        RECT  1.830 -0.115 2.100 0.115 ;
        RECT  1.760 -0.115 1.830 0.450 ;
        RECT  1.090 -0.115 1.760 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.315 -0.115 1.010 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.145 2.240 1.375 ;
        RECT  2.100 0.985 2.200 1.375 ;
        RECT  1.830 1.145 2.100 1.375 ;
        RECT  1.760 0.800 1.830 1.375 ;
        RECT  1.470 1.145 1.760 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.545 1.910 0.620 ;
        RECT  1.620 0.205 1.690 1.050 ;
        RECT  1.510 0.205 1.620 0.275 ;
        RECT  1.550 0.980 1.620 1.050 ;
        RECT  1.460 0.345 1.540 0.910 ;
        RECT  1.330 0.345 1.460 0.415 ;
        RECT  1.290 0.840 1.460 0.910 ;
        RECT  1.210 0.840 1.290 1.055 ;
        RECT  0.850 0.980 1.210 1.055 ;
        RECT  1.000 0.540 1.200 0.620 ;
        RECT  0.930 0.540 1.000 0.900 ;
        RECT  0.810 0.540 0.930 0.610 ;
        RECT  0.570 0.830 0.930 0.900 ;
        RECT  0.665 0.680 0.850 0.755 ;
        RECT  0.740 0.185 0.810 0.610 ;
        RECT  0.610 0.185 0.740 0.265 ;
        RECT  0.595 0.345 0.665 0.755 ;
        RECT  0.130 0.345 0.595 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSNQD2BWP

MACRO LNSNQD4BWP
    CLASS CORE ;
    FOREIGN LNSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.495 1.365 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.275 0.355 2.350 0.485 ;
        RECT  2.275 0.760 2.350 0.905 ;
        RECT  2.065 0.355 2.275 0.905 ;
        RECT  2.035 0.355 2.065 0.485 ;
        RECT  2.030 0.760 2.065 0.905 ;
        RECT  1.950 0.185 2.035 0.485 ;
        RECT  1.950 0.760 2.030 1.040 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.980 0.610 1.075 ;
        RECT  0.275 0.980 0.480 1.050 ;
        RECT  0.245 0.825 0.275 1.050 ;
        RECT  0.205 0.495 0.245 1.050 ;
        RECT  0.175 0.495 0.205 0.905 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.0238 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.340 0.545 0.455 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.465 ;
        RECT  2.250 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.250 0.275 ;
        RECT  1.840 -0.115 2.150 0.115 ;
        RECT  1.760 -0.115 1.840 0.460 ;
        RECT  1.090 -0.115 1.760 0.115 ;
        RECT  1.010 -0.115 1.090 0.310 ;
        RECT  0.315 -0.115 1.010 0.115 ;
        RECT  0.235 -0.115 0.315 0.260 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.685 2.610 1.375 ;
        RECT  2.250 1.145 2.530 1.375 ;
        RECT  2.150 0.985 2.250 1.375 ;
        RECT  1.840 1.145 2.150 1.375 ;
        RECT  1.760 0.750 1.840 1.375 ;
        RECT  1.470 1.145 1.760 1.375 ;
        RECT  1.390 0.980 1.470 1.375 ;
        RECT  0.340 1.145 1.390 1.375 ;
        RECT  0.220 1.130 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.185 2.430 0.485 ;
        RECT  2.350 0.760 2.430 1.040 ;
        RECT  2.345 0.355 2.350 0.485 ;
        RECT  2.345 0.760 2.350 0.905 ;
        RECT  1.950 0.185 1.995 0.485 ;
        RECT  1.950 0.760 1.995 1.040 ;
        RECT  1.670 0.555 1.960 0.625 ;
        RECT  1.600 0.205 1.670 1.050 ;
        RECT  1.530 0.205 1.600 0.275 ;
        RECT  1.550 0.980 1.600 1.050 ;
        RECT  1.460 0.345 1.530 0.910 ;
        RECT  1.350 0.345 1.460 0.415 ;
        RECT  1.270 0.840 1.460 0.910 ;
        RECT  1.190 0.840 1.270 1.055 ;
        RECT  1.020 0.540 1.190 0.620 ;
        RECT  0.850 0.980 1.190 1.055 ;
        RECT  0.950 0.540 1.020 0.900 ;
        RECT  0.810 0.540 0.950 0.610 ;
        RECT  0.580 0.830 0.950 0.900 ;
        RECT  0.665 0.680 0.870 0.755 ;
        RECT  0.740 0.185 0.810 0.610 ;
        RECT  0.610 0.185 0.740 0.265 ;
        RECT  0.595 0.345 0.665 0.755 ;
        RECT  0.130 0.345 0.595 0.415 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.105 0.955 0.125 1.075 ;
        RECT  0.035 0.185 0.105 1.075 ;
    END
END LNSNQD4BWP

MACRO LVLHLD1BWP
    CLASS CORE ;
    FOREIGN LVLHLD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 1.045 ;
        RECT  0.435 0.185 0.455 0.465 ;
        RECT  0.435 0.755 0.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.355 0.520 0.385 0.640 ;
        RECT  0.285 0.340 0.355 0.925 ;
        RECT  0.130 0.340 0.285 0.410 ;
        RECT  0.130 0.855 0.285 0.925 ;
        RECT  0.050 0.205 0.130 0.410 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END LVLHLD1BWP

MACRO LVLHLD2BWP
    CLASS CORE ;
    FOREIGN LVLHLD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.820 ;
        RECT  0.575 0.355 0.595 0.465 ;
        RECT  0.575 0.750 0.595 0.820 ;
        RECT  0.505 0.185 0.575 0.465 ;
        RECT  0.505 0.750 0.575 1.050 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.140 0.495 0.175 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 -0.115 0.840 0.115 ;
        RECT  0.690 -0.115 0.770 0.280 ;
        RECT  0.380 -0.115 0.690 0.115 ;
        RECT  0.260 -0.115 0.380 0.270 ;
        RECT  0.000 -0.115 0.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.145 0.840 1.375 ;
        RECT  0.690 0.950 0.770 1.375 ;
        RECT  0.380 1.145 0.690 1.375 ;
        RECT  0.260 0.995 0.380 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.340 0.435 0.925 ;
        RECT  0.150 0.340 0.365 0.410 ;
        RECT  0.150 0.855 0.365 0.925 ;
        RECT  0.070 0.240 0.150 0.410 ;
        RECT  0.070 0.855 0.150 1.025 ;
    END
END LVLHLD2BWP

MACRO LVLHLD4BWP
    CLASS CORE ;
    FOREIGN LVLHLD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.030 0.465 ;
        RECT  1.015 0.755 1.030 1.045 ;
        RECT  0.950 0.185 1.015 1.045 ;
        RECT  0.805 0.355 0.950 0.905 ;
        RECT  0.670 0.355 0.805 0.465 ;
        RECT  0.670 0.755 0.805 0.905 ;
        RECT  0.590 0.185 0.670 0.465 ;
        RECT  0.590 0.755 0.670 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.470 ;
        RECT  0.870 -0.115 1.130 0.115 ;
        RECT  0.750 -0.115 0.870 0.280 ;
        RECT  0.490 -0.115 0.750 0.115 ;
        RECT  0.410 -0.115 0.490 0.310 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.330 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.670 1.210 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.750 0.980 0.870 1.375 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.910 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.910 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.670 0.355 0.735 0.465 ;
        RECT  0.670 0.755 0.735 0.905 ;
        RECT  0.590 0.185 0.670 0.465 ;
        RECT  0.590 0.755 0.670 1.045 ;
        RECT  0.400 0.545 0.640 0.615 ;
        RECT  0.330 0.390 0.400 0.790 ;
        RECT  0.305 0.390 0.330 0.460 ;
        RECT  0.305 0.720 0.330 0.790 ;
        RECT  0.235 0.200 0.305 0.460 ;
        RECT  0.235 0.720 0.305 1.050 ;
    END
END LVLHLD4BWP

MACRO LVLHLD8BWP
    CLASS CORE ;
    FOREIGN LVLHLD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.725 2.030 0.955 ;
        RECT  1.935 0.185 2.005 0.465 ;
        RECT  1.625 0.355 1.935 0.465 ;
        RECT  1.575 0.185 1.625 0.465 ;
        RECT  1.555 0.185 1.575 0.955 ;
        RECT  1.365 0.355 1.555 0.955 ;
        RECT  1.245 0.355 1.365 0.465 ;
        RECT  0.770 0.725 1.365 0.955 ;
        RECT  1.175 0.185 1.245 0.465 ;
        RECT  0.865 0.355 1.175 0.465 ;
        RECT  0.795 0.185 0.865 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.475 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.720 -0.115 1.840 0.275 ;
        RECT  1.460 -0.115 1.720 0.115 ;
        RECT  1.340 -0.115 1.460 0.275 ;
        RECT  1.080 -0.115 1.340 0.115 ;
        RECT  0.960 -0.115 1.080 0.275 ;
        RECT  0.690 -0.115 0.960 0.115 ;
        RECT  0.610 -0.115 0.690 0.465 ;
        RECT  0.340 -0.115 0.610 0.115 ;
        RECT  0.220 -0.115 0.340 0.230 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.675 2.190 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.720 1.025 1.840 1.375 ;
        RECT  1.460 1.145 1.720 1.375 ;
        RECT  1.340 1.025 1.460 1.375 ;
        RECT  1.080 1.145 1.340 1.375 ;
        RECT  0.960 1.025 1.080 1.375 ;
        RECT  0.690 1.145 0.960 1.375 ;
        RECT  0.610 0.750 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.985 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.725 2.030 0.955 ;
        RECT  1.935 0.185 2.005 0.465 ;
        RECT  1.645 0.355 1.935 0.465 ;
        RECT  1.245 0.355 1.295 0.465 ;
        RECT  0.770 0.725 1.295 0.955 ;
        RECT  1.175 0.185 1.245 0.465 ;
        RECT  0.865 0.355 1.175 0.465 ;
        RECT  0.795 0.185 0.865 0.465 ;
        RECT  1.680 0.540 1.980 0.620 ;
        RECT  0.515 0.545 1.120 0.615 ;
        RECT  0.425 0.185 0.515 1.070 ;
        RECT  0.125 0.300 0.425 0.390 ;
        RECT  0.125 0.845 0.425 0.915 ;
        RECT  0.055 0.220 0.125 0.390 ;
        RECT  0.055 0.845 0.125 0.995 ;
    END
END LVLHLD8BWP

MACRO LVLLHCD1BWP
    CLASS CORE ;
    FOREIGN LVLLHCD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.0924 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.655 1.475 0.725 1.745 ;
        RECT  0.385 1.675 0.655 1.745 ;
        RECT  0.315 1.475 0.385 2.335 ;
        RECT  0.275 1.475 0.315 1.760 ;
        RECT  0.275 2.055 0.315 2.335 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1040 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 1.615 0.945 1.975 ;
        RECT  0.700 1.905 0.875 1.975 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.265 0.495 2.355 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.115 3.640 0.115 ;
        RECT  3.130 -0.115 3.270 0.420 ;
        RECT  0.000 -0.115 3.130 0.115 ;
        RECT  3.270 2.405 3.640 2.635 ;
        RECT  3.130 2.100 3.270 2.635 ;
        RECT  1.810 2.405 3.130 2.635 ;
        RECT  1.730 2.215 1.810 2.635 ;
        RECT  1.450 2.405 1.730 2.635 ;
        RECT  1.370 2.215 1.450 2.635 ;
        RECT  1.090 2.405 1.370 2.635 ;
        RECT  1.010 2.215 1.090 2.635 ;
        RECT  0.730 2.405 1.010 2.635 ;
        RECT  0.650 2.215 0.730 2.635 ;
        RECT  0.000 2.405 0.650 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.655 1.495 2.145 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.360 1.145 3.640 1.375 ;
        RECT  3.240 0.855 3.360 1.675 ;
        RECT  0.535 1.145 3.240 1.375 ;
        RECT  0.525 1.145 0.535 1.600 ;
        RECT  0.465 0.915 0.525 1.600 ;
        RECT  0.455 0.915 0.465 1.375 ;
        RECT  0.000 1.145 0.455 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.985 0.205 3.055 1.055 ;
        RECT  2.725 0.205 2.985 0.275 ;
        RECT  2.240 0.985 2.985 1.055 ;
        RECT  2.835 0.350 2.905 0.915 ;
        RECT  2.035 0.845 2.835 0.915 ;
        RECT  2.655 0.205 2.725 0.470 ;
        RECT  1.645 0.205 2.655 0.275 ;
        RECT  1.825 0.350 2.570 0.420 ;
        RECT  2.280 1.455 2.360 2.125 ;
        RECT  1.985 2.055 2.280 2.125 ;
        RECT  1.965 0.755 2.035 1.055 ;
        RECT  1.915 2.055 1.985 2.335 ;
        RECT  1.430 0.755 1.965 0.825 ;
        RECT  1.630 2.055 1.915 2.125 ;
        RECT  1.755 0.350 1.825 0.635 ;
        RECT  0.890 0.565 1.755 0.635 ;
        RECT  1.575 0.205 1.645 0.470 ;
        RECT  1.550 2.055 1.630 2.335 ;
        RECT  0.820 0.205 1.575 0.275 ;
        RECT  1.270 2.055 1.550 2.125 ;
        RECT  0.665 0.375 1.495 0.445 ;
        RECT  1.190 2.055 1.270 2.335 ;
        RECT  0.910 2.055 1.190 2.125 ;
        RECT  0.830 2.055 0.910 2.335 ;
        RECT  0.820 0.565 0.890 0.835 ;
        RECT  0.535 2.055 0.830 2.125 ;
        RECT  0.465 0.765 0.820 0.835 ;
        RECT  0.595 0.375 0.665 0.690 ;
        RECT  0.325 0.375 0.595 0.445 ;
        RECT  0.465 2.055 0.535 2.335 ;
        RECT  0.395 0.560 0.465 0.835 ;
        RECT  0.325 0.915 0.345 1.045 ;
        RECT  0.255 0.375 0.325 1.045 ;
    END
END LVLLHCD1BWP

MACRO LVLLHCD2BWP
    CLASS CORE ;
    FOREIGN LVLLHCD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1283 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 1.475 0.885 1.745 ;
        RECT  0.525 1.675 0.815 1.745 ;
        RECT  0.455 1.475 0.525 2.165 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1092 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.615 1.090 1.975 ;
        RECT  0.775 1.905 1.010 1.975 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.495 2.075 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.410 -0.115 3.780 0.115 ;
        RECT  3.270 -0.115 3.410 0.420 ;
        RECT  0.000 -0.115 3.270 0.115 ;
        RECT  3.410 2.405 3.780 2.635 ;
        RECT  3.270 2.100 3.410 2.635 ;
        RECT  1.965 2.405 3.270 2.635 ;
        RECT  1.895 2.215 1.965 2.635 ;
        RECT  1.605 2.405 1.895 2.635 ;
        RECT  1.535 2.215 1.605 2.635 ;
        RECT  1.245 2.405 1.535 2.635 ;
        RECT  1.175 2.215 1.245 2.635 ;
        RECT  0.885 2.405 1.175 2.635 ;
        RECT  0.815 2.215 0.885 2.635 ;
        RECT  0.000 2.405 0.815 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 1.495 2.285 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.145 3.780 1.375 ;
        RECT  3.380 0.855 3.500 1.675 ;
        RECT  0.710 1.145 3.380 1.375 ;
        RECT  0.630 1.145 0.710 1.600 ;
        RECT  0.530 1.145 0.630 1.375 ;
        RECT  0.450 0.915 0.530 1.375 ;
        RECT  0.350 1.145 0.450 1.375 ;
        RECT  0.270 1.145 0.350 1.760 ;
        RECT  0.000 1.145 0.270 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.015 0.205 3.085 1.055 ;
        RECT  2.755 0.205 3.015 0.275 ;
        RECT  2.400 0.985 3.015 1.055 ;
        RECT  2.865 0.350 2.935 0.820 ;
        RECT  2.215 0.740 2.865 0.820 ;
        RECT  2.685 0.205 2.755 0.470 ;
        RECT  1.675 0.205 2.685 0.275 ;
        RECT  1.855 0.350 2.600 0.420 ;
        RECT  2.420 1.455 2.500 2.135 ;
        RECT  2.150 2.055 2.420 2.135 ;
        RECT  2.145 0.740 2.215 1.055 ;
        RECT  2.070 2.055 2.150 2.325 ;
        RECT  1.605 0.985 2.145 1.055 ;
        RECT  1.790 2.055 2.070 2.135 ;
        RECT  1.785 0.350 1.855 0.635 ;
        RECT  1.710 2.055 1.790 2.325 ;
        RECT  1.240 0.565 1.785 0.635 ;
        RECT  1.430 2.055 1.710 2.135 ;
        RECT  1.605 0.205 1.675 0.470 ;
        RECT  0.850 0.205 1.605 0.275 ;
        RECT  1.535 0.730 1.605 1.055 ;
        RECT  0.665 0.375 1.520 0.445 ;
        RECT  1.350 2.055 1.430 2.325 ;
        RECT  1.070 2.055 1.350 2.135 ;
        RECT  1.170 0.565 1.240 0.835 ;
        RECT  0.465 0.765 1.170 0.835 ;
        RECT  0.990 2.055 1.070 2.335 ;
        RECT  0.745 2.055 0.990 2.135 ;
        RECT  0.675 2.055 0.745 2.325 ;
        RECT  0.350 2.245 0.675 2.325 ;
        RECT  0.595 0.375 0.665 0.690 ;
        RECT  0.325 0.375 0.595 0.445 ;
        RECT  0.395 0.560 0.465 0.835 ;
        RECT  0.270 2.045 0.350 2.325 ;
        RECT  0.325 0.915 0.345 1.045 ;
        RECT  0.255 0.375 0.325 1.045 ;
    END
END LVLLHCD2BWP

MACRO LVLLHCD4BWP
    CLASS CORE ;
    FOREIGN LVLLHCD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.2467 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.465 1.305 1.745 ;
        RECT  0.945 1.615 1.235 1.745 ;
        RECT  0.735 2.055 0.970 2.175 ;
        RECT  0.875 1.465 0.945 1.745 ;
        RECT  0.735 1.615 0.875 1.745 ;
        RECT  0.585 1.615 0.735 2.175 ;
        RECT  0.525 1.465 0.585 2.175 ;
        RECT  0.515 1.465 0.525 1.745 ;
        RECT  0.515 2.055 0.525 2.175 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1156 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 1.905 2.100 1.975 ;
        RECT  1.715 1.615 1.785 1.975 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.405 0.495 2.495 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 -0.115 4.060 0.115 ;
        RECT  3.550 -0.115 3.690 0.420 ;
        RECT  0.000 -0.115 3.550 0.115 ;
        RECT  3.690 2.405 4.060 2.635 ;
        RECT  3.550 2.100 3.690 2.635 ;
        RECT  2.390 2.405 3.550 2.635 ;
        RECT  2.310 2.215 2.390 2.635 ;
        RECT  2.030 2.405 2.310 2.635 ;
        RECT  1.950 2.215 2.030 2.635 ;
        RECT  1.670 2.405 1.950 2.635 ;
        RECT  1.590 2.215 1.670 2.635 ;
        RECT  1.310 2.405 1.590 2.635 ;
        RECT  1.230 2.215 1.310 2.635 ;
        RECT  0.000 2.405 1.230 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.495 2.765 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.780 1.145 4.060 1.375 ;
        RECT  3.660 0.855 3.780 1.675 ;
        RECT  1.150 1.145 3.660 1.375 ;
        RECT  1.030 1.145 1.150 1.535 ;
        RECT  0.790 1.145 1.030 1.375 ;
        RECT  0.670 1.145 0.790 1.535 ;
        RECT  0.590 1.145 0.670 1.375 ;
        RECT  0.510 0.915 0.590 1.375 ;
        RECT  0.410 1.145 0.510 1.375 ;
        RECT  0.330 1.145 0.410 1.755 ;
        RECT  0.000 1.145 0.330 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.235 1.465 1.305 1.745 ;
        RECT  0.945 1.615 1.235 1.745 ;
        RECT  0.805 2.055 0.970 2.175 ;
        RECT  0.875 1.465 0.945 1.745 ;
        RECT  0.805 1.615 0.875 1.745 ;
        RECT  3.265 0.205 3.335 1.055 ;
        RECT  2.995 0.205 3.265 0.275 ;
        RECT  2.870 0.985 3.265 1.055 ;
        RECT  3.105 0.350 3.175 0.720 ;
        RECT  2.655 0.650 3.105 0.720 ;
        RECT  2.925 0.205 2.995 0.470 ;
        RECT  2.900 1.455 2.980 2.125 ;
        RECT  1.915 0.205 2.925 0.275 ;
        RECT  2.570 2.045 2.900 2.125 ;
        RECT  2.095 0.350 2.840 0.420 ;
        RECT  2.585 0.650 2.655 1.055 ;
        RECT  1.845 0.985 2.585 1.055 ;
        RECT  2.490 2.045 2.570 2.325 ;
        RECT  2.210 2.045 2.490 2.125 ;
        RECT  2.130 2.045 2.210 2.325 ;
        RECT  1.850 2.045 2.130 2.125 ;
        RECT  2.025 0.350 2.095 0.635 ;
        RECT  1.650 0.565 2.025 0.635 ;
        RECT  1.845 0.205 1.915 0.470 ;
        RECT  1.770 2.045 1.850 2.325 ;
        RECT  1.450 0.205 1.845 0.275 ;
        RECT  1.775 0.730 1.845 1.055 ;
        RECT  1.490 2.045 1.770 2.125 ;
        RECT  0.725 0.375 1.765 0.445 ;
        RECT  1.575 0.565 1.650 1.065 ;
        RECT  1.570 1.455 1.645 1.975 ;
        RECT  1.570 0.765 1.575 1.065 ;
        RECT  0.525 0.765 1.570 0.835 ;
        RECT  0.890 1.905 1.570 1.975 ;
        RECT  1.410 2.045 1.490 2.325 ;
        RECT  1.130 2.045 1.410 2.125 ;
        RECT  1.050 2.045 1.130 2.325 ;
        RECT  0.410 2.255 1.050 2.325 ;
        RECT  0.655 0.375 0.725 0.690 ;
        RECT  0.375 0.375 0.655 0.445 ;
        RECT  0.455 0.560 0.525 0.835 ;
        RECT  0.330 2.045 0.410 2.325 ;
        RECT  0.375 0.915 0.405 1.045 ;
        RECT  0.305 0.375 0.375 1.045 ;
    END
END LVLLHCD4BWP

MACRO LVLLHCD8BWP
    CLASS CORE ;
    FOREIGN LVLLHCD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.4606 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.895 1.465 1.965 1.745 ;
        RECT  1.605 1.615 1.895 1.745 ;
        RECT  1.155 2.055 1.630 2.175 ;
        RECT  1.535 1.465 1.605 1.745 ;
        RECT  1.245 1.615 1.535 1.745 ;
        RECT  1.165 1.465 1.245 1.745 ;
        RECT  1.155 1.615 1.165 1.745 ;
        RECT  0.945 1.615 1.155 2.175 ;
        RECT  0.885 1.615 0.945 1.745 ;
        RECT  0.430 2.055 0.945 2.175 ;
        RECT  0.815 1.465 0.885 1.745 ;
        RECT  0.525 1.615 0.815 1.745 ;
        RECT  0.455 1.465 0.525 1.745 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.2188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 1.905 3.160 1.975 ;
        RECT  2.555 1.615 2.625 1.975 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.545 3.185 0.905 ;
        RECT  2.865 0.545 3.115 0.615 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 -0.115 5.180 0.115 ;
        RECT  4.680 -0.115 4.810 0.420 ;
        RECT  0.000 -0.115 4.680 0.115 ;
        RECT  4.810 2.405 5.180 2.635 ;
        RECT  4.680 2.100 4.810 2.635 ;
        RECT  4.490 2.405 4.680 2.635 ;
        RECT  4.410 2.035 4.490 2.635 ;
        RECT  4.130 2.405 4.410 2.635 ;
        RECT  4.050 2.205 4.130 2.635 ;
        RECT  3.770 2.405 4.050 2.635 ;
        RECT  3.690 2.205 3.770 2.635 ;
        RECT  3.410 2.405 3.690 2.635 ;
        RECT  3.330 2.205 3.410 2.635 ;
        RECT  3.050 2.405 3.330 2.635 ;
        RECT  2.970 2.205 3.050 2.635 ;
        RECT  2.690 2.405 2.970 2.635 ;
        RECT  2.610 2.205 2.690 2.635 ;
        RECT  2.330 2.405 2.610 2.635 ;
        RECT  2.250 2.205 2.330 2.635 ;
        RECT  1.970 2.405 2.250 2.635 ;
        RECT  1.890 2.205 1.970 2.635 ;
        RECT  0.000 2.405 1.890 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.055 1.495 3.545 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.900 1.145 5.180 1.375 ;
        RECT  4.780 0.855 4.900 1.675 ;
        RECT  2.150 1.145 4.780 1.375 ;
        RECT  2.070 1.145 2.150 1.745 ;
        RECT  1.810 1.145 2.070 1.375 ;
        RECT  1.690 1.145 1.810 1.535 ;
        RECT  1.450 1.145 1.690 1.375 ;
        RECT  1.330 1.145 1.450 1.535 ;
        RECT  1.090 1.145 1.330 1.375 ;
        RECT  0.970 1.145 1.090 1.535 ;
        RECT  0.730 1.145 0.970 1.375 ;
        RECT  0.610 1.145 0.730 1.535 ;
        RECT  0.530 1.145 0.610 1.375 ;
        RECT  0.450 0.915 0.530 1.375 ;
        RECT  0.350 1.145 0.450 1.375 ;
        RECT  0.270 1.145 0.350 1.755 ;
        RECT  0.000 1.145 0.270 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.895 1.465 1.965 1.745 ;
        RECT  1.605 1.615 1.895 1.745 ;
        RECT  1.225 2.055 1.630 2.175 ;
        RECT  1.535 1.465 1.605 1.745 ;
        RECT  1.245 1.615 1.535 1.745 ;
        RECT  1.225 1.465 1.245 1.745 ;
        RECT  0.815 1.465 0.875 1.745 ;
        RECT  0.430 2.055 0.875 2.175 ;
        RECT  0.525 1.615 0.815 1.745 ;
        RECT  0.455 1.465 0.525 1.745 ;
        RECT  4.230 2.045 4.310 2.325 ;
        RECT  3.950 2.045 4.230 2.125 ;
        RECT  3.870 2.045 3.950 2.325 ;
        RECT  3.875 0.205 3.945 1.055 ;
        RECT  3.615 0.205 3.875 0.275 ;
        RECT  3.640 0.985 3.875 1.055 ;
        RECT  3.760 2.045 3.870 2.125 ;
        RECT  3.725 0.350 3.795 0.810 ;
        RECT  3.680 1.455 3.760 2.125 ;
        RECT  3.440 0.740 3.725 0.810 ;
        RECT  3.590 2.045 3.680 2.125 ;
        RECT  3.545 0.205 3.615 0.470 ;
        RECT  3.510 2.045 3.590 2.325 ;
        RECT  2.540 0.205 3.545 0.275 ;
        RECT  3.230 2.045 3.510 2.125 ;
        RECT  2.680 0.375 3.460 0.445 ;
        RECT  3.360 0.740 3.440 1.055 ;
        RECT  2.665 0.985 3.360 1.055 ;
        RECT  3.150 2.045 3.230 2.325 ;
        RECT  2.870 2.045 3.150 2.125 ;
        RECT  2.790 2.045 2.870 2.325 ;
        RECT  2.510 2.045 2.790 2.125 ;
        RECT  2.610 0.375 2.680 0.635 ;
        RECT  2.595 0.755 2.665 1.055 ;
        RECT  2.245 0.565 2.610 0.635 ;
        RECT  2.390 0.755 2.595 0.825 ;
        RECT  2.460 0.205 2.540 0.470 ;
        RECT  2.430 2.045 2.510 2.325 ;
        RECT  2.080 0.205 2.460 0.275 ;
        RECT  2.245 0.970 2.460 1.040 ;
        RECT  2.150 2.045 2.430 2.125 ;
        RECT  2.355 1.455 2.425 1.975 ;
        RECT  1.995 0.375 2.380 0.445 ;
        RECT  1.270 1.905 2.355 1.975 ;
        RECT  2.175 0.565 2.245 1.040 ;
        RECT  0.465 0.765 2.175 0.835 ;
        RECT  2.070 2.045 2.150 2.325 ;
        RECT  1.790 2.045 2.070 2.125 ;
        RECT  1.925 0.185 1.995 0.445 ;
        RECT  0.665 0.375 1.925 0.445 ;
        RECT  1.710 2.045 1.790 2.325 ;
        RECT  0.350 2.255 1.710 2.325 ;
        RECT  0.480 1.900 0.780 1.980 ;
        RECT  0.595 0.375 0.665 0.690 ;
        RECT  0.325 0.375 0.595 0.445 ;
        RECT  0.395 0.560 0.465 0.835 ;
        RECT  0.270 2.045 0.350 2.325 ;
        RECT  0.325 0.915 0.345 1.045 ;
        RECT  0.255 0.375 0.325 1.045 ;
    END
END LVLLHCD8BWP

MACRO LVLLHCLOD1BWP
    CLASS CORE ;
    FOREIGN LVLLHCLOD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.185 0.565 0.445 ;
        RECT  0.525 0.765 0.565 1.045 ;
        RECT  0.455 0.185 0.525 1.045 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.905 2.375 1.975 ;
        RECT  1.155 1.565 1.225 1.975 ;
        RECT  0.725 1.565 1.155 1.635 ;
        RECT  0.655 1.565 0.725 1.835 ;
        RECT  0.495 1.765 0.655 1.835 ;
        RECT  0.425 1.765 0.495 2.000 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.495 2.915 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.920 -0.115 4.340 0.115 ;
        RECT  3.780 -0.115 3.920 0.420 ;
        RECT  0.745 -0.115 3.780 0.115 ;
        RECT  0.675 -0.115 0.745 0.440 ;
        RECT  0.000 -0.115 0.675 0.115 ;
        RECT  3.920 2.405 4.340 2.635 ;
        RECT  3.780 2.100 3.920 2.635 ;
        RECT  2.410 2.405 3.780 2.635 ;
        RECT  2.330 2.215 2.410 2.635 ;
        RECT  2.050 2.405 2.330 2.635 ;
        RECT  1.970 2.215 2.050 2.635 ;
        RECT  1.690 2.405 1.970 2.635 ;
        RECT  1.610 2.215 1.690 2.635 ;
        RECT  1.330 2.405 1.610 2.635 ;
        RECT  1.250 2.215 1.330 2.635 ;
        RECT  0.000 2.405 1.250 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.495 2.765 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.145 4.340 1.375 ;
        RECT  3.940 0.855 4.060 1.675 ;
        RECT  1.150 1.145 3.940 1.375 ;
        RECT  1.125 1.145 1.150 1.495 ;
        RECT  1.055 0.915 1.125 1.495 ;
        RECT  1.030 1.145 1.055 1.495 ;
        RECT  0.770 1.145 1.030 1.375 ;
        RECT  0.750 1.145 0.770 1.495 ;
        RECT  0.670 0.755 0.750 1.495 ;
        RECT  0.650 1.145 0.670 1.495 ;
        RECT  0.390 1.145 0.650 1.375 ;
        RECT  0.310 1.145 0.390 1.550 ;
        RECT  0.000 1.145 0.310 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.595 0.205 3.665 1.055 ;
        RECT  3.325 0.205 3.595 0.275 ;
        RECT  2.840 0.985 3.595 1.055 ;
        RECT  3.435 0.350 3.505 0.915 ;
        RECT  2.635 0.845 3.435 0.915 ;
        RECT  3.255 0.205 3.325 0.470 ;
        RECT  2.245 0.205 3.255 0.275 ;
        RECT  2.425 0.350 3.170 0.420 ;
        RECT  2.880 1.455 2.960 2.125 ;
        RECT  2.590 2.055 2.880 2.125 ;
        RECT  2.565 0.755 2.635 1.055 ;
        RECT  2.510 2.055 2.590 2.335 ;
        RECT  2.030 0.755 2.565 0.825 ;
        RECT  2.230 2.055 2.510 2.125 ;
        RECT  2.355 0.350 2.425 0.635 ;
        RECT  1.490 0.565 2.355 0.635 ;
        RECT  2.175 0.205 2.245 0.470 ;
        RECT  2.150 2.055 2.230 2.335 ;
        RECT  1.420 0.205 2.175 0.275 ;
        RECT  1.870 2.055 2.150 2.125 ;
        RECT  1.265 0.375 2.095 0.445 ;
        RECT  1.790 2.055 1.870 2.335 ;
        RECT  1.510 2.055 1.790 2.125 ;
        RECT  1.430 2.055 1.510 2.335 ;
        RECT  1.420 0.565 1.490 0.835 ;
        RECT  1.140 2.055 1.430 2.125 ;
        RECT  1.065 0.765 1.420 0.835 ;
        RECT  1.195 0.375 1.265 0.690 ;
        RECT  0.925 0.375 1.195 0.445 ;
        RECT  1.060 2.055 1.140 2.315 ;
        RECT  0.995 0.560 1.065 0.835 ;
        RECT  0.290 2.245 1.060 2.315 ;
        RECT  0.870 1.705 0.950 2.165 ;
        RECT  0.925 0.915 0.945 1.045 ;
        RECT  0.855 0.375 0.925 1.045 ;
        RECT  0.580 1.905 0.870 1.975 ;
        RECT  0.320 2.095 0.770 2.165 ;
        RECT  0.495 1.470 0.565 1.695 ;
        RECT  0.320 1.625 0.495 1.695 ;
        RECT  0.240 1.625 0.320 2.165 ;
    END
END LVLLHCLOD1BWP

MACRO LVLLHCLOD2BWP
    CLASS CORE ;
    FOREIGN LVLLHCLOD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.185 0.565 0.445 ;
        RECT  0.525 0.765 0.565 1.045 ;
        RECT  0.495 0.185 0.525 1.045 ;
        RECT  0.455 0.375 0.495 0.835 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.905 2.375 1.975 ;
        RECT  1.155 1.565 1.225 1.975 ;
        RECT  0.725 1.565 1.155 1.635 ;
        RECT  0.655 1.565 0.725 1.835 ;
        RECT  0.495 1.765 0.655 1.835 ;
        RECT  0.425 1.765 0.495 2.000 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.495 2.915 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.920 -0.115 4.340 0.115 ;
        RECT  3.780 -0.115 3.920 0.420 ;
        RECT  0.745 -0.115 3.780 0.115 ;
        RECT  0.675 -0.115 0.745 0.440 ;
        RECT  0.390 -0.115 0.675 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        RECT  3.920 2.405 4.340 2.635 ;
        RECT  3.780 2.100 3.920 2.635 ;
        RECT  2.410 2.405 3.780 2.635 ;
        RECT  2.330 2.215 2.410 2.635 ;
        RECT  2.050 2.405 2.330 2.635 ;
        RECT  1.970 2.215 2.050 2.635 ;
        RECT  1.690 2.405 1.970 2.635 ;
        RECT  1.610 2.215 1.690 2.635 ;
        RECT  1.330 2.405 1.610 2.635 ;
        RECT  1.250 2.215 1.330 2.635 ;
        RECT  0.000 2.405 1.250 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.495 2.765 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.145 4.340 1.375 ;
        RECT  3.940 0.855 4.060 1.675 ;
        RECT  1.150 1.145 3.940 1.375 ;
        RECT  1.125 1.145 1.150 1.495 ;
        RECT  1.055 0.915 1.125 1.495 ;
        RECT  1.030 1.145 1.055 1.495 ;
        RECT  0.770 1.145 1.030 1.375 ;
        RECT  0.750 1.145 0.770 1.495 ;
        RECT  0.670 0.755 0.750 1.495 ;
        RECT  0.650 1.145 0.670 1.495 ;
        RECT  0.390 1.145 0.650 1.375 ;
        RECT  0.310 0.915 0.390 1.550 ;
        RECT  0.000 1.145 0.310 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.595 0.205 3.665 1.055 ;
        RECT  3.325 0.205 3.595 0.275 ;
        RECT  2.840 0.985 3.595 1.055 ;
        RECT  3.435 0.350 3.505 0.915 ;
        RECT  2.635 0.845 3.435 0.915 ;
        RECT  3.255 0.205 3.325 0.470 ;
        RECT  2.245 0.205 3.255 0.275 ;
        RECT  2.425 0.350 3.170 0.420 ;
        RECT  2.880 1.455 2.960 2.125 ;
        RECT  2.590 2.055 2.880 2.125 ;
        RECT  2.565 0.755 2.635 1.055 ;
        RECT  2.510 2.055 2.590 2.335 ;
        RECT  2.030 0.755 2.565 0.825 ;
        RECT  2.230 2.055 2.510 2.125 ;
        RECT  2.355 0.350 2.425 0.635 ;
        RECT  1.490 0.565 2.355 0.635 ;
        RECT  2.175 0.205 2.245 0.470 ;
        RECT  2.150 2.055 2.230 2.335 ;
        RECT  1.420 0.205 2.175 0.275 ;
        RECT  1.870 2.055 2.150 2.125 ;
        RECT  1.265 0.375 2.095 0.445 ;
        RECT  1.790 2.055 1.870 2.335 ;
        RECT  1.510 2.055 1.790 2.125 ;
        RECT  1.430 2.055 1.510 2.335 ;
        RECT  1.420 0.565 1.490 0.835 ;
        RECT  1.140 2.055 1.430 2.125 ;
        RECT  1.065 0.765 1.420 0.835 ;
        RECT  1.195 0.375 1.265 0.690 ;
        RECT  0.925 0.375 1.195 0.445 ;
        RECT  1.060 2.055 1.140 2.315 ;
        RECT  0.995 0.560 1.065 0.835 ;
        RECT  0.290 2.245 1.060 2.315 ;
        RECT  0.870 1.705 0.950 2.165 ;
        RECT  0.925 0.915 0.945 1.045 ;
        RECT  0.855 0.375 0.925 1.045 ;
        RECT  0.580 1.905 0.870 1.975 ;
        RECT  0.320 2.095 0.770 2.165 ;
        RECT  0.495 1.470 0.565 1.695 ;
        RECT  0.320 1.625 0.495 1.695 ;
        RECT  0.240 1.625 0.320 2.165 ;
    END
END LVLLHCLOD2BWP

MACRO LVLLHCLOD4BWP
    CLASS CORE ;
    FOREIGN LVLLHCLOD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.185 0.665 0.495 ;
        RECT  0.595 0.735 0.665 1.045 ;
        RECT  0.455 0.375 0.595 0.495 ;
        RECT  0.455 0.735 0.595 0.835 ;
        RECT  0.305 0.375 0.455 0.835 ;
        RECT  0.245 0.185 0.305 1.045 ;
        RECT  0.235 0.185 0.245 0.495 ;
        RECT  0.235 0.735 0.245 1.045 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.1280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 1.905 2.475 1.975 ;
        RECT  1.295 1.565 1.365 1.975 ;
        RECT  0.825 1.565 1.295 1.635 ;
        RECT  0.755 1.565 0.825 1.835 ;
        RECT  0.595 1.765 0.755 1.835 ;
        RECT  0.525 1.765 0.595 2.000 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.495 2.915 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.990 -0.115 4.340 0.115 ;
        RECT  3.850 -0.115 3.990 0.420 ;
        RECT  0.845 -0.115 3.850 0.115 ;
        RECT  0.775 -0.115 0.845 0.440 ;
        RECT  0.490 -0.115 0.775 0.115 ;
        RECT  0.410 -0.115 0.490 0.300 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.440 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        RECT  3.990 2.405 4.340 2.635 ;
        RECT  3.850 2.100 3.990 2.635 ;
        RECT  2.510 2.405 3.850 2.635 ;
        RECT  2.430 2.215 2.510 2.635 ;
        RECT  2.150 2.405 2.430 2.635 ;
        RECT  2.070 2.215 2.150 2.635 ;
        RECT  1.790 2.405 2.070 2.635 ;
        RECT  1.710 2.215 1.790 2.635 ;
        RECT  1.430 2.405 1.710 2.635 ;
        RECT  1.350 2.215 1.430 2.635 ;
        RECT  0.000 2.405 1.350 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 1.495 2.905 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.145 4.340 1.375 ;
        RECT  3.940 0.855 4.060 1.675 ;
        RECT  1.250 1.145 3.940 1.375 ;
        RECT  1.225 1.145 1.250 1.495 ;
        RECT  1.155 0.915 1.225 1.495 ;
        RECT  1.130 1.145 1.155 1.495 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.850 1.145 0.870 1.495 ;
        RECT  0.770 0.755 0.850 1.495 ;
        RECT  0.750 1.145 0.770 1.495 ;
        RECT  0.490 1.145 0.750 1.375 ;
        RECT  0.410 0.915 0.490 1.550 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.755 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.595 0.185 0.665 0.495 ;
        RECT  0.595 0.735 0.665 1.045 ;
        RECT  0.525 0.375 0.595 0.495 ;
        RECT  0.525 0.735 0.595 0.835 ;
        RECT  3.685 0.205 3.755 1.055 ;
        RECT  3.425 0.205 3.685 0.275 ;
        RECT  2.940 0.985 3.685 1.055 ;
        RECT  3.535 0.350 3.605 0.915 ;
        RECT  2.735 0.845 3.535 0.915 ;
        RECT  3.355 0.205 3.425 0.470 ;
        RECT  2.345 0.205 3.355 0.275 ;
        RECT  2.525 0.350 3.270 0.420 ;
        RECT  2.980 1.455 3.060 2.125 ;
        RECT  2.685 2.055 2.980 2.125 ;
        RECT  2.665 0.755 2.735 1.055 ;
        RECT  2.615 2.055 2.685 2.335 ;
        RECT  2.130 0.755 2.665 0.825 ;
        RECT  2.330 2.055 2.615 2.125 ;
        RECT  2.455 0.350 2.525 0.635 ;
        RECT  1.590 0.565 2.455 0.635 ;
        RECT  2.275 0.205 2.345 0.470 ;
        RECT  2.250 2.055 2.330 2.335 ;
        RECT  1.530 0.205 2.275 0.275 ;
        RECT  1.970 2.055 2.250 2.125 ;
        RECT  1.445 0.375 2.195 0.445 ;
        RECT  1.890 2.055 1.970 2.335 ;
        RECT  1.610 2.055 1.890 2.125 ;
        RECT  1.530 2.055 1.610 2.335 ;
        RECT  1.520 0.565 1.590 0.835 ;
        RECT  1.240 2.055 1.530 2.125 ;
        RECT  1.165 0.765 1.520 0.835 ;
        RECT  1.375 0.210 1.445 0.445 ;
        RECT  1.365 0.375 1.375 0.445 ;
        RECT  1.295 0.375 1.365 0.690 ;
        RECT  1.025 0.375 1.295 0.445 ;
        RECT  1.160 2.055 1.240 2.315 ;
        RECT  1.095 0.560 1.165 0.835 ;
        RECT  0.390 2.245 1.160 2.315 ;
        RECT  1.025 0.915 1.045 1.045 ;
        RECT  0.975 1.705 1.045 2.165 ;
        RECT  0.955 0.375 1.025 1.045 ;
        RECT  0.680 1.905 0.975 1.975 ;
        RECT  0.415 2.095 0.870 2.165 ;
        RECT  0.595 1.470 0.665 1.695 ;
        RECT  0.415 1.625 0.595 1.695 ;
        RECT  0.345 1.625 0.415 2.165 ;
    END
END LVLLHCLOD4BWP

MACRO LVLLHCLOD8BWP
    CLASS CORE ;
    FOREIGN LVLLHCLOD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.315 0.185 1.385 0.475 ;
        RECT  1.315 0.735 1.385 1.045 ;
        RECT  1.025 0.375 1.315 0.475 ;
        RECT  1.025 0.735 1.315 0.835 ;
        RECT  0.955 0.185 1.025 0.475 ;
        RECT  0.955 0.735 1.025 1.045 ;
        RECT  0.875 0.375 0.955 0.475 ;
        RECT  0.875 0.735 0.955 0.835 ;
        RECT  0.665 0.375 0.875 0.835 ;
        RECT  0.595 0.185 0.665 0.475 ;
        RECT  0.595 0.735 0.665 1.045 ;
        RECT  0.305 0.375 0.595 0.475 ;
        RECT  0.305 0.735 0.595 0.835 ;
        RECT  0.235 0.185 0.305 0.475 ;
        RECT  0.235 0.735 0.305 1.045 ;
        END
    END Z
    PIN NSLEEP
        ANTENNAGATEAREA 0.2436 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 1.905 3.195 1.975 ;
        RECT  1.995 1.565 2.065 1.975 ;
        RECT  1.565 1.565 1.995 1.635 ;
        RECT  1.495 1.565 1.565 1.835 ;
        RECT  1.230 1.765 1.495 1.835 ;
        RECT  1.110 1.765 1.230 1.905 ;
        END
    END NSLEEP
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.495 3.755 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 -0.115 5.180 0.115 ;
        RECT  4.690 -0.115 4.830 0.420 ;
        RECT  1.565 -0.115 4.690 0.115 ;
        RECT  1.495 -0.115 1.565 0.440 ;
        RECT  1.210 -0.115 1.495 0.115 ;
        RECT  1.130 -0.115 1.210 0.300 ;
        RECT  0.850 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.850 0.300 ;
        RECT  0.490 -0.115 0.770 0.115 ;
        RECT  0.410 -0.115 0.490 0.300 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.440 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        RECT  4.670 2.405 5.180 2.635 ;
        RECT  4.590 2.055 4.670 2.635 ;
        RECT  4.310 2.405 4.590 2.635 ;
        RECT  4.230 2.215 4.310 2.635 ;
        RECT  3.950 2.405 4.230 2.635 ;
        RECT  3.870 2.215 3.950 2.635 ;
        RECT  3.590 2.405 3.870 2.635 ;
        RECT  3.510 2.215 3.590 2.635 ;
        RECT  3.230 2.405 3.510 2.635 ;
        RECT  3.150 2.215 3.230 2.635 ;
        RECT  2.870 2.405 3.150 2.635 ;
        RECT  2.790 2.215 2.870 2.635 ;
        RECT  2.510 2.405 2.790 2.635 ;
        RECT  2.430 2.215 2.510 2.635 ;
        RECT  2.150 2.405 2.430 2.635 ;
        RECT  2.070 2.215 2.150 2.635 ;
        RECT  0.450 2.405 2.070 2.635 ;
        RECT  0.310 2.100 0.450 2.635 ;
        RECT  0.000 2.405 0.310 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.115 1.495 3.605 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.900 1.145 5.180 1.375 ;
        RECT  4.780 0.855 4.900 1.675 ;
        RECT  1.970 1.145 4.780 1.375 ;
        RECT  1.945 1.145 1.970 1.495 ;
        RECT  1.875 0.915 1.945 1.495 ;
        RECT  1.850 1.145 1.875 1.495 ;
        RECT  1.570 1.145 1.850 1.375 ;
        RECT  1.565 0.755 1.570 1.375 ;
        RECT  1.495 0.755 1.565 1.490 ;
        RECT  1.490 0.755 1.495 1.375 ;
        RECT  1.210 1.145 1.490 1.375 ;
        RECT  1.205 0.915 1.210 1.375 ;
        RECT  1.135 0.915 1.205 1.540 ;
        RECT  1.130 0.915 1.135 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.845 0.915 0.850 1.375 ;
        RECT  0.775 0.915 0.845 1.540 ;
        RECT  0.770 0.915 0.775 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.915 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.755 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.315 0.185 1.385 0.475 ;
        RECT  1.315 0.735 1.385 1.045 ;
        RECT  1.025 0.375 1.315 0.475 ;
        RECT  1.025 0.735 1.315 0.835 ;
        RECT  0.955 0.185 1.025 0.475 ;
        RECT  0.955 0.735 1.025 1.045 ;
        RECT  0.945 0.375 0.955 0.475 ;
        RECT  0.945 0.735 0.955 0.835 ;
        RECT  0.305 0.375 0.595 0.475 ;
        RECT  0.305 0.735 0.595 0.835 ;
        RECT  0.235 0.185 0.305 0.475 ;
        RECT  0.235 0.735 0.305 1.045 ;
        RECT  4.410 2.055 4.490 2.335 ;
        RECT  4.415 0.205 4.485 1.055 ;
        RECT  4.145 0.205 4.415 0.275 ;
        RECT  3.660 0.985 4.415 1.055 ;
        RECT  4.130 2.055 4.410 2.125 ;
        RECT  4.255 0.350 4.325 0.915 ;
        RECT  3.455 0.845 4.255 0.915 ;
        RECT  4.075 0.205 4.145 0.470 ;
        RECT  4.050 2.055 4.130 2.335 ;
        RECT  3.065 0.205 4.075 0.275 ;
        RECT  3.780 2.055 4.050 2.125 ;
        RECT  3.245 0.350 3.990 0.420 ;
        RECT  3.770 1.455 3.780 2.125 ;
        RECT  3.700 1.455 3.770 2.335 ;
        RECT  3.690 2.055 3.700 2.335 ;
        RECT  3.410 2.055 3.690 2.125 ;
        RECT  3.385 0.755 3.455 1.055 ;
        RECT  3.330 2.055 3.410 2.335 ;
        RECT  2.850 0.755 3.385 0.825 ;
        RECT  3.050 2.055 3.330 2.125 ;
        RECT  3.175 0.350 3.245 0.635 ;
        RECT  2.310 0.565 3.175 0.635 ;
        RECT  2.995 0.205 3.065 0.470 ;
        RECT  2.970 2.055 3.050 2.335 ;
        RECT  2.250 0.205 2.995 0.275 ;
        RECT  2.690 2.055 2.970 2.125 ;
        RECT  2.165 0.375 2.915 0.445 ;
        RECT  2.610 2.055 2.690 2.335 ;
        RECT  2.330 2.055 2.610 2.125 ;
        RECT  2.250 2.055 2.330 2.335 ;
        RECT  2.240 0.565 2.310 0.835 ;
        RECT  1.960 2.055 2.250 2.125 ;
        RECT  1.885 0.765 2.240 0.835 ;
        RECT  2.095 0.210 2.165 0.445 ;
        RECT  2.085 0.375 2.095 0.445 ;
        RECT  2.015 0.375 2.085 0.690 ;
        RECT  1.745 0.375 2.015 0.445 ;
        RECT  1.880 2.055 1.960 2.325 ;
        RECT  1.815 0.560 1.885 0.835 ;
        RECT  1.110 2.255 1.880 2.325 ;
        RECT  1.745 0.915 1.765 1.045 ;
        RECT  1.695 1.705 1.765 2.165 ;
        RECT  1.675 0.375 1.745 1.045 ;
        RECT  1.520 1.975 1.695 2.045 ;
        RECT  0.740 2.115 1.590 2.185 ;
        RECT  1.400 1.905 1.520 2.045 ;
        RECT  1.300 1.455 1.400 1.695 ;
        RECT  0.955 1.975 1.400 2.045 ;
        RECT  1.040 1.625 1.300 1.695 ;
        RECT  0.940 1.455 1.040 1.695 ;
        RECT  0.885 1.880 0.955 2.045 ;
        RECT  0.740 1.625 0.940 1.695 ;
        RECT  0.660 1.625 0.740 2.185 ;
        RECT  0.300 1.905 0.660 1.980 ;
    END
END LVLLHCLOD8BWP

MACRO LVLLHD1BWP
    CLASS CORE ;
    FOREIGN LVLLHD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 1.475 0.405 2.335 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.545 2.345 0.615 ;
        RECT  1.855 0.545 1.925 0.905 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 -0.115 3.500 0.115 ;
        RECT  2.990 -0.115 3.130 0.420 ;
        RECT  2.770 -0.115 2.990 0.115 ;
        RECT  2.690 -0.115 2.770 0.465 ;
        RECT  2.230 -0.115 2.690 0.115 ;
        RECT  2.150 -0.115 2.230 0.305 ;
        RECT  1.870 -0.115 2.150 0.115 ;
        RECT  1.790 -0.115 1.870 0.305 ;
        RECT  1.510 -0.115 1.790 0.115 ;
        RECT  1.430 -0.115 1.510 0.465 ;
        RECT  1.150 -0.115 1.430 0.115 ;
        RECT  1.070 -0.115 1.150 0.305 ;
        RECT  0.790 -0.115 1.070 0.115 ;
        RECT  0.710 -0.115 0.790 0.305 ;
        RECT  0.000 -0.115 0.710 0.115 ;
        RECT  3.130 2.405 3.500 2.635 ;
        RECT  2.990 2.100 3.130 2.635 ;
        RECT  0.585 2.405 2.990 2.635 ;
        RECT  0.515 2.055 0.585 2.635 ;
        RECT  0.000 2.405 0.515 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.495 2.205 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.145 3.500 1.375 ;
        RECT  3.105 0.855 3.225 1.675 ;
        RECT  0.590 1.145 3.105 1.375 ;
        RECT  0.585 0.915 0.590 1.375 ;
        RECT  0.515 0.915 0.585 1.760 ;
        RECT  0.510 0.915 0.515 1.375 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.510 0.185 2.590 0.840 ;
        RECT  2.100 0.760 2.510 0.840 ;
        RECT  2.335 0.185 2.405 0.465 ;
        RECT  2.045 0.395 2.335 0.465 ;
        RECT  2.020 0.760 2.100 1.055 ;
        RECT  1.975 0.185 2.045 0.465 ;
        RECT  1.460 0.985 2.020 1.055 ;
        RECT  1.685 0.395 1.975 0.465 ;
        RECT  1.615 0.185 1.685 0.635 ;
        RECT  0.955 0.565 1.615 0.635 ;
        RECT  1.380 0.730 1.460 1.055 ;
        RECT  1.255 0.185 1.325 0.465 ;
        RECT  0.965 0.395 1.255 0.465 ;
        RECT  0.895 0.185 0.965 0.465 ;
        RECT  0.885 0.565 0.955 0.835 ;
        RECT  0.715 0.395 0.895 0.465 ;
        RECT  0.525 0.765 0.885 0.835 ;
        RECT  0.645 0.395 0.715 0.690 ;
        RECT  0.375 0.395 0.645 0.465 ;
        RECT  0.455 0.560 0.525 0.835 ;
        RECT  0.375 0.915 0.405 1.045 ;
        RECT  0.305 0.395 0.375 1.045 ;
    END
END LVLLHD1BWP

MACRO LVLLHD2BWP
    CLASS CORE ;
    FOREIGN LVLLHD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 1.475 0.585 1.760 ;
        RECT  0.525 2.055 0.585 2.335 ;
        RECT  0.515 1.475 0.525 2.335 ;
        RECT  0.455 1.690 0.515 2.125 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.545 2.345 0.615 ;
        RECT  1.855 0.545 1.925 0.905 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 -0.115 3.500 0.115 ;
        RECT  2.990 -0.115 3.130 0.420 ;
        RECT  2.750 -0.115 2.990 0.115 ;
        RECT  2.670 -0.115 2.750 0.465 ;
        RECT  2.210 -0.115 2.670 0.115 ;
        RECT  2.130 -0.115 2.210 0.305 ;
        RECT  1.850 -0.115 2.130 0.115 ;
        RECT  1.770 -0.115 1.850 0.305 ;
        RECT  1.490 -0.115 1.770 0.115 ;
        RECT  1.410 -0.115 1.490 0.465 ;
        RECT  1.130 -0.115 1.410 0.115 ;
        RECT  1.050 -0.115 1.130 0.305 ;
        RECT  0.000 -0.115 1.050 0.115 ;
        RECT  3.130 2.405 3.500 2.635 ;
        RECT  2.990 2.100 3.130 2.635 ;
        RECT  0.770 2.405 2.990 2.635 ;
        RECT  0.690 2.055 0.770 2.635 ;
        RECT  0.410 2.405 0.690 2.635 ;
        RECT  0.330 2.210 0.410 2.635 ;
        RECT  0.000 2.405 0.330 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.495 2.205 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.145 3.500 1.375 ;
        RECT  3.105 0.855 3.225 1.675 ;
        RECT  0.800 1.145 3.105 1.375 ;
        RECT  0.770 0.970 0.800 1.375 ;
        RECT  0.720 0.970 0.770 1.770 ;
        RECT  0.690 1.145 0.720 1.770 ;
        RECT  0.590 1.145 0.690 1.375 ;
        RECT  0.510 0.915 0.590 1.375 ;
        RECT  0.410 1.145 0.510 1.375 ;
        RECT  0.330 1.145 0.410 1.570 ;
        RECT  0.000 1.145 0.330 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.185 2.570 0.840 ;
        RECT  2.100 0.760 2.490 0.840 ;
        RECT  2.315 0.185 2.385 0.465 ;
        RECT  2.025 0.395 2.315 0.465 ;
        RECT  2.020 0.760 2.100 1.055 ;
        RECT  1.955 0.185 2.025 0.465 ;
        RECT  1.440 0.985 2.020 1.055 ;
        RECT  1.665 0.395 1.955 0.465 ;
        RECT  1.595 0.185 1.665 0.635 ;
        RECT  0.955 0.565 1.595 0.635 ;
        RECT  1.360 0.730 1.440 1.055 ;
        RECT  1.235 0.185 1.305 0.465 ;
        RECT  0.945 0.395 1.235 0.465 ;
        RECT  0.885 0.565 0.955 0.835 ;
        RECT  0.870 0.185 0.945 0.465 ;
        RECT  0.525 0.765 0.885 0.835 ;
        RECT  0.725 0.395 0.870 0.465 ;
        RECT  0.655 0.395 0.725 0.690 ;
        RECT  0.375 0.395 0.655 0.465 ;
        RECT  0.455 0.560 0.525 0.835 ;
        RECT  0.375 0.915 0.405 1.045 ;
        RECT  0.305 0.395 0.375 1.045 ;
    END
END LVLLHD2BWP

MACRO LVLLHD4BWP
    CLASS CORE ;
    FOREIGN LVLLHD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 1.465 0.945 1.745 ;
        RECT  0.875 2.045 0.945 2.330 ;
        RECT  0.735 1.615 0.875 1.745 ;
        RECT  0.735 2.045 0.875 2.165 ;
        RECT  0.585 1.615 0.735 2.165 ;
        RECT  0.525 1.465 0.585 2.330 ;
        RECT  0.515 1.465 0.525 1.745 ;
        RECT  0.515 2.045 0.525 2.330 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0908 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.545 2.665 0.615 ;
        RECT  2.135 0.545 2.205 0.905 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.410 -0.115 3.780 0.115 ;
        RECT  3.270 -0.115 3.410 0.420 ;
        RECT  3.025 -0.115 3.270 0.115 ;
        RECT  2.955 -0.115 3.025 0.465 ;
        RECT  2.450 -0.115 2.955 0.115 ;
        RECT  2.370 -0.115 2.450 0.305 ;
        RECT  2.090 -0.115 2.370 0.115 ;
        RECT  2.010 -0.115 2.090 0.305 ;
        RECT  1.730 -0.115 2.010 0.115 ;
        RECT  1.650 -0.115 1.730 0.465 ;
        RECT  1.360 -0.115 1.650 0.115 ;
        RECT  1.280 -0.115 1.360 0.305 ;
        RECT  0.000 -0.115 1.280 0.115 ;
        RECT  3.410 2.405 3.780 2.635 ;
        RECT  3.270 2.100 3.410 2.635 ;
        RECT  1.130 2.405 3.270 2.635 ;
        RECT  1.050 2.055 1.130 2.635 ;
        RECT  0.790 2.405 1.050 2.635 ;
        RECT  0.670 2.245 0.790 2.635 ;
        RECT  0.410 2.405 0.670 2.635 ;
        RECT  0.330 2.055 0.410 2.635 ;
        RECT  0.000 2.405 0.330 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.995 1.495 2.485 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.145 3.780 1.375 ;
        RECT  3.380 0.855 3.500 1.675 ;
        RECT  1.130 1.145 3.380 1.375 ;
        RECT  1.050 1.145 1.130 1.755 ;
        RECT  0.790 1.145 1.050 1.375 ;
        RECT  0.670 1.145 0.790 1.535 ;
        RECT  0.590 1.145 0.670 1.375 ;
        RECT  0.510 0.915 0.590 1.375 ;
        RECT  0.410 1.145 0.510 1.375 ;
        RECT  0.330 1.145 0.410 1.755 ;
        RECT  0.000 1.145 0.330 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.875 1.465 0.945 1.745 ;
        RECT  0.875 2.045 0.945 2.330 ;
        RECT  0.805 1.615 0.875 1.745 ;
        RECT  0.805 2.045 0.875 2.165 ;
        RECT  2.770 0.185 2.850 0.840 ;
        RECT  2.380 0.760 2.770 0.840 ;
        RECT  2.555 0.185 2.625 0.465 ;
        RECT  2.265 0.395 2.555 0.465 ;
        RECT  2.300 0.760 2.380 1.055 ;
        RECT  1.675 0.985 2.300 1.055 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  1.905 0.395 2.195 0.465 ;
        RECT  1.835 0.185 1.905 0.635 ;
        RECT  1.440 0.565 1.835 0.635 ;
        RECT  1.605 0.730 1.675 1.055 ;
        RECT  1.475 0.185 1.545 0.465 ;
        RECT  1.165 0.395 1.475 0.465 ;
        RECT  1.360 0.565 1.440 1.065 ;
        RECT  1.360 1.455 1.440 1.975 ;
        RECT  0.525 0.765 1.360 0.835 ;
        RECT  0.890 1.905 1.360 1.975 ;
        RECT  1.095 0.185 1.165 0.465 ;
        RECT  0.725 0.395 1.095 0.465 ;
        RECT  0.655 0.395 0.725 0.690 ;
        RECT  0.375 0.395 0.655 0.465 ;
        RECT  0.455 0.560 0.525 0.835 ;
        RECT  0.375 0.915 0.405 1.045 ;
        RECT  0.305 0.395 0.375 1.045 ;
    END
END LVLLHD4BWP

MACRO LVLLHD8BWP
    CLASS CORE ;
    FOREIGN LVLLHD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE bcore ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.535 1.465 1.605 1.745 ;
        RECT  1.535 2.055 1.605 2.335 ;
        RECT  1.245 1.615 1.535 1.745 ;
        RECT  1.245 2.055 1.535 2.165 ;
        RECT  1.175 1.465 1.245 1.745 ;
        RECT  1.175 2.055 1.245 2.335 ;
        RECT  1.155 1.615 1.175 1.745 ;
        RECT  1.155 2.055 1.175 2.165 ;
        RECT  0.945 1.615 1.155 2.165 ;
        RECT  0.885 1.615 0.945 1.745 ;
        RECT  0.885 2.055 0.945 2.165 ;
        RECT  0.815 1.465 0.885 1.745 ;
        RECT  0.815 2.055 0.885 2.335 ;
        RECT  0.525 1.615 0.815 1.745 ;
        RECT  0.525 2.055 0.815 2.165 ;
        RECT  0.455 1.465 0.525 1.745 ;
        RECT  0.455 2.055 0.525 2.335 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1032 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.545 2.765 0.905 ;
        RECT  2.450 0.545 2.695 0.615 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.110 -0.115 4.480 0.115 ;
        RECT  3.970 -0.115 4.110 0.420 ;
        RECT  3.240 -0.115 3.970 0.115 ;
        RECT  3.160 -0.115 3.240 0.465 ;
        RECT  2.880 -0.115 3.160 0.115 ;
        RECT  2.800 -0.115 2.880 0.305 ;
        RECT  2.520 -0.115 2.800 0.115 ;
        RECT  2.440 -0.115 2.520 0.305 ;
        RECT  2.160 -0.115 2.440 0.115 ;
        RECT  2.080 -0.115 2.160 0.465 ;
        RECT  1.800 -0.115 2.080 0.115 ;
        RECT  1.720 -0.115 1.800 0.305 ;
        RECT  0.000 -0.115 1.720 0.115 ;
        RECT  4.110 2.405 4.480 2.635 ;
        RECT  3.970 2.100 4.110 2.635 ;
        RECT  1.790 2.405 3.970 2.635 ;
        RECT  1.710 2.055 1.790 2.635 ;
        RECT  1.450 2.405 1.710 2.635 ;
        RECT  1.330 2.245 1.450 2.635 ;
        RECT  1.090 2.405 1.330 2.635 ;
        RECT  0.970 2.245 1.090 2.635 ;
        RECT  0.730 2.405 0.970 2.635 ;
        RECT  0.610 2.245 0.730 2.635 ;
        RECT  0.350 2.405 0.610 2.635 ;
        RECT  0.270 2.055 0.350 2.635 ;
        RECT  0.000 2.405 0.270 2.635 ;
        END
    END VSS
    PIN VDDL
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.635 1.495 3.125 1.745 ;
        END
    END VDDL
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.145 4.480 1.375 ;
        RECT  4.080 0.855 4.200 1.675 ;
        RECT  1.790 1.145 4.080 1.375 ;
        RECT  1.710 1.145 1.790 1.745 ;
        RECT  1.450 1.145 1.710 1.375 ;
        RECT  1.330 1.145 1.450 1.535 ;
        RECT  1.090 1.145 1.330 1.375 ;
        RECT  0.970 1.145 1.090 1.535 ;
        RECT  0.730 1.145 0.970 1.375 ;
        RECT  0.610 1.145 0.730 1.535 ;
        RECT  0.530 1.145 0.610 1.375 ;
        RECT  0.450 0.915 0.530 1.375 ;
        RECT  0.350 1.145 0.450 1.375 ;
        RECT  0.270 1.145 0.350 1.745 ;
        RECT  0.000 1.145 0.270 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 1.465 1.605 1.745 ;
        RECT  1.535 2.055 1.605 2.335 ;
        RECT  1.245 1.615 1.535 1.745 ;
        RECT  1.245 2.055 1.535 2.165 ;
        RECT  1.225 1.465 1.245 1.745 ;
        RECT  1.225 2.055 1.245 2.335 ;
        RECT  0.815 1.465 0.875 1.745 ;
        RECT  0.815 2.055 0.875 2.335 ;
        RECT  0.525 1.615 0.815 1.745 ;
        RECT  0.525 2.055 0.815 2.165 ;
        RECT  0.455 1.465 0.525 1.745 ;
        RECT  0.455 2.055 0.525 2.335 ;
        RECT  3.340 0.185 3.420 0.840 ;
        RECT  3.055 0.760 3.340 0.840 ;
        RECT  2.985 0.185 3.055 0.465 ;
        RECT  2.985 0.760 3.055 1.055 ;
        RECT  2.695 0.395 2.985 0.465 ;
        RECT  2.285 0.985 2.985 1.055 ;
        RECT  2.625 0.185 2.695 0.465 ;
        RECT  2.335 0.395 2.625 0.465 ;
        RECT  2.265 0.185 2.335 0.635 ;
        RECT  2.215 0.755 2.285 1.055 ;
        RECT  1.865 0.565 2.265 0.635 ;
        RECT  2.010 0.755 2.215 0.825 ;
        RECT  1.865 0.970 2.110 1.040 ;
        RECT  2.000 1.455 2.080 1.975 ;
        RECT  1.270 1.905 2.000 1.975 ;
        RECT  1.905 0.185 1.975 0.465 ;
        RECT  1.615 0.395 1.905 0.465 ;
        RECT  1.795 0.565 1.865 1.040 ;
        RECT  0.465 0.765 1.795 0.835 ;
        RECT  1.545 0.185 1.615 0.465 ;
        RECT  0.655 0.395 1.545 0.465 ;
        RECT  0.460 1.900 0.780 1.980 ;
        RECT  0.585 0.395 0.655 0.690 ;
        RECT  0.325 0.395 0.585 0.465 ;
        RECT  0.395 0.560 0.465 0.835 ;
        RECT  0.325 0.915 0.345 1.045 ;
        RECT  0.255 0.395 0.325 1.045 ;
    END
END LVLLHD8BWP

MACRO MAOI222D0BWP
    CLASS CORE ;
    FOREIGN MAOI222D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1138 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.795 ;
        RECT  0.770 0.355 1.015 0.425 ;
        RECT  0.880 0.725 1.015 0.795 ;
        RECT  0.810 0.725 0.880 0.915 ;
        RECT  0.130 0.845 0.810 0.915 ;
        RECT  0.105 0.845 0.130 1.055 ;
        RECT  0.105 0.215 0.125 0.375 ;
        RECT  0.035 0.215 0.105 1.055 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.705 0.730 0.775 ;
        RECT  0.490 0.635 0.670 0.775 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.495 0.945 0.630 ;
        RECT  0.420 0.495 0.750 0.565 ;
        RECT  0.385 0.495 0.420 0.635 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.115 1.120 0.115 ;
        RECT  0.420 -0.115 0.520 0.415 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 1.120 1.375 ;
        RECT  0.430 0.985 0.510 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 0.185 1.080 0.285 ;
        RECT  0.990 0.895 1.070 1.055 ;
        RECT  0.590 0.985 0.990 1.055 ;
        RECT  0.690 0.205 0.980 0.275 ;
        RECT  0.610 0.205 0.690 0.425 ;
    END
END MAOI222D0BWP

MACRO MAOI222D1BWP
    CLASS CORE ;
    FOREIGN MAOI222D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1770 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.795 ;
        RECT  0.790 0.355 1.015 0.425 ;
        RECT  0.885 0.725 1.015 0.795 ;
        RECT  0.815 0.725 0.885 0.925 ;
        RECT  0.130 0.855 0.815 0.925 ;
        RECT  0.105 0.855 0.130 1.055 ;
        RECT  0.105 0.215 0.125 0.375 ;
        RECT  0.035 0.215 0.105 1.055 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.715 0.730 0.785 ;
        RECT  0.490 0.635 0.670 0.785 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0438 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.495 0.820 0.645 ;
        RECT  0.420 0.495 0.750 0.565 ;
        RECT  0.385 0.495 0.420 0.765 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.540 -0.115 1.120 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 1.120 1.375 ;
        RECT  0.430 0.995 0.510 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 0.185 1.080 0.285 ;
        RECT  0.990 0.895 1.070 1.065 ;
        RECT  0.590 0.995 0.990 1.065 ;
        RECT  0.710 0.205 0.980 0.275 ;
        RECT  0.630 0.205 0.710 0.425 ;
    END
END MAOI222D1BWP

MACRO MAOI222D2BWP
    CLASS CORE ;
    FOREIGN MAOI222D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.355 1.645 0.905 ;
        RECT  1.575 0.185 1.590 1.045 ;
        RECT  1.515 0.185 1.575 0.465 ;
        RECT  1.515 0.755 1.575 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.785 ;
        RECT  0.640 0.715 0.875 0.785 ;
        RECT  0.520 0.625 0.640 0.785 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.485 0.805 0.645 ;
        RECT  0.440 0.485 0.715 0.555 ;
        RECT  0.385 0.485 0.440 0.640 ;
        RECT  0.315 0.485 0.385 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.300 ;
        RECT  1.410 -0.115 1.690 0.115 ;
        RECT  1.330 -0.115 1.410 0.315 ;
        RECT  0.520 -0.115 1.330 0.115 ;
        RECT  0.420 -0.115 0.520 0.410 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.960 1.770 1.375 ;
        RECT  1.410 1.145 1.690 1.375 ;
        RECT  1.330 0.905 1.410 1.375 ;
        RECT  0.510 1.145 1.330 1.375 ;
        RECT  0.430 0.995 0.510 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.435 0.545 1.500 0.615 ;
        RECT  1.365 0.395 1.435 0.825 ;
        RECT  1.230 0.395 1.365 0.465 ;
        RECT  1.230 0.755 1.365 0.825 ;
        RECT  1.085 0.545 1.285 0.615 ;
        RECT  1.155 0.185 1.230 0.465 ;
        RECT  1.155 0.755 1.230 1.045 ;
        RECT  0.690 0.195 1.070 0.265 ;
        RECT  0.590 0.995 1.070 1.065 ;
        RECT  0.770 0.335 1.015 0.405 ;
        RECT  0.125 0.855 1.015 0.925 ;
        RECT  0.610 0.195 0.690 0.415 ;
        RECT  0.105 0.200 0.125 0.345 ;
        RECT  0.105 0.855 0.125 1.045 ;
        RECT  0.035 0.200 0.105 1.045 ;
        RECT  1.015 0.335 1.085 0.925 ;
    END
END MAOI222D2BWP

MACRO MAOI222D4BWP
    CLASS CORE ;
    FOREIGN MAOI222D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.005 0.465 ;
        RECT  1.995 0.775 2.005 1.055 ;
        RECT  1.935 0.185 1.995 1.055 ;
        RECT  1.785 0.355 1.935 0.905 ;
        RECT  1.605 0.355 1.785 0.465 ;
        RECT  1.605 0.775 1.785 0.905 ;
        RECT  1.535 0.185 1.605 0.465 ;
        RECT  1.535 0.775 1.605 1.055 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0218 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.945 0.785 ;
        RECT  0.640 0.715 0.870 0.785 ;
        RECT  0.520 0.625 0.640 0.785 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0454 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.485 0.790 0.645 ;
        RECT  0.440 0.485 0.720 0.555 ;
        RECT  0.385 0.485 0.440 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.485 ;
        RECT  1.810 -0.115 2.110 0.115 ;
        RECT  1.710 -0.115 1.810 0.275 ;
        RECT  1.430 -0.115 1.710 0.115 ;
        RECT  1.350 -0.115 1.430 0.295 ;
        RECT  0.540 -0.115 1.350 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.665 2.190 1.375 ;
        RECT  1.810 1.145 2.110 1.375 ;
        RECT  1.710 0.985 1.810 1.375 ;
        RECT  1.430 1.145 1.710 1.375 ;
        RECT  1.350 0.905 1.430 1.375 ;
        RECT  0.520 1.145 1.350 1.375 ;
        RECT  0.440 0.995 0.520 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.605 0.355 1.715 0.465 ;
        RECT  1.605 0.775 1.715 0.905 ;
        RECT  1.535 0.185 1.605 0.465 ;
        RECT  1.535 0.775 1.605 1.055 ;
        RECT  1.465 0.545 1.680 0.615 ;
        RECT  1.395 0.375 1.465 0.825 ;
        RECT  1.250 0.375 1.395 0.445 ;
        RECT  1.250 0.755 1.395 0.825 ;
        RECT  1.105 0.530 1.325 0.635 ;
        RECT  1.175 0.185 1.250 0.445 ;
        RECT  1.175 0.755 1.250 1.045 ;
        RECT  1.035 0.335 1.105 0.925 ;
        RECT  0.710 0.195 1.090 0.265 ;
        RECT  0.610 0.995 1.090 1.065 ;
        RECT  0.125 0.855 1.035 0.925 ;
        RECT  0.630 0.195 0.710 0.415 ;
        RECT  0.105 0.200 0.125 0.345 ;
        RECT  0.105 0.855 0.125 1.045 ;
        RECT  0.035 0.200 0.105 1.045 ;
        RECT  0.790 0.335 1.035 0.405 ;
    END
END MAOI222D4BWP

MACRO MAOI22D0BWP
    CLASS CORE ;
    FOREIGN MAOI22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0601 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.840 0.910 0.915 ;
        RECT  0.805 0.415 0.860 0.915 ;
        RECT  0.790 0.195 0.805 0.915 ;
        RECT  0.735 0.195 0.790 0.485 ;
        RECT  0.760 0.840 0.790 0.915 ;
        RECT  0.600 0.195 0.735 0.295 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0140 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0140 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.930 0.495 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0140 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.635 0.720 0.755 ;
        RECT  0.595 0.635 0.665 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.115 1.120 0.115 ;
        RECT  0.980 -0.115 1.080 0.275 ;
        RECT  0.130 -0.115 0.980 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.145 1.120 1.375 ;
        RECT  0.400 0.995 0.500 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.905 1.070 1.055 ;
        RECT  0.590 0.985 0.990 1.055 ;
        RECT  0.525 0.395 0.560 0.515 ;
        RECT  0.455 0.205 0.525 0.915 ;
        RECT  0.210 0.205 0.455 0.275 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.065 ;
    END
END MAOI22D0BWP

MACRO MAOI22D1BWP
    CLASS CORE ;
    FOREIGN MAOI22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1276 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.765 0.955 0.905 ;
        RECT  0.875 0.195 0.945 0.905 ;
        RECT  0.595 0.195 0.875 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.640 ;
        RECT  1.015 0.520 1.155 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.150 -0.115 1.260 0.115 ;
        RECT  1.070 -0.115 1.150 0.275 ;
        RECT  0.130 -0.115 1.070 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.145 1.260 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.075 0.765 1.145 1.055 ;
        RECT  0.640 0.985 1.075 1.055 ;
        RECT  0.525 0.520 0.600 0.640 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.210 0.215 0.455 0.285 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END MAOI22D1BWP

MACRO MAOI22D2BWP
    CLASS CORE ;
    FOREIGN MAOI22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.355 1.505 0.905 ;
        RECT  1.435 0.185 1.450 1.045 ;
        RECT  1.370 0.185 1.435 0.465 ;
        RECT  1.370 0.765 1.435 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.835 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.300 ;
        RECT  1.270 -0.115 1.550 0.115 ;
        RECT  1.190 -0.115 1.270 0.285 ;
        RECT  0.000 -0.115 1.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.960 1.630 1.375 ;
        RECT  1.200 1.145 1.550 1.375 ;
        RECT  1.200 0.985 1.290 1.055 ;
        RECT  1.080 0.985 1.200 1.375 ;
        RECT  0.990 0.985 1.080 1.055 ;
        RECT  0.540 1.145 1.080 1.375 ;
        RECT  0.420 0.995 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.290 0.540 1.350 0.620 ;
        RECT  1.220 0.355 1.290 0.915 ;
        RECT  0.790 0.355 1.220 0.425 ;
        RECT  0.610 0.845 1.220 0.915 ;
        RECT  0.620 0.205 1.110 0.275 ;
        RECT  0.525 0.545 0.640 0.615 ;
        RECT  0.455 0.205 0.525 0.915 ;
        RECT  0.130 0.205 0.455 0.275 ;
        RECT  0.210 0.845 0.455 0.915 ;
        RECT  0.050 0.205 0.130 0.345 ;
    END
END MAOI22D2BWP

MACRO MAOI22D4BWP
    CLASS CORE ;
    FOREIGN MAOI22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2304 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.865 0.465 ;
        RECT  1.855 0.775 1.865 1.055 ;
        RECT  1.795 0.185 1.855 1.055 ;
        RECT  1.645 0.355 1.795 0.905 ;
        RECT  1.465 0.355 1.645 0.465 ;
        RECT  1.465 0.775 1.645 0.905 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.835 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.470 ;
        RECT  1.670 -0.115 1.970 0.115 ;
        RECT  1.570 -0.115 1.670 0.275 ;
        RECT  1.270 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.270 0.285 ;
        RECT  0.000 -0.115 1.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.665 2.050 1.375 ;
        RECT  1.670 1.145 1.970 1.375 ;
        RECT  1.570 0.985 1.670 1.375 ;
        RECT  1.200 1.145 1.570 1.375 ;
        RECT  1.200 0.985 1.290 1.055 ;
        RECT  1.080 0.985 1.200 1.375 ;
        RECT  0.990 0.985 1.080 1.055 ;
        RECT  0.540 1.145 1.080 1.375 ;
        RECT  0.420 0.995 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.465 0.355 1.575 0.465 ;
        RECT  1.465 0.775 1.575 0.905 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        RECT  1.290 0.540 1.555 0.620 ;
        RECT  1.220 0.355 1.290 0.915 ;
        RECT  0.790 0.355 1.220 0.425 ;
        RECT  0.610 0.845 1.220 0.915 ;
        RECT  0.620 0.205 1.110 0.275 ;
        RECT  0.525 0.545 0.640 0.615 ;
        RECT  0.455 0.205 0.525 0.915 ;
        RECT  0.130 0.205 0.455 0.275 ;
        RECT  0.210 0.845 0.455 0.915 ;
        RECT  0.050 0.205 0.130 0.345 ;
    END
END MAOI22D4BWP

MACRO MOAI22D0BWP
    CLASS CORE ;
    FOREIGN MOAI22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0619 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.345 0.910 0.420 ;
        RECT  0.805 0.345 0.860 0.845 ;
        RECT  0.790 0.345 0.805 1.045 ;
        RECT  0.760 0.345 0.790 0.420 ;
        RECT  0.735 0.775 0.790 1.045 ;
        RECT  0.595 0.915 0.735 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.930 0.495 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.505 0.720 0.625 ;
        RECT  0.595 0.355 0.665 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.500 -0.115 1.120 0.115 ;
        RECT  0.400 -0.115 0.500 0.265 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.940 1.070 1.375 ;
        RECT  0.130 1.145 0.990 1.375 ;
        RECT  0.050 0.940 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.205 1.070 0.355 ;
        RECT  0.590 0.205 0.990 0.275 ;
        RECT  0.525 0.755 0.590 0.835 ;
        RECT  0.455 0.345 0.525 1.055 ;
        RECT  0.130 0.345 0.455 0.415 ;
        RECT  0.210 0.985 0.455 1.055 ;
        RECT  0.050 0.195 0.130 0.415 ;
    END
END MOAI22D0BWP

MACRO MOAI22D1BWP
    CLASS CORE ;
    FOREIGN MOAI22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1316 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.955 1.065 ;
        RECT  0.640 0.985 0.875 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.025 0.495 1.155 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.145 1.260 1.375 ;
        RECT  1.070 0.845 1.150 1.375 ;
        RECT  0.530 1.145 1.070 1.375 ;
        RECT  0.430 0.985 0.530 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.940 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.205 1.150 0.355 ;
        RECT  0.640 0.205 1.070 0.275 ;
        RECT  0.525 0.520 0.600 0.640 ;
        RECT  0.455 0.205 0.525 0.885 ;
        RECT  0.130 0.205 0.455 0.275 ;
        RECT  0.310 0.815 0.455 0.885 ;
        RECT  0.230 0.815 0.310 1.075 ;
        RECT  0.050 0.205 0.130 0.345 ;
    END
END MOAI22D1BWP

MACRO MOAI22D2BWP
    CLASS CORE ;
    FOREIGN MOAI22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.355 1.505 0.905 ;
        RECT  1.435 0.185 1.450 1.045 ;
        RECT  1.370 0.185 1.435 0.465 ;
        RECT  1.370 0.765 1.435 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.835 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.300 ;
        RECT  1.200 -0.115 1.550 0.115 ;
        RECT  1.200 0.205 1.290 0.275 ;
        RECT  1.080 -0.115 1.200 0.275 ;
        RECT  0.140 -0.115 1.080 0.115 ;
        RECT  0.990 0.205 1.080 0.275 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.960 1.630 1.375 ;
        RECT  1.270 1.145 1.550 1.375 ;
        RECT  1.190 0.975 1.270 1.375 ;
        RECT  0.530 1.145 1.190 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.290 0.540 1.350 0.620 ;
        RECT  1.220 0.345 1.290 0.905 ;
        RECT  0.750 0.345 1.220 0.415 ;
        RECT  0.790 0.835 1.220 0.905 ;
        RECT  0.610 0.985 1.110 1.055 ;
        RECT  0.630 0.205 0.750 0.415 ;
        RECT  0.525 0.545 0.640 0.615 ;
        RECT  0.455 0.205 0.525 0.915 ;
        RECT  0.210 0.205 0.455 0.275 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.025 ;
    END
END MOAI22D2BWP

MACRO MOAI22D4BWP
    CLASS CORE ;
    FOREIGN MOAI22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2304 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.865 0.465 ;
        RECT  1.855 0.775 1.865 1.055 ;
        RECT  1.795 0.185 1.855 1.055 ;
        RECT  1.645 0.355 1.795 0.905 ;
        RECT  1.465 0.355 1.645 0.465 ;
        RECT  1.465 0.775 1.645 0.905 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.835 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.470 ;
        RECT  1.670 -0.115 1.970 0.115 ;
        RECT  1.570 -0.115 1.670 0.275 ;
        RECT  1.200 -0.115 1.570 0.115 ;
        RECT  1.200 0.205 1.290 0.275 ;
        RECT  1.080 -0.115 1.200 0.275 ;
        RECT  0.140 -0.115 1.080 0.115 ;
        RECT  0.990 0.205 1.080 0.275 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.665 2.050 1.375 ;
        RECT  1.670 1.145 1.970 1.375 ;
        RECT  1.570 0.985 1.670 1.375 ;
        RECT  1.270 1.145 1.570 1.375 ;
        RECT  1.190 0.975 1.270 1.375 ;
        RECT  0.530 1.145 1.190 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.465 0.355 1.575 0.465 ;
        RECT  1.465 0.775 1.575 0.905 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        RECT  1.290 0.540 1.555 0.620 ;
        RECT  1.220 0.345 1.290 0.905 ;
        RECT  0.750 0.345 1.220 0.415 ;
        RECT  0.790 0.835 1.220 0.905 ;
        RECT  0.610 0.985 1.110 1.055 ;
        RECT  0.630 0.205 0.750 0.415 ;
        RECT  0.525 0.545 0.640 0.615 ;
        RECT  0.455 0.205 0.525 0.915 ;
        RECT  0.210 0.205 0.455 0.275 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.025 ;
    END
END MOAI22D4BWP

MACRO MUX2D0BWP
    CLASS CORE ;
    FOREIGN MUX2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.060 ;
        RECT  1.275 0.185 1.295 0.305 ;
        RECT  1.275 0.900 1.295 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.510 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.145 1.400 1.375 ;
        RECT  1.070 0.980 1.170 1.375 ;
        RECT  0.330 1.145 1.070 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.505 1.225 0.770 ;
        RECT  1.155 0.505 1.190 0.910 ;
        RECT  1.120 0.700 1.155 0.910 ;
        RECT  0.750 0.840 1.120 0.910 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.670 0.305 0.750 0.910 ;
        RECT  0.560 0.985 0.740 1.055 ;
        RECT  0.490 0.870 0.560 1.055 ;
        RECT  0.125 0.870 0.490 0.940 ;
        RECT  0.105 0.205 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.205 0.105 1.040 ;
    END
END MUX2D0BWP

MACRO MUX2D1BWP
    CLASS CORE ;
    FOREIGN MUX2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.060 ;
        RECT  1.275 0.185 1.295 0.465 ;
        RECT  1.275 0.900 1.295 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.510 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.420 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.145 1.400 1.375 ;
        RECT  1.070 0.990 1.170 1.375 ;
        RECT  0.330 1.145 1.070 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.515 1.225 0.770 ;
        RECT  1.155 0.515 1.190 0.920 ;
        RECT  1.120 0.700 1.155 0.920 ;
        RECT  0.760 0.850 1.120 0.920 ;
        RECT  0.900 0.195 1.000 0.275 ;
        RECT  0.900 0.710 1.000 0.780 ;
        RECT  0.830 0.195 0.900 0.780 ;
        RECT  0.740 0.995 0.900 1.075 ;
        RECT  0.660 0.335 0.760 0.920 ;
        RECT  0.560 0.995 0.740 1.065 ;
        RECT  0.490 0.315 0.560 0.790 ;
        RECT  0.490 0.870 0.560 1.065 ;
        RECT  0.125 0.870 0.490 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D1BWP

MACRO MUX2D2BWP
    CLASS CORE ;
    FOREIGN MUX2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.395 1.505 0.910 ;
        RECT  1.305 0.395 1.435 0.465 ;
        RECT  1.210 0.840 1.435 0.910 ;
        RECT  1.235 0.195 1.305 0.465 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.930 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.420 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.300 ;
        RECT  0.330 -0.115 1.410 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.990 1.500 1.375 ;
        RECT  1.130 1.145 1.400 1.375 ;
        RECT  1.050 0.990 1.130 1.375 ;
        RECT  0.330 1.145 1.050 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.545 1.310 0.615 ;
        RECT  1.155 0.545 1.225 0.770 ;
        RECT  1.120 0.700 1.155 0.770 ;
        RECT  1.050 0.700 1.120 0.920 ;
        RECT  0.710 0.850 1.050 0.920 ;
        RECT  0.850 0.710 0.970 0.780 ;
        RECT  0.850 0.225 0.920 0.345 ;
        RECT  0.720 0.995 0.880 1.075 ;
        RECT  0.780 0.225 0.850 0.780 ;
        RECT  0.490 0.995 0.720 1.065 ;
        RECT  0.640 0.315 0.710 0.920 ;
        RECT  0.490 0.315 0.560 0.780 ;
        RECT  0.460 0.315 0.490 0.455 ;
        RECT  0.390 0.710 0.490 0.780 ;
        RECT  0.420 0.850 0.490 1.065 ;
        RECT  0.125 0.850 0.420 0.920 ;
        RECT  0.105 0.195 0.125 0.315 ;
        RECT  0.105 0.850 0.125 1.020 ;
        RECT  0.035 0.195 0.105 1.020 ;
    END
END MUX2D2BWP

MACRO MUX2D4BWP
    CLASS CORE ;
    FOREIGN MUX2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.185 2.145 0.465 ;
        RECT  2.135 0.775 2.145 1.055 ;
        RECT  2.075 0.185 2.135 1.055 ;
        RECT  1.925 0.355 2.075 0.905 ;
        RECT  1.785 0.355 1.925 0.465 ;
        RECT  1.785 0.775 1.925 0.905 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.715 0.775 1.785 1.055 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.0342 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.640 ;
        RECT  1.090 0.520 1.155 0.640 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.350 1.505 0.670 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.495 0.385 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.485 ;
        RECT  1.990 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.990 0.270 ;
        RECT  1.620 -0.115 1.870 0.115 ;
        RECT  1.520 -0.115 1.620 0.270 ;
        RECT  0.320 -0.115 1.520 0.115 ;
        RECT  0.220 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.145 2.380 1.375 ;
        RECT  2.250 0.680 2.330 1.375 ;
        RECT  1.980 1.145 2.250 1.375 ;
        RECT  1.880 0.985 1.980 1.375 ;
        RECT  1.630 1.145 1.880 1.375 ;
        RECT  1.510 1.030 1.630 1.375 ;
        RECT  1.270 1.145 1.510 1.375 ;
        RECT  1.150 1.030 1.270 1.375 ;
        RECT  0.310 1.145 1.150 1.375 ;
        RECT  0.230 0.980 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.355 1.855 0.465 ;
        RECT  1.785 0.775 1.855 0.905 ;
        RECT  1.715 0.185 1.785 0.465 ;
        RECT  1.715 0.775 1.785 1.055 ;
        RECT  1.645 0.545 1.820 0.615 ;
        RECT  1.575 0.545 1.645 0.960 ;
        RECT  0.675 0.890 1.575 0.960 ;
        RECT  1.365 0.750 1.470 0.820 ;
        RECT  1.365 0.195 1.450 0.265 ;
        RECT  1.295 0.195 1.365 0.820 ;
        RECT  0.815 0.205 1.295 0.275 ;
        RECT  1.010 0.750 1.090 0.820 ;
        RECT  1.010 0.350 1.060 0.450 ;
        RECT  0.940 0.350 1.010 0.820 ;
        RECT  0.890 0.500 0.940 0.620 ;
        RECT  0.815 0.690 0.865 0.810 ;
        RECT  0.745 0.205 0.815 0.810 ;
        RECT  0.605 0.240 0.675 0.960 ;
        RECT  0.415 0.240 0.485 0.415 ;
        RECT  0.415 0.840 0.485 1.045 ;
        RECT  0.125 0.345 0.415 0.415 ;
        RECT  0.125 0.840 0.415 0.910 ;
        RECT  0.055 0.230 0.125 1.070 ;
    END
END MUX2D4BWP

MACRO MUX2ND0BWP
    CLASS CORE ;
    FOREIGN MUX2ND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0796 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.215 0.735 0.295 ;
        RECT  0.665 0.825 0.720 0.925 ;
        RECT  0.595 0.215 0.665 0.485 ;
        RECT  0.595 0.705 0.665 0.925 ;
        RECT  0.580 0.405 0.595 0.485 ;
        RECT  0.580 0.705 0.595 0.775 ;
        RECT  0.510 0.405 0.580 0.775 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.470 0.245 0.785 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.930 0.495 1.015 0.640 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.440 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.115 1.120 0.115 ;
        RECT  0.990 -0.115 1.070 0.410 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.860 1.070 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 1.005 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.790 0.555 0.860 1.065 ;
        RECT  0.660 0.555 0.790 0.635 ;
        RECT  0.480 0.995 0.790 1.065 ;
        RECT  0.410 0.865 0.480 1.065 ;
        RECT  0.130 0.865 0.410 0.935 ;
        RECT  0.105 0.865 0.130 1.055 ;
        RECT  0.105 0.285 0.120 0.425 ;
        RECT  0.035 0.285 0.105 1.055 ;
    END
END MUX2ND0BWP

MACRO MUX2ND1BWP
    CLASS CORE ;
    FOREIGN MUX2ND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.185 1.785 1.070 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.625 ;
        RECT  0.970 0.520 1.015 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.420 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.590 -0.115 1.820 0.115 ;
        RECT  1.510 -0.115 1.590 0.315 ;
        RECT  1.210 -0.115 1.510 0.115 ;
        RECT  1.110 -0.115 1.210 0.275 ;
        RECT  0.360 -0.115 1.110 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.585 1.145 1.820 1.375 ;
        RECT  1.515 0.925 1.585 1.375 ;
        RECT  1.200 1.145 1.515 1.375 ;
        RECT  1.120 0.980 1.200 1.375 ;
        RECT  0.330 1.145 1.120 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.545 0.395 1.615 0.845 ;
        RECT  1.405 0.395 1.545 0.465 ;
        RECT  1.405 0.775 1.545 0.845 ;
        RECT  1.335 0.185 1.405 0.465 ;
        RECT  1.335 0.775 1.405 1.055 ;
        RECT  1.225 0.545 1.340 0.620 ;
        RECT  1.155 0.545 1.225 0.910 ;
        RECT  0.750 0.840 1.155 0.910 ;
        RECT  0.900 0.700 1.030 0.770 ;
        RECT  0.900 0.205 1.020 0.275 ;
        RECT  0.760 0.995 0.920 1.075 ;
        RECT  0.830 0.205 0.900 0.770 ;
        RECT  0.560 0.995 0.760 1.065 ;
        RECT  0.670 0.325 0.750 0.910 ;
        RECT  0.510 0.335 0.580 0.770 ;
        RECT  0.490 0.850 0.560 1.065 ;
        RECT  0.480 0.335 0.510 0.455 ;
        RECT  0.460 0.700 0.510 0.770 ;
        RECT  0.125 0.850 0.490 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND1BWP

MACRO MUX2ND2BWP
    CLASS CORE ;
    FOREIGN MUX2ND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.355 1.785 0.905 ;
        RECT  1.715 0.185 1.730 1.055 ;
        RECT  1.650 0.185 1.715 0.465 ;
        RECT  1.650 0.795 1.715 1.055 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.625 ;
        RECT  0.970 0.520 1.015 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.420 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.830 -0.115 1.910 0.300 ;
        RECT  1.550 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.550 0.315 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.360 -0.115 1.090 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.830 0.960 1.910 1.375 ;
        RECT  1.550 1.145 1.830 1.375 ;
        RECT  1.470 0.915 1.550 1.375 ;
        RECT  1.180 1.145 1.470 1.375 ;
        RECT  1.100 0.980 1.180 1.375 ;
        RECT  0.330 1.145 1.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.395 1.575 0.805 ;
        RECT  1.370 0.395 1.505 0.465 ;
        RECT  1.370 0.735 1.505 0.805 ;
        RECT  1.290 0.185 1.370 0.465 ;
        RECT  1.295 0.735 1.370 1.055 ;
        RECT  1.225 0.545 1.290 0.615 ;
        RECT  1.155 0.545 1.225 0.910 ;
        RECT  0.750 0.840 1.155 0.910 ;
        RECT  0.900 0.700 1.030 0.770 ;
        RECT  0.900 0.205 1.020 0.275 ;
        RECT  0.760 0.995 0.920 1.075 ;
        RECT  0.830 0.205 0.900 0.770 ;
        RECT  0.560 0.995 0.760 1.065 ;
        RECT  0.670 0.325 0.750 0.910 ;
        RECT  0.510 0.335 0.580 0.770 ;
        RECT  0.490 0.850 0.560 1.065 ;
        RECT  0.480 0.335 0.510 0.455 ;
        RECT  0.460 0.700 0.510 0.770 ;
        RECT  0.125 0.850 0.490 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND2BWP

MACRO MUX2ND4BWP
    CLASS CORE ;
    FOREIGN MUX2ND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.565 0.465 ;
        RECT  2.555 0.775 2.565 1.055 ;
        RECT  2.495 0.185 2.555 1.055 ;
        RECT  2.345 0.355 2.495 0.905 ;
        RECT  2.205 0.355 2.345 0.465 ;
        RECT  2.205 0.775 2.345 0.905 ;
        RECT  2.135 0.185 2.205 0.465 ;
        RECT  2.135 0.775 2.205 1.055 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.0342 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.090 0.495 1.155 0.640 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.350 1.505 0.670 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.495 0.385 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.485 ;
        RECT  2.410 -0.115 2.670 0.115 ;
        RECT  2.290 -0.115 2.410 0.270 ;
        RECT  2.030 -0.115 2.290 0.115 ;
        RECT  1.950 -0.115 2.030 0.305 ;
        RECT  1.650 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.650 0.270 ;
        RECT  0.320 -0.115 1.550 0.115 ;
        RECT  0.220 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.680 2.750 1.375 ;
        RECT  2.400 1.145 2.670 1.375 ;
        RECT  2.300 0.985 2.400 1.375 ;
        RECT  2.030 1.145 2.300 1.375 ;
        RECT  1.950 0.850 2.030 1.375 ;
        RECT  1.660 1.145 1.950 1.375 ;
        RECT  1.540 1.030 1.660 1.375 ;
        RECT  1.270 1.145 1.540 1.375 ;
        RECT  1.150 1.030 1.270 1.375 ;
        RECT  0.310 1.145 1.150 1.375 ;
        RECT  0.230 0.980 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.355 2.275 0.465 ;
        RECT  2.205 0.775 2.275 0.905 ;
        RECT  2.135 0.185 2.205 0.465 ;
        RECT  2.135 0.775 2.205 1.055 ;
        RECT  2.060 0.545 2.240 0.615 ;
        RECT  1.980 0.395 2.060 0.770 ;
        RECT  1.850 0.395 1.980 0.465 ;
        RECT  1.850 0.700 1.980 0.770 ;
        RECT  1.655 0.545 1.890 0.615 ;
        RECT  1.770 0.185 1.850 0.465 ;
        RECT  1.770 0.700 1.850 1.020 ;
        RECT  1.585 0.545 1.655 0.960 ;
        RECT  0.675 0.890 1.585 0.960 ;
        RECT  1.365 0.750 1.470 0.820 ;
        RECT  1.365 0.195 1.450 0.265 ;
        RECT  1.295 0.195 1.365 0.820 ;
        RECT  0.815 0.205 1.295 0.275 ;
        RECT  1.010 0.350 1.070 0.420 ;
        RECT  1.010 0.750 1.070 0.820 ;
        RECT  0.940 0.350 1.010 0.820 ;
        RECT  0.890 0.500 0.940 0.620 ;
        RECT  0.815 0.690 0.865 0.810 ;
        RECT  0.745 0.205 0.815 0.810 ;
        RECT  0.605 0.240 0.675 0.960 ;
        RECT  0.415 0.240 0.485 0.415 ;
        RECT  0.415 0.840 0.485 1.045 ;
        RECT  0.125 0.345 0.415 0.415 ;
        RECT  0.125 0.840 0.415 0.910 ;
        RECT  0.055 0.195 0.125 1.070 ;
    END
END MUX2ND4BWP

MACRO MUX3D0BWP
    CLASS CORE ;
    FOREIGN MUX3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.215 2.345 1.070 ;
        RECT  2.255 0.215 2.275 0.425 ;
        RECT  2.240 0.970 2.275 1.070 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.250 0.650 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.775 2.205 0.905 ;
        RECT  1.930 0.500 2.000 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0146 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.625 ;
        RECT  0.990 0.500 1.015 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 2.380 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.145 2.380 1.375 ;
        RECT  2.020 0.985 2.140 1.375 ;
        RECT  0.330 1.145 2.020 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.175 0.520 2.195 0.640 ;
        RECT  2.105 0.205 2.175 0.640 ;
        RECT  1.720 0.205 2.105 0.275 ;
        RECT  1.860 0.350 1.950 0.420 ;
        RECT  1.860 0.985 1.950 1.065 ;
        RECT  1.790 0.350 1.860 1.065 ;
        RECT  1.650 0.205 1.720 1.045 ;
        RECT  1.510 0.320 1.580 1.045 ;
        RECT  1.460 0.320 1.510 0.480 ;
        RECT  1.085 0.975 1.510 1.045 ;
        RECT  1.390 0.570 1.440 0.690 ;
        RECT  1.320 0.230 1.390 0.905 ;
        RECT  1.250 0.230 1.320 0.300 ;
        RECT  1.250 0.835 1.320 0.905 ;
        RECT  1.005 0.845 1.085 1.045 ;
        RECT  0.910 0.705 1.020 0.775 ;
        RECT  0.745 0.845 1.005 0.915 ;
        RECT  0.910 0.195 0.975 0.275 ;
        RECT  0.800 0.985 0.920 1.075 ;
        RECT  0.840 0.195 0.910 0.775 ;
        RECT  0.560 0.985 0.800 1.055 ;
        RECT  0.675 0.325 0.745 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.490 0.850 0.560 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.490 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D0BWP

MACRO MUX3D1BWP
    CLASS CORE ;
    FOREIGN MUX3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.195 2.345 1.070 ;
        RECT  2.255 0.195 2.275 0.475 ;
        RECT  2.240 0.970 2.275 1.070 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.250 0.650 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.775 2.205 0.905 ;
        RECT  1.930 0.500 2.000 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 2.380 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 2.380 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.175 0.520 2.195 0.640 ;
        RECT  2.105 0.205 2.175 0.640 ;
        RECT  1.720 0.205 2.105 0.275 ;
        RECT  1.860 0.350 1.950 0.420 ;
        RECT  1.860 0.985 1.950 1.065 ;
        RECT  1.790 0.350 1.860 1.065 ;
        RECT  1.650 0.205 1.720 1.045 ;
        RECT  1.510 0.320 1.580 1.045 ;
        RECT  1.460 0.320 1.510 0.480 ;
        RECT  1.085 0.975 1.510 1.045 ;
        RECT  1.390 0.570 1.440 0.690 ;
        RECT  1.320 0.225 1.390 0.905 ;
        RECT  1.250 0.225 1.320 0.295 ;
        RECT  1.230 0.835 1.320 0.905 ;
        RECT  1.005 0.845 1.085 1.045 ;
        RECT  0.750 0.845 1.005 0.915 ;
        RECT  0.890 0.705 0.990 0.775 ;
        RECT  0.890 0.195 0.975 0.275 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.820 0.195 0.890 0.775 ;
        RECT  0.670 0.325 0.750 0.915 ;
        RECT  0.530 0.985 0.740 1.055 ;
        RECT  0.630 0.835 0.670 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.460 0.850 0.530 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.460 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D1BWP

MACRO MUX3D2BWP
    CLASS CORE ;
    FOREIGN MUX3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.355 2.345 0.905 ;
        RECT  2.275 0.185 2.290 1.055 ;
        RECT  2.220 0.185 2.275 0.465 ;
        RECT  2.210 0.795 2.275 1.055 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.250 0.650 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.775 2.080 1.045 ;
        RECT  1.990 0.500 2.000 1.045 ;
        RECT  1.930 0.500 1.990 0.885 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.300 ;
        RECT  1.170 -0.115 2.390 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.960 2.470 1.375 ;
        RECT  0.330 1.145 2.390 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.140 0.530 2.190 0.630 ;
        RECT  2.070 0.210 2.140 0.630 ;
        RECT  1.720 0.210 2.070 0.280 ;
        RECT  1.860 0.350 1.950 0.420 ;
        RECT  1.860 0.965 1.920 1.065 ;
        RECT  1.790 0.350 1.860 1.065 ;
        RECT  1.650 0.210 1.720 1.045 ;
        RECT  1.510 0.320 1.580 1.045 ;
        RECT  1.460 0.320 1.510 0.480 ;
        RECT  1.085 0.975 1.510 1.045 ;
        RECT  1.390 0.590 1.440 0.710 ;
        RECT  1.320 0.225 1.390 0.905 ;
        RECT  1.250 0.225 1.320 0.295 ;
        RECT  1.230 0.835 1.320 0.905 ;
        RECT  1.005 0.845 1.085 1.045 ;
        RECT  0.750 0.845 1.005 0.915 ;
        RECT  0.890 0.705 0.990 0.775 ;
        RECT  0.890 0.195 0.975 0.275 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.820 0.195 0.890 0.775 ;
        RECT  0.670 0.325 0.750 0.915 ;
        RECT  0.530 0.985 0.740 1.055 ;
        RECT  0.630 0.835 0.670 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.460 0.850 0.530 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.460 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D2BWP

MACRO MUX3D4BWP
    CLASS CORE ;
    FOREIGN MUX3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.185 3.405 0.465 ;
        RECT  3.395 0.775 3.405 1.055 ;
        RECT  3.335 0.185 3.395 1.055 ;
        RECT  3.185 0.355 3.335 0.905 ;
        RECT  3.045 0.355 3.185 0.465 ;
        RECT  3.045 0.775 3.185 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.405 0.355 2.485 0.640 ;
        RECT  2.370 0.520 2.405 0.640 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.640 ;
        RECT  1.090 0.520 1.155 0.640 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.350 2.765 0.670 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.525 0.640 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.495 0.385 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.640 0.115 ;
        RECT  3.510 -0.115 3.590 0.485 ;
        RECT  3.250 -0.115 3.510 0.115 ;
        RECT  3.130 -0.115 3.250 0.270 ;
        RECT  2.880 -0.115 3.130 0.115 ;
        RECT  2.780 -0.115 2.880 0.270 ;
        RECT  1.600 -0.115 2.780 0.115 ;
        RECT  1.500 -0.115 1.600 0.285 ;
        RECT  0.320 -0.115 1.500 0.115 ;
        RECT  0.220 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.665 3.590 1.375 ;
        RECT  3.240 1.145 3.510 1.375 ;
        RECT  3.140 0.985 3.240 1.375 ;
        RECT  2.890 1.145 3.140 1.375 ;
        RECT  2.770 1.030 2.890 1.375 ;
        RECT  0.310 1.145 2.770 1.375 ;
        RECT  0.230 0.980 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.355 3.115 0.465 ;
        RECT  3.045 0.775 3.115 0.905 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.775 3.045 1.055 ;
        RECT  2.905 0.545 3.080 0.615 ;
        RECT  2.835 0.545 2.905 0.960 ;
        RECT  1.950 0.890 2.835 0.960 ;
        RECT  2.625 0.750 2.730 0.820 ;
        RECT  2.625 0.195 2.710 0.265 ;
        RECT  2.555 0.195 2.625 0.820 ;
        RECT  2.100 0.205 2.555 0.275 ;
        RECT  2.300 0.730 2.370 0.810 ;
        RECT  2.300 0.345 2.325 0.465 ;
        RECT  2.230 0.345 2.300 0.810 ;
        RECT  2.180 0.500 2.230 0.640 ;
        RECT  2.100 0.710 2.160 0.810 ;
        RECT  2.030 0.205 2.100 0.810 ;
        RECT  1.870 0.195 1.950 0.960 ;
        RECT  1.690 0.195 1.770 1.065 ;
        RECT  0.670 0.995 1.690 1.065 ;
        RECT  1.225 0.855 1.610 0.925 ;
        RECT  1.365 0.715 1.450 0.785 ;
        RECT  1.365 0.185 1.420 0.285 ;
        RECT  1.305 0.185 1.365 0.785 ;
        RECT  1.295 0.205 1.305 0.785 ;
        RECT  0.820 0.205 1.295 0.275 ;
        RECT  1.150 0.745 1.225 0.925 ;
        RECT  1.020 0.350 1.070 0.450 ;
        RECT  1.020 0.775 1.070 0.855 ;
        RECT  0.950 0.350 1.020 0.855 ;
        RECT  0.900 0.520 0.950 0.640 ;
        RECT  0.820 0.755 0.870 0.875 ;
        RECT  0.750 0.205 0.820 0.875 ;
        RECT  0.590 0.230 0.670 1.065 ;
        RECT  0.410 0.230 0.490 0.415 ;
        RECT  0.410 0.840 0.490 1.025 ;
        RECT  0.125 0.345 0.410 0.415 ;
        RECT  0.125 0.840 0.410 0.910 ;
        RECT  0.055 0.195 0.125 1.070 ;
    END
END MUX3D4BWP

MACRO MUX3ND0BWP
    CLASS CORE ;
    FOREIGN MUX3ND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0945 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.215 1.790 1.065 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.445 1.245 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.205 0.765 ;
        RECT  2.040 0.495 2.135 0.645 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.965 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.420 ;
        RECT  0.360 -0.115 2.110 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.200 1.145 2.240 1.375 ;
        RECT  2.100 0.850 2.200 1.375 ;
        RECT  0.330 1.145 2.100 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 0.185 1.985 0.445 ;
        RECT  1.940 0.735 1.985 1.035 ;
        RECT  1.915 0.185 1.940 1.035 ;
        RECT  1.870 0.375 1.915 0.805 ;
        RECT  1.520 0.285 1.590 1.055 ;
        RECT  1.495 0.285 1.520 0.435 ;
        RECT  1.085 0.985 1.520 1.055 ;
        RECT  1.390 0.510 1.450 0.630 ;
        RECT  1.315 0.195 1.390 0.855 ;
        RECT  1.005 0.845 1.085 1.055 ;
        RECT  0.750 0.845 1.005 0.915 ;
        RECT  0.890 0.195 0.995 0.275 ;
        RECT  0.890 0.705 0.990 0.775 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.820 0.195 0.890 0.775 ;
        RECT  0.670 0.325 0.750 0.915 ;
        RECT  0.530 0.985 0.740 1.055 ;
        RECT  0.630 0.835 0.670 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.460 0.850 0.530 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.460 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND0BWP

MACRO MUX3ND1BWP
    CLASS CORE ;
    FOREIGN MUX3ND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.185 2.625 1.070 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0328 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.065 0.640 ;
        RECT  1.930 0.520 1.995 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.965 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.115 2.660 0.115 ;
        RECT  2.350 -0.115 2.430 0.300 ;
        RECT  2.080 -0.115 2.350 0.115 ;
        RECT  1.980 -0.115 2.080 0.275 ;
        RECT  1.160 -0.115 1.980 0.115 ;
        RECT  1.060 -0.115 1.160 0.275 ;
        RECT  0.360 -0.115 1.060 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.145 2.660 1.375 ;
        RECT  2.330 1.005 2.450 1.375 ;
        RECT  2.090 1.145 2.330 1.375 ;
        RECT  1.970 1.030 2.090 1.375 ;
        RECT  0.330 1.145 1.970 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.380 2.465 0.930 ;
        RECT  2.250 0.380 2.390 0.450 ;
        RECT  2.245 0.860 2.390 0.930 ;
        RECT  2.150 0.190 2.250 0.450 ;
        RECT  2.175 0.860 2.245 1.020 ;
        RECT  2.145 0.520 2.215 0.780 ;
        RECT  2.100 0.710 2.145 0.780 ;
        RECT  2.030 0.710 2.100 0.960 ;
        RECT  1.720 0.890 2.030 0.960 ;
        RECT  1.860 0.750 1.930 0.820 ;
        RECT  1.860 0.280 1.900 0.380 ;
        RECT  1.790 0.280 1.860 0.820 ;
        RECT  1.640 0.285 1.720 1.045 ;
        RECT  1.500 0.320 1.570 1.045 ;
        RECT  1.440 0.320 1.500 0.480 ;
        RECT  1.085 0.975 1.500 1.045 ;
        RECT  1.370 0.570 1.430 0.690 ;
        RECT  1.300 0.205 1.370 0.905 ;
        RECT  1.230 0.205 1.300 0.275 ;
        RECT  1.250 0.835 1.300 0.905 ;
        RECT  1.005 0.845 1.085 1.045 ;
        RECT  0.750 0.845 1.005 0.915 ;
        RECT  0.890 0.705 0.990 0.775 ;
        RECT  0.890 0.195 0.975 0.275 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.820 0.195 0.890 0.775 ;
        RECT  0.670 0.325 0.750 0.915 ;
        RECT  0.530 0.985 0.740 1.055 ;
        RECT  0.630 0.835 0.670 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.460 0.850 0.530 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.460 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND1BWP

MACRO MUX3ND2BWP
    CLASS CORE ;
    FOREIGN MUX3ND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.710 0.355 2.765 0.905 ;
        RECT  2.705 0.185 2.710 0.905 ;
        RECT  2.695 0.185 2.705 1.055 ;
        RECT  2.635 0.185 2.695 0.485 ;
        RECT  2.635 0.795 2.695 1.055 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.250 0.650 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.065 0.640 ;
        RECT  1.950 0.530 1.995 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.530 1.015 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0174 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.480 0.430 0.630 ;
        RECT  0.315 0.355 0.385 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.300 ;
        RECT  2.530 -0.115 2.810 0.115 ;
        RECT  2.450 -0.115 2.530 0.315 ;
        RECT  1.170 -0.115 2.450 0.115 ;
        RECT  1.070 -0.115 1.170 0.275 ;
        RECT  0.360 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.960 2.890 1.375 ;
        RECT  2.530 1.145 2.810 1.375 ;
        RECT  2.450 0.915 2.530 1.375 ;
        RECT  2.130 1.145 2.450 1.375 ;
        RECT  2.050 0.745 2.130 1.375 ;
        RECT  0.330 1.145 2.050 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.395 2.565 0.805 ;
        RECT  2.365 0.395 2.490 0.465 ;
        RECT  2.350 0.735 2.490 0.805 ;
        RECT  2.275 0.185 2.365 0.465 ;
        RECT  2.270 0.735 2.350 1.055 ;
        RECT  2.205 0.540 2.320 0.620 ;
        RECT  2.135 0.195 2.205 0.620 ;
        RECT  1.720 0.195 2.135 0.265 ;
        RECT  1.860 0.345 1.920 0.445 ;
        RECT  1.860 0.745 1.905 1.065 ;
        RECT  1.835 0.345 1.860 1.065 ;
        RECT  1.790 0.345 1.835 0.815 ;
        RECT  1.650 0.195 1.720 1.065 ;
        RECT  1.510 0.330 1.580 1.045 ;
        RECT  1.460 0.330 1.510 0.480 ;
        RECT  1.085 0.975 1.510 1.045 ;
        RECT  1.390 0.570 1.440 0.690 ;
        RECT  1.320 0.220 1.390 0.905 ;
        RECT  1.250 0.220 1.320 0.290 ;
        RECT  1.230 0.835 1.320 0.905 ;
        RECT  1.005 0.845 1.085 1.045 ;
        RECT  0.750 0.845 1.005 0.915 ;
        RECT  0.890 0.705 0.990 0.775 ;
        RECT  0.890 0.195 0.975 0.275 ;
        RECT  0.740 0.985 0.900 1.075 ;
        RECT  0.820 0.195 0.890 0.775 ;
        RECT  0.670 0.325 0.750 0.915 ;
        RECT  0.530 0.985 0.740 1.055 ;
        RECT  0.630 0.835 0.670 0.915 ;
        RECT  0.500 0.325 0.580 0.770 ;
        RECT  0.460 0.850 0.530 1.055 ;
        RECT  0.460 0.700 0.500 0.770 ;
        RECT  0.125 0.850 0.460 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND2BWP

MACRO MUX3ND4BWP
    CLASS CORE ;
    FOREIGN MUX3ND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.710 3.460 0.800 ;
        RECT  3.395 0.185 3.425 0.465 ;
        RECT  3.350 0.185 3.395 0.800 ;
        RECT  3.185 0.355 3.350 0.800 ;
        RECT  3.070 0.355 3.185 0.485 ;
        RECT  2.970 0.710 3.185 0.800 ;
        RECT  2.990 0.185 3.070 0.485 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.405 0.355 2.485 0.640 ;
        RECT  2.370 0.520 2.405 0.640 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.640 ;
        RECT  1.090 0.520 1.155 0.640 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.350 2.785 0.670 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.525 0.640 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.495 0.385 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.670 -0.115 3.920 0.115 ;
        RECT  3.570 -0.115 3.670 0.290 ;
        RECT  3.260 -0.115 3.570 0.115 ;
        RECT  3.160 -0.115 3.260 0.275 ;
        RECT  2.890 -0.115 3.160 0.115 ;
        RECT  2.790 -0.115 2.890 0.275 ;
        RECT  1.600 -0.115 2.790 0.115 ;
        RECT  1.500 -0.115 1.600 0.285 ;
        RECT  0.320 -0.115 1.500 0.115 ;
        RECT  0.220 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.680 1.145 3.920 1.375 ;
        RECT  3.560 1.020 3.680 1.375 ;
        RECT  3.270 1.145 3.560 1.375 ;
        RECT  3.150 1.020 3.270 1.375 ;
        RECT  2.900 1.145 3.150 1.375 ;
        RECT  2.780 1.020 2.900 1.375 ;
        RECT  0.310 1.145 2.780 1.375 ;
        RECT  0.230 0.980 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.070 0.355 3.115 0.485 ;
        RECT  2.970 0.710 3.115 0.800 ;
        RECT  2.990 0.185 3.070 0.485 ;
        RECT  3.865 0.370 3.885 1.055 ;
        RECT  3.815 0.260 3.865 1.055 ;
        RECT  3.790 0.260 3.815 0.440 ;
        RECT  3.795 0.735 3.815 1.055 ;
        RECT  3.575 0.370 3.790 0.440 ;
        RECT  3.715 0.515 3.745 0.650 ;
        RECT  3.645 0.515 3.715 0.950 ;
        RECT  1.950 0.880 3.645 0.950 ;
        RECT  3.505 0.370 3.575 0.640 ;
        RECT  3.485 0.520 3.505 0.640 ;
        RECT  2.625 0.740 2.730 0.810 ;
        RECT  2.625 0.195 2.710 0.265 ;
        RECT  2.555 0.195 2.625 0.810 ;
        RECT  2.100 0.205 2.555 0.275 ;
        RECT  2.300 0.730 2.370 0.810 ;
        RECT  2.300 0.345 2.325 0.465 ;
        RECT  2.230 0.345 2.300 0.810 ;
        RECT  2.180 0.500 2.230 0.640 ;
        RECT  2.100 0.710 2.160 0.810 ;
        RECT  2.030 0.205 2.100 0.810 ;
        RECT  1.870 0.195 1.950 0.950 ;
        RECT  1.690 0.195 1.770 1.065 ;
        RECT  0.670 0.995 1.690 1.065 ;
        RECT  1.225 0.855 1.610 0.925 ;
        RECT  1.365 0.715 1.450 0.785 ;
        RECT  1.365 0.185 1.420 0.285 ;
        RECT  1.305 0.185 1.365 0.785 ;
        RECT  1.295 0.205 1.305 0.785 ;
        RECT  0.820 0.205 1.295 0.275 ;
        RECT  1.150 0.745 1.225 0.925 ;
        RECT  1.020 0.350 1.070 0.450 ;
        RECT  1.020 0.775 1.070 0.855 ;
        RECT  0.950 0.350 1.020 0.855 ;
        RECT  0.900 0.520 0.950 0.640 ;
        RECT  0.820 0.755 0.870 0.875 ;
        RECT  0.750 0.205 0.820 0.875 ;
        RECT  0.590 0.230 0.670 1.065 ;
        RECT  0.410 0.230 0.490 0.415 ;
        RECT  0.410 0.840 0.490 1.025 ;
        RECT  0.125 0.345 0.410 0.415 ;
        RECT  0.125 0.840 0.410 0.910 ;
        RECT  0.055 0.195 0.125 1.070 ;
    END
END MUX3ND4BWP

MACRO MUX4D0BWP
    CLASS CORE ;
    FOREIGN MUX4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.195 3.325 0.960 ;
        RECT  3.235 0.195 3.255 0.335 ;
        RECT  3.240 0.840 3.255 0.960 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0306 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.355 3.045 0.655 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.615 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.770 0.495 0.875 0.650 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.905 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.410 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.115 3.360 0.115 ;
        RECT  3.040 -0.115 3.140 0.275 ;
        RECT  1.290 -0.115 3.040 0.115 ;
        RECT  1.200 -0.115 1.290 0.260 ;
        RECT  0.990 -0.115 1.200 0.115 ;
        RECT  0.920 -0.115 0.990 0.235 ;
        RECT  0.140 -0.115 0.920 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 3.360 1.375 ;
        RECT  1.200 1.050 1.320 1.375 ;
        RECT  0.960 1.145 1.200 1.375 ;
        RECT  0.840 1.050 0.960 1.375 ;
        RECT  0.130 1.145 0.840 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.170 0.605 3.185 0.785 ;
        RECT  3.115 0.605 3.170 1.050 ;
        RECT  3.100 0.725 3.115 1.050 ;
        RECT  2.570 0.980 3.100 1.050 ;
        RECT  2.900 0.195 2.970 0.275 ;
        RECT  2.900 0.820 2.970 0.900 ;
        RECT  2.830 0.195 2.900 0.900 ;
        RECT  2.780 0.590 2.830 0.710 ;
        RECT  2.710 0.350 2.760 0.470 ;
        RECT  2.710 0.790 2.730 0.910 ;
        RECT  2.640 0.200 2.710 0.910 ;
        RECT  1.765 0.200 2.640 0.270 ;
        RECT  2.480 0.350 2.570 1.050 ;
        RECT  2.340 0.350 2.410 1.055 ;
        RECT  2.290 0.350 2.340 0.420 ;
        RECT  1.470 0.985 2.340 1.055 ;
        RECT  1.960 0.845 2.010 0.915 ;
        RECT  1.960 0.345 1.990 0.445 ;
        RECT  1.890 0.345 1.960 0.915 ;
        RECT  1.765 0.835 1.810 0.915 ;
        RECT  1.695 0.200 1.765 0.915 ;
        RECT  1.690 0.370 1.695 0.915 ;
        RECT  1.660 0.370 1.690 0.470 ;
        RECT  1.430 0.205 1.625 0.275 ;
        RECT  1.500 0.370 1.570 0.835 ;
        RECT  1.445 0.755 1.500 0.835 ;
        RECT  1.400 0.910 1.470 1.055 ;
        RECT  1.360 0.205 1.430 0.400 ;
        RECT  0.500 0.910 1.400 0.980 ;
        RECT  1.085 0.330 1.360 0.400 ;
        RECT  1.015 0.330 1.085 0.830 ;
        RECT  0.840 0.330 1.015 0.400 ;
        RECT  0.770 0.200 0.840 0.400 ;
        RECT  0.510 0.200 0.770 0.270 ;
        RECT  0.690 0.740 0.740 0.810 ;
        RECT  0.620 0.355 0.690 0.810 ;
        RECT  0.400 0.345 0.500 0.980 ;
        RECT  0.260 0.205 0.330 0.990 ;
        RECT  0.210 0.205 0.260 0.285 ;
        RECT  0.210 0.910 0.260 0.990 ;
    END
END MUX4D0BWP

MACRO MUX4D1BWP
    CLASS CORE ;
    FOREIGN MUX4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.195 3.325 1.070 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.520 2.250 0.640 ;
        RECT  2.135 0.355 2.205 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.770 0.495 0.875 0.650 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.485 2.065 0.775 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0178 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.430 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 -0.115 3.360 0.115 ;
        RECT  3.050 -0.115 3.130 0.290 ;
        RECT  1.290 -0.115 3.050 0.115 ;
        RECT  1.200 -0.115 1.290 0.260 ;
        RECT  1.010 -0.115 1.200 0.115 ;
        RECT  0.940 -0.115 1.010 0.235 ;
        RECT  0.140 -0.115 0.940 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.145 3.360 1.375 ;
        RECT  3.050 0.890 3.130 1.375 ;
        RECT  1.320 1.145 3.050 1.375 ;
        RECT  1.200 1.040 1.320 1.375 ;
        RECT  0.940 1.145 1.200 1.375 ;
        RECT  0.820 1.040 0.940 1.375 ;
        RECT  0.140 1.145 0.820 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.090 0.370 3.160 0.810 ;
        RECT  2.910 0.370 3.090 0.440 ;
        RECT  2.950 0.740 3.090 0.810 ;
        RECT  2.760 0.540 3.020 0.660 ;
        RECT  2.870 0.740 2.950 1.065 ;
        RECT  2.840 0.195 2.910 0.440 ;
        RECT  1.765 0.195 2.840 0.265 ;
        RECT  2.690 0.345 2.760 1.065 ;
        RECT  2.570 0.350 2.610 0.915 ;
        RECT  2.540 0.350 2.570 1.065 ;
        RECT  2.470 0.350 2.540 0.420 ;
        RECT  2.490 0.755 2.540 1.065 ;
        RECT  1.470 0.995 2.490 1.065 ;
        RECT  2.390 0.555 2.470 0.675 ;
        RECT  2.320 0.350 2.390 0.915 ;
        RECT  1.915 0.335 2.010 0.405 ;
        RECT  1.915 0.855 2.000 0.925 ;
        RECT  1.845 0.335 1.915 0.925 ;
        RECT  1.695 0.195 1.765 0.925 ;
        RECT  1.430 0.200 1.620 0.280 ;
        RECT  1.500 0.365 1.570 0.830 ;
        RECT  1.445 0.755 1.500 0.830 ;
        RECT  1.400 0.900 1.470 1.065 ;
        RECT  1.360 0.200 1.430 0.400 ;
        RECT  0.485 0.900 1.400 0.970 ;
        RECT  1.085 0.330 1.360 0.400 ;
        RECT  1.015 0.330 1.085 0.820 ;
        RECT  0.860 0.330 1.015 0.400 ;
        RECT  0.790 0.205 0.860 0.400 ;
        RECT  0.530 0.205 0.790 0.275 ;
        RECT  0.630 0.355 0.700 0.830 ;
        RECT  0.485 0.380 0.550 0.460 ;
        RECT  0.415 0.380 0.485 1.060 ;
        RECT  0.305 0.215 0.330 0.880 ;
        RECT  0.260 0.215 0.305 1.060 ;
        RECT  0.210 0.215 0.260 0.295 ;
        RECT  0.235 0.800 0.260 1.060 ;
    END
END MUX4D1BWP

MACRO MUX4D2BWP
    CLASS CORE ;
    FOREIGN MUX4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.355 4.585 0.905 ;
        RECT  4.515 0.185 4.530 1.055 ;
        RECT  4.460 0.185 4.515 0.455 ;
        RECT  4.450 0.795 4.515 1.055 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.520 3.490 0.640 ;
        RECT  3.455 0.355 3.465 0.640 ;
        RECT  3.385 0.355 3.455 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 0.995 2.480 1.075 ;
        RECT  1.230 0.995 2.340 1.065 ;
        RECT  1.110 0.995 1.230 1.075 ;
        RECT  1.010 0.995 1.110 1.065 ;
        RECT  0.940 0.845 1.010 1.065 ;
        RECT  0.630 0.845 0.940 0.915 ;
        RECT  0.560 0.840 0.630 0.915 ;
        RECT  0.320 0.840 0.560 0.910 ;
        RECT  0.250 0.740 0.320 0.910 ;
        RECT  0.240 0.485 0.250 0.910 ;
        RECT  0.175 0.485 0.240 0.810 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.215 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.205 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.790 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.300 ;
        RECT  0.000 -0.115 4.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.960 4.710 1.375 ;
        RECT  4.350 1.145 4.630 1.375 ;
        RECT  4.270 0.740 4.350 1.375 ;
        RECT  0.000 1.145 4.270 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.380 0.530 4.430 0.630 ;
        RECT  4.300 0.195 4.380 0.630 ;
        RECT  3.980 0.195 4.300 0.265 ;
        RECT  4.090 0.345 4.170 1.055 ;
        RECT  2.630 0.985 4.090 1.055 ;
        RECT  3.910 0.195 3.980 0.900 ;
        RECT  3.760 0.195 3.830 0.900 ;
        RECT  2.680 0.195 3.760 0.265 ;
        RECT  3.720 0.740 3.760 0.900 ;
        RECT  3.650 0.520 3.680 0.640 ;
        RECT  3.580 0.335 3.650 0.860 ;
        RECT  3.540 0.335 3.580 0.455 ;
        RECT  3.540 0.720 3.580 0.860 ;
        RECT  2.850 0.335 3.270 0.415 ;
        RECT  2.850 0.845 3.270 0.915 ;
        RECT  2.770 0.335 2.850 0.915 ;
        RECT  2.610 0.195 2.680 0.785 ;
        RECT  2.560 0.855 2.630 1.055 ;
        RECT  2.540 0.715 2.610 0.785 ;
        RECT  1.150 0.855 2.560 0.925 ;
        RECT  2.420 0.185 2.540 0.280 ;
        RECT  2.430 0.350 2.510 0.430 ;
        RECT  2.360 0.350 2.430 0.780 ;
        RECT  1.700 0.210 2.420 0.280 ;
        RECT  1.990 0.350 2.360 0.420 ;
        RECT  1.930 0.710 2.360 0.780 ;
        RECT  1.320 0.350 1.770 0.420 ;
        RECT  1.320 0.710 1.710 0.780 ;
        RECT  1.630 0.195 1.700 0.280 ;
        RECT  1.310 0.195 1.630 0.265 ;
        RECT  1.250 0.350 1.320 0.780 ;
        RECT  1.190 0.185 1.310 0.265 ;
        RECT  1.220 0.680 1.250 0.780 ;
        RECT  0.125 0.195 1.190 0.265 ;
        RECT  1.150 0.335 1.160 0.620 ;
        RECT  1.080 0.335 1.150 0.925 ;
        RECT  1.020 0.335 1.080 0.405 ;
        RECT  0.960 0.685 1.080 0.775 ;
        RECT  0.890 0.335 0.910 0.495 ;
        RECT  0.820 0.335 0.890 0.775 ;
        RECT  0.490 0.995 0.870 1.065 ;
        RECT  0.430 0.335 0.820 0.415 ;
        RECT  0.770 0.700 0.820 0.775 ;
        RECT  0.400 0.700 0.770 0.770 ;
        RECT  0.420 0.980 0.490 1.065 ;
        RECT  0.125 0.980 0.420 1.050 ;
        RECT  0.105 0.195 0.125 0.380 ;
        RECT  0.105 0.890 0.125 1.050 ;
        RECT  0.035 0.195 0.105 1.050 ;
    END
END MUX4D2BWP

MACRO MUX4D4BWP
    CLASS CORE ;
    FOREIGN MUX4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.865 0.185 4.955 0.465 ;
        RECT  4.865 0.775 4.955 1.055 ;
        RECT  4.795 0.345 4.865 0.465 ;
        RECT  4.795 0.775 4.865 0.905 ;
        RECT  4.595 0.345 4.795 0.905 ;
        RECT  4.585 0.185 4.595 1.055 ;
        RECT  4.515 0.185 4.585 0.465 ;
        RECT  4.515 0.775 4.585 1.055 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.495 3.570 0.640 ;
        RECT  3.395 0.495 3.465 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0434 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.420 0.995 2.560 1.075 ;
        RECT  1.270 0.995 2.420 1.065 ;
        RECT  1.150 0.995 1.270 1.075 ;
        RECT  1.050 0.995 1.150 1.065 ;
        RECT  0.980 0.845 1.050 1.065 ;
        RECT  0.320 0.845 0.980 0.915 ;
        RECT  0.250 0.740 0.320 0.915 ;
        RECT  0.240 0.485 0.250 0.915 ;
        RECT  0.175 0.485 0.240 0.810 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.325 0.625 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.205 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.675 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.790 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.485 ;
        RECT  4.775 -0.115 5.050 0.115 ;
        RECT  4.685 -0.115 4.775 0.265 ;
        RECT  0.000 -0.115 4.685 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.145 5.180 1.375 ;
        RECT  5.050 0.665 5.130 1.375 ;
        RECT  4.770 1.145 5.050 1.375 ;
        RECT  4.690 0.985 4.770 1.375 ;
        RECT  4.410 1.145 4.690 1.375 ;
        RECT  4.330 0.755 4.410 1.375 ;
        RECT  3.500 1.145 4.330 1.375 ;
        RECT  3.380 1.030 3.500 1.375 ;
        RECT  3.140 1.145 3.380 1.375 ;
        RECT  3.000 1.025 3.140 1.375 ;
        RECT  0.000 1.145 3.000 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.185 4.955 0.465 ;
        RECT  4.865 0.775 4.955 1.055 ;
        RECT  4.425 0.545 4.505 0.620 ;
        RECT  4.355 0.195 4.425 0.620 ;
        RECT  4.040 0.195 4.355 0.265 ;
        RECT  4.150 0.345 4.230 1.055 ;
        RECT  3.685 0.985 4.150 1.055 ;
        RECT  3.960 0.195 4.040 0.885 ;
        RECT  3.820 0.195 3.890 0.870 ;
        RECT  2.760 0.195 3.820 0.265 ;
        RECT  3.780 0.710 3.820 0.870 ;
        RECT  3.710 0.510 3.750 0.630 ;
        RECT  3.640 0.345 3.710 0.815 ;
        RECT  3.615 0.885 3.685 1.055 ;
        RECT  3.580 0.345 3.640 0.415 ;
        RECT  3.565 0.730 3.640 0.815 ;
        RECT  2.710 0.885 3.615 0.955 ;
        RECT  2.940 0.335 3.360 0.415 ;
        RECT  2.940 0.725 3.325 0.815 ;
        RECT  2.840 0.335 2.940 0.815 ;
        RECT  2.680 0.195 2.760 0.785 ;
        RECT  2.640 0.855 2.710 0.955 ;
        RECT  2.620 0.715 2.680 0.785 ;
        RECT  1.190 0.855 2.640 0.925 ;
        RECT  2.450 0.185 2.590 0.280 ;
        RECT  2.510 0.350 2.570 0.430 ;
        RECT  2.440 0.350 2.510 0.780 ;
        RECT  1.740 0.210 2.450 0.280 ;
        RECT  2.030 0.350 2.440 0.420 ;
        RECT  2.010 0.700 2.440 0.780 ;
        RECT  1.360 0.350 1.810 0.420 ;
        RECT  1.360 0.700 1.750 0.780 ;
        RECT  1.670 0.195 1.740 0.280 ;
        RECT  1.350 0.195 1.670 0.265 ;
        RECT  1.290 0.350 1.360 0.780 ;
        RECT  1.230 0.185 1.350 0.265 ;
        RECT  1.260 0.680 1.290 0.780 ;
        RECT  0.125 0.195 1.230 0.265 ;
        RECT  1.120 0.335 1.190 0.925 ;
        RECT  1.000 0.335 1.120 0.425 ;
        RECT  1.000 0.685 1.120 0.775 ;
        RECT  0.830 0.335 0.930 0.775 ;
        RECT  0.125 0.995 0.910 1.065 ;
        RECT  0.105 0.890 0.125 1.065 ;
        RECT  0.035 0.195 0.105 1.065 ;
        RECT  0.430 0.335 0.830 0.415 ;
        RECT  0.440 0.700 0.830 0.775 ;
        RECT  0.105 0.195 0.125 0.380 ;
    END
END MUX4D4BWP

MACRO MUX4ND0BWP
    CLASS CORE ;
    FOREIGN MUX4ND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1076 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.420 2.905 0.800 ;
        RECT  2.835 0.420 2.840 0.925 ;
        RECT  2.830 0.420 2.835 0.500 ;
        RECT  2.760 0.730 2.835 0.925 ;
        RECT  2.760 0.195 2.830 0.500 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0348 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.495 2.290 0.640 ;
        RECT  2.135 0.355 2.205 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.770 0.495 0.875 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.980 0.495 2.065 0.765 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.395 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 -0.115 3.080 0.115 ;
        RECT  1.200 -0.115 1.290 0.260 ;
        RECT  0.990 -0.115 1.200 0.115 ;
        RECT  0.920 -0.115 0.990 0.250 ;
        RECT  0.125 -0.115 0.920 0.115 ;
        RECT  0.055 -0.115 0.125 0.280 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 3.080 1.375 ;
        RECT  1.200 1.050 1.320 1.375 ;
        RECT  0.960 1.145 1.200 1.375 ;
        RECT  0.840 1.050 0.960 1.375 ;
        RECT  0.130 1.145 0.840 1.375 ;
        RECT  0.050 0.990 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.975 0.215 3.045 1.065 ;
        RECT  2.940 0.215 2.975 0.315 ;
        RECT  2.940 0.865 2.975 1.065 ;
        RECT  1.470 0.995 2.940 1.065 ;
        RECT  2.600 0.205 2.670 0.925 ;
        RECT  2.540 0.205 2.600 0.435 ;
        RECT  2.510 0.855 2.600 0.925 ;
        RECT  1.770 0.205 2.540 0.275 ;
        RECT  2.430 0.520 2.530 0.640 ;
        RECT  2.360 0.350 2.430 0.860 ;
        RECT  1.910 0.345 2.030 0.415 ;
        RECT  1.910 0.845 2.030 0.915 ;
        RECT  1.840 0.345 1.910 0.915 ;
        RECT  1.700 0.205 1.770 0.915 ;
        RECT  1.650 0.375 1.700 0.445 ;
        RECT  1.430 0.205 1.620 0.275 ;
        RECT  1.500 0.370 1.570 0.810 ;
        RECT  1.435 0.740 1.500 0.810 ;
        RECT  1.400 0.910 1.470 1.065 ;
        RECT  1.360 0.205 1.430 0.400 ;
        RECT  0.460 0.910 1.400 0.980 ;
        RECT  1.085 0.330 1.360 0.400 ;
        RECT  1.015 0.330 1.085 0.830 ;
        RECT  0.840 0.330 1.015 0.400 ;
        RECT  0.770 0.215 0.840 0.400 ;
        RECT  0.510 0.215 0.770 0.285 ;
        RECT  0.700 0.755 0.760 0.830 ;
        RECT  0.620 0.370 0.700 0.830 ;
        RECT  0.460 0.375 0.540 0.460 ;
        RECT  0.390 0.375 0.460 0.980 ;
        RECT  0.230 0.185 0.310 0.425 ;
        RECT  0.230 0.845 0.310 1.040 ;
        RECT  0.105 0.355 0.230 0.425 ;
        RECT  0.105 0.845 0.230 0.915 ;
        RECT  0.035 0.355 0.105 0.915 ;
    END
END MUX4ND0BWP

MACRO MUX4ND1BWP
    CLASS CORE ;
    FOREIGN MUX4ND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.195 3.745 1.045 ;
        RECT  3.660 0.195 3.675 0.475 ;
        RECT  3.650 0.725 3.675 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.625 0.770 ;
        RECT  2.530 0.495 2.555 0.640 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.770 0.495 0.875 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.065 0.630 ;
        RECT  1.970 0.510 1.995 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0178 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.430 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.180 -0.115 3.780 0.115 ;
        RECT  2.060 -0.115 2.180 0.275 ;
        RECT  1.270 -0.115 2.060 0.115 ;
        RECT  1.200 -0.115 1.270 0.260 ;
        RECT  1.010 -0.115 1.200 0.115 ;
        RECT  0.940 -0.115 1.010 0.235 ;
        RECT  0.140 -0.115 0.940 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 3.780 1.375 ;
        RECT  1.200 1.050 1.320 1.375 ;
        RECT  0.940 1.145 1.200 1.375 ;
        RECT  0.820 1.040 0.940 1.375 ;
        RECT  0.140 1.145 0.820 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.590 0.520 3.605 0.640 ;
        RECT  3.515 0.195 3.590 0.640 ;
        RECT  3.490 0.710 3.560 1.065 ;
        RECT  3.150 0.195 3.515 0.265 ;
        RECT  3.435 0.710 3.490 0.780 ;
        RECT  1.470 0.995 3.490 1.065 ;
        RECT  3.360 0.500 3.435 0.780 ;
        RECT  3.290 0.850 3.390 0.920 ;
        RECT  3.290 0.335 3.320 0.435 ;
        RECT  3.220 0.335 3.290 0.920 ;
        RECT  3.080 0.195 3.150 0.910 ;
        RECT  3.010 0.195 3.080 0.275 ;
        RECT  2.850 0.195 2.920 0.900 ;
        RECT  2.350 0.195 2.850 0.265 ;
        RECT  2.710 0.345 2.780 0.920 ;
        RECT  2.590 0.345 2.710 0.415 ;
        RECT  2.610 0.850 2.710 0.920 ;
        RECT  2.280 0.195 2.350 0.900 ;
        RECT  2.140 0.500 2.210 0.910 ;
        RECT  1.760 0.840 2.140 0.910 ;
        RECT  1.900 0.700 1.990 0.770 ;
        RECT  1.900 0.195 1.980 0.275 ;
        RECT  1.830 0.195 1.900 0.770 ;
        RECT  1.690 0.195 1.760 0.910 ;
        RECT  1.645 0.840 1.690 0.910 ;
        RECT  1.430 0.200 1.620 0.280 ;
        RECT  1.500 0.365 1.570 0.830 ;
        RECT  1.445 0.750 1.500 0.830 ;
        RECT  1.400 0.900 1.470 1.065 ;
        RECT  1.360 0.200 1.430 0.400 ;
        RECT  0.485 0.900 1.400 0.970 ;
        RECT  1.085 0.330 1.360 0.400 ;
        RECT  1.015 0.330 1.085 0.820 ;
        RECT  0.860 0.330 1.015 0.400 ;
        RECT  0.790 0.200 0.860 0.400 ;
        RECT  0.530 0.200 0.790 0.270 ;
        RECT  0.630 0.355 0.700 0.830 ;
        RECT  0.485 0.380 0.550 0.460 ;
        RECT  0.415 0.380 0.485 1.060 ;
        RECT  0.260 0.215 0.330 1.065 ;
        RECT  0.210 0.215 0.260 0.295 ;
        RECT  0.230 0.745 0.260 1.065 ;
    END
END MUX4ND1BWP

MACRO MUX4ND2BWP
    CLASS CORE ;
    FOREIGN MUX4ND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1152 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.355 3.885 0.905 ;
        RECT  3.795 0.355 3.815 0.470 ;
        RECT  3.795 0.785 3.815 0.905 ;
        RECT  3.725 0.190 3.795 0.470 ;
        RECT  3.725 0.785 3.795 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.625 0.770 ;
        RECT  2.530 0.495 2.555 0.640 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.770 0.495 0.875 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.065 0.630 ;
        RECT  1.970 0.510 1.995 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0178 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.430 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.990 -0.115 4.060 0.115 ;
        RECT  3.910 -0.115 3.990 0.285 ;
        RECT  2.180 -0.115 3.910 0.115 ;
        RECT  2.060 -0.115 2.180 0.275 ;
        RECT  1.270 -0.115 2.060 0.115 ;
        RECT  1.200 -0.115 1.270 0.260 ;
        RECT  1.010 -0.115 1.200 0.115 ;
        RECT  0.940 -0.115 1.010 0.235 ;
        RECT  0.140 -0.115 0.940 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.990 1.145 4.060 1.375 ;
        RECT  3.910 0.975 3.990 1.375 ;
        RECT  1.320 1.145 3.910 1.375 ;
        RECT  1.200 1.050 1.320 1.375 ;
        RECT  0.940 1.145 1.200 1.375 ;
        RECT  0.820 1.040 0.940 1.375 ;
        RECT  0.140 1.145 0.820 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.630 0.545 3.730 0.615 ;
        RECT  3.580 0.710 3.650 1.065 ;
        RECT  3.555 0.195 3.630 0.615 ;
        RECT  3.475 0.710 3.580 0.780 ;
        RECT  1.470 0.995 3.580 1.065 ;
        RECT  3.190 0.195 3.555 0.265 ;
        RECT  3.400 0.500 3.475 0.780 ;
        RECT  3.330 0.850 3.430 0.920 ;
        RECT  3.330 0.335 3.380 0.405 ;
        RECT  3.260 0.335 3.330 0.920 ;
        RECT  3.120 0.195 3.190 0.910 ;
        RECT  3.050 0.195 3.120 0.275 ;
        RECT  2.890 0.195 2.960 0.910 ;
        RECT  2.350 0.195 2.890 0.265 ;
        RECT  2.710 0.345 2.780 0.920 ;
        RECT  2.590 0.345 2.710 0.415 ;
        RECT  2.590 0.850 2.710 0.920 ;
        RECT  2.280 0.195 2.350 0.900 ;
        RECT  2.140 0.500 2.210 0.910 ;
        RECT  1.760 0.840 2.140 0.910 ;
        RECT  1.900 0.700 1.990 0.770 ;
        RECT  1.900 0.195 1.980 0.275 ;
        RECT  1.830 0.195 1.900 0.770 ;
        RECT  1.690 0.195 1.760 0.910 ;
        RECT  1.645 0.840 1.690 0.910 ;
        RECT  1.430 0.200 1.620 0.280 ;
        RECT  1.500 0.365 1.570 0.830 ;
        RECT  1.445 0.750 1.500 0.830 ;
        RECT  1.400 0.900 1.470 1.065 ;
        RECT  1.360 0.200 1.430 0.400 ;
        RECT  0.485 0.900 1.400 0.970 ;
        RECT  1.085 0.330 1.360 0.400 ;
        RECT  1.015 0.330 1.085 0.820 ;
        RECT  0.860 0.330 1.015 0.400 ;
        RECT  0.790 0.205 0.860 0.400 ;
        RECT  0.530 0.205 0.790 0.275 ;
        RECT  0.630 0.355 0.700 0.830 ;
        RECT  0.485 0.380 0.550 0.460 ;
        RECT  0.415 0.380 0.485 1.060 ;
        RECT  0.305 0.215 0.330 0.815 ;
        RECT  0.260 0.215 0.305 1.065 ;
        RECT  0.210 0.215 0.260 0.295 ;
        RECT  0.235 0.745 0.260 1.065 ;
    END
END MUX4ND2BWP

MACRO MUX4ND4BWP
    CLASS CORE ;
    FOREIGN MUX4ND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.575 0.185 5.645 0.485 ;
        RECT  5.575 0.775 5.645 1.055 ;
        RECT  5.495 0.355 5.575 0.485 ;
        RECT  5.495 0.775 5.575 0.905 ;
        RECT  5.285 0.355 5.495 0.905 ;
        RECT  5.215 0.185 5.285 0.465 ;
        RECT  5.215 0.775 5.285 1.055 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.545 3.920 0.615 ;
        RECT  3.675 0.495 3.745 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.0440 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 0.995 2.480 1.075 ;
        RECT  1.230 0.995 2.340 1.065 ;
        RECT  1.110 0.995 1.230 1.075 ;
        RECT  1.010 0.995 1.110 1.065 ;
        RECT  0.940 0.845 1.010 1.065 ;
        RECT  0.320 0.845 0.940 0.915 ;
        RECT  0.250 0.740 0.320 0.915 ;
        RECT  0.240 0.485 0.250 0.915 ;
        RECT  0.175 0.485 0.240 0.810 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.110 0.495 3.210 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.205 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.790 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 -0.115 5.880 0.115 ;
        RECT  5.750 -0.115 5.830 0.485 ;
        RECT  5.480 -0.115 5.750 0.115 ;
        RECT  5.380 -0.115 5.480 0.275 ;
        RECT  0.000 -0.115 5.380 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.145 5.880 1.375 ;
        RECT  5.750 0.665 5.830 1.375 ;
        RECT  5.480 1.145 5.750 1.375 ;
        RECT  5.380 0.985 5.480 1.375 ;
        RECT  5.120 1.145 5.380 1.375 ;
        RECT  5.020 0.870 5.120 1.375 ;
        RECT  0.000 1.145 5.020 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.575 0.185 5.645 0.485 ;
        RECT  5.575 0.775 5.645 1.055 ;
        RECT  5.565 0.355 5.575 0.485 ;
        RECT  5.565 0.775 5.575 0.905 ;
        RECT  5.120 0.545 5.200 0.615 ;
        RECT  5.050 0.210 5.120 0.615 ;
        RECT  4.380 0.210 5.050 0.280 ;
        RECT  4.930 0.360 4.970 0.805 ;
        RECT  4.900 0.360 4.930 1.055 ;
        RECT  4.520 0.360 4.900 0.430 ;
        RECT  4.850 0.735 4.900 1.055 ;
        RECT  4.740 0.545 4.830 0.615 ;
        RECT  4.670 0.545 4.740 1.065 ;
        RECT  4.045 0.995 4.670 1.065 ;
        RECT  4.520 0.855 4.590 0.925 ;
        RECT  4.450 0.360 4.520 0.925 ;
        RECT  4.280 0.210 4.380 0.925 ;
        RECT  4.140 0.210 4.210 0.910 ;
        RECT  3.625 0.210 4.140 0.280 ;
        RECT  3.500 0.840 4.140 0.910 ;
        RECT  4.000 0.375 4.070 0.770 ;
        RECT  3.975 0.980 4.045 1.065 ;
        RECT  3.900 0.375 4.000 0.445 ;
        RECT  3.870 0.700 4.000 0.770 ;
        RECT  2.630 0.980 3.975 1.050 ;
        RECT  3.550 0.210 3.625 0.395 ;
        RECT  3.460 0.545 3.595 0.615 ;
        RECT  3.390 0.195 3.460 0.615 ;
        RECT  2.680 0.195 3.390 0.265 ;
        RECT  2.850 0.335 3.290 0.405 ;
        RECT  2.850 0.840 3.260 0.910 ;
        RECT  2.770 0.335 2.850 0.910 ;
        RECT  2.610 0.195 2.680 0.785 ;
        RECT  2.560 0.855 2.630 1.050 ;
        RECT  2.540 0.715 2.610 0.785 ;
        RECT  1.150 0.855 2.560 0.925 ;
        RECT  2.420 0.185 2.540 0.280 ;
        RECT  2.430 0.350 2.510 0.430 ;
        RECT  2.360 0.350 2.430 0.780 ;
        RECT  1.700 0.210 2.420 0.280 ;
        RECT  2.000 0.350 2.360 0.420 ;
        RECT  1.940 0.710 2.360 0.780 ;
        RECT  1.320 0.350 1.760 0.420 ;
        RECT  1.630 0.195 1.700 0.280 ;
        RECT  1.320 0.710 1.700 0.780 ;
        RECT  1.310 0.195 1.630 0.265 ;
        RECT  1.250 0.350 1.320 0.780 ;
        RECT  1.190 0.185 1.310 0.265 ;
        RECT  1.220 0.680 1.250 0.780 ;
        RECT  0.125 0.195 1.190 0.265 ;
        RECT  1.150 0.335 1.160 0.620 ;
        RECT  1.080 0.335 1.150 0.925 ;
        RECT  1.020 0.335 1.080 0.405 ;
        RECT  0.960 0.685 1.080 0.775 ;
        RECT  0.890 0.335 0.910 0.495 ;
        RECT  0.820 0.335 0.890 0.775 ;
        RECT  0.125 0.995 0.870 1.065 ;
        RECT  0.430 0.335 0.820 0.415 ;
        RECT  0.770 0.700 0.820 0.775 ;
        RECT  0.400 0.700 0.770 0.770 ;
        RECT  0.105 0.195 0.125 0.380 ;
        RECT  0.105 0.890 0.125 1.065 ;
        RECT  0.035 0.195 0.105 1.065 ;
    END
END MUX4ND4BWP

MACRO ND2D0BWP
    CLASS CORE ;
    FOREIGN ND2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0498 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 0.915 ;
        RECT  0.435 0.185 0.455 0.305 ;
        RECT  0.315 0.845 0.455 0.915 ;
        RECT  0.245 0.845 0.315 1.060 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.450 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.560 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.145 0.560 1.375 ;
        RECT  0.420 0.985 0.520 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END ND2D0BWP

MACRO ND2D1BWP
    CLASS CORE ;
    FOREIGN ND2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0997 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.215 0.525 0.905 ;
        RECT  0.435 0.215 0.455 0.345 ;
        RECT  0.315 0.835 0.455 0.905 ;
        RECT  0.245 0.835 0.315 1.050 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.560 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 0.560 1.375 ;
        RECT  0.430 0.980 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.770 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END ND2D1BWP

MACRO ND2D2BWP
    CLASS CORE ;
    FOREIGN ND2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1582 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.835 0.730 1.035 ;
        RECT  0.390 0.835 0.650 0.915 ;
        RECT  0.385 0.345 0.390 0.915 ;
        RECT  0.315 0.345 0.385 1.045 ;
        RECT  0.270 0.345 0.315 0.415 ;
        RECT  0.290 0.705 0.315 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.495 0.805 0.765 ;
        RECT  0.630 0.495 0.730 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.740 0.275 ;
        RECT  0.000 -0.115 0.640 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.835 0.910 1.375 ;
        RECT  0.560 1.145 0.830 1.375 ;
        RECT  0.460 0.990 0.560 1.375 ;
        RECT  0.185 1.145 0.460 1.375 ;
        RECT  0.115 0.705 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 0.255 0.910 0.415 ;
        RECT  0.560 0.345 0.830 0.415 ;
        RECT  0.490 0.205 0.560 0.415 ;
        RECT  0.070 0.205 0.490 0.275 ;
    END
END ND2D2BWP

MACRO ND2D3BWP
    CLASS CORE ;
    FOREIGN ND2D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2497 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.835 1.030 0.950 ;
        RECT  0.525 0.835 0.950 0.905 ;
        RECT  0.455 0.350 0.525 0.905 ;
        RECT  0.130 0.350 0.455 0.420 ;
        RECT  0.310 0.835 0.455 0.905 ;
        RECT  0.230 0.835 0.310 0.950 ;
        RECT  0.050 0.215 0.130 0.420 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.495 1.020 0.625 ;
        RECT  0.730 0.495 0.810 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.625 ;
        RECT  0.145 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.260 0.115 ;
        RECT  1.120 -0.115 1.220 0.430 ;
        RECT  0.860 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.860 0.275 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.260 1.375 ;
        RECT  1.120 0.685 1.220 1.375 ;
        RECT  0.860 1.145 1.120 1.375 ;
        RECT  0.760 0.990 0.860 1.375 ;
        RECT  0.500 1.145 0.760 1.375 ;
        RECT  0.400 0.990 0.500 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.840 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.665 0.355 0.940 0.425 ;
        RECT  0.595 0.210 0.665 0.425 ;
        RECT  0.210 0.210 0.595 0.280 ;
    END
END ND2D3BWP

MACRO ND2D4BWP
    CLASS CORE ;
    FOREIGN ND2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3164 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.775 1.445 1.075 ;
        RECT  1.085 0.775 1.375 0.935 ;
        RECT  1.015 0.775 1.085 1.075 ;
        RECT  0.665 0.775 1.015 0.935 ;
        RECT  0.595 0.335 0.690 0.415 ;
        RECT  0.595 0.775 0.665 1.075 ;
        RECT  0.385 0.335 0.595 0.935 ;
        RECT  0.210 0.335 0.385 0.415 ;
        RECT  0.305 0.775 0.385 0.935 ;
        RECT  0.235 0.775 0.305 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.505 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.250 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 1.680 0.115 ;
        RECT  1.360 -0.115 1.460 0.270 ;
        RECT  1.100 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.100 0.270 ;
        RECT  0.000 -0.115 1.000 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.790 1.630 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 1.005 1.290 1.375 ;
        RECT  0.900 1.145 1.170 1.375 ;
        RECT  0.780 1.025 0.900 1.375 ;
        RECT  0.510 1.145 0.780 1.375 ;
        RECT  0.390 1.005 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.375 0.775 1.445 1.075 ;
        RECT  1.085 0.775 1.375 0.935 ;
        RECT  1.015 0.775 1.085 1.075 ;
        RECT  0.665 0.775 1.015 0.935 ;
        RECT  0.665 0.335 0.690 0.415 ;
        RECT  0.210 0.335 0.315 0.415 ;
        RECT  0.305 0.775 0.315 0.935 ;
        RECT  0.235 0.775 0.305 1.075 ;
        RECT  1.555 0.230 1.625 0.415 ;
        RECT  0.880 0.345 1.555 0.415 ;
        RECT  0.800 0.195 0.880 0.415 ;
        RECT  0.125 0.195 0.800 0.265 ;
        RECT  0.055 0.195 0.125 0.375 ;
    END
END ND2D4BWP

MACRO ND2D8BWP
    CLASS CORE ;
    FOREIGN ND2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6328 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.780 2.845 1.075 ;
        RECT  2.485 0.780 2.775 0.935 ;
        RECT  2.415 0.780 2.485 1.075 ;
        RECT  2.125 0.780 2.415 0.935 ;
        RECT  2.055 0.780 2.125 1.075 ;
        RECT  1.765 0.780 2.055 0.935 ;
        RECT  1.695 0.780 1.765 1.075 ;
        RECT  1.385 0.780 1.695 0.935 ;
        RECT  1.295 0.335 1.410 0.425 ;
        RECT  1.315 0.780 1.385 1.075 ;
        RECT  1.295 0.780 1.315 0.935 ;
        RECT  1.085 0.335 1.295 0.935 ;
        RECT  0.210 0.335 1.085 0.425 ;
        RECT  1.025 0.780 1.085 0.935 ;
        RECT  0.955 0.780 1.025 1.075 ;
        RECT  0.665 0.780 0.955 0.935 ;
        RECT  0.595 0.780 0.665 1.075 ;
        RECT  0.305 0.780 0.595 0.935 ;
        RECT  0.235 0.780 0.305 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.635 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.955 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 -0.115 3.080 0.115 ;
        RECT  2.760 -0.115 2.860 0.270 ;
        RECT  2.500 -0.115 2.760 0.115 ;
        RECT  2.400 -0.115 2.500 0.270 ;
        RECT  2.140 -0.115 2.400 0.115 ;
        RECT  2.040 -0.115 2.140 0.270 ;
        RECT  1.780 -0.115 2.040 0.115 ;
        RECT  1.680 -0.115 1.780 0.270 ;
        RECT  0.000 -0.115 1.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.780 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 1.005 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 1.005 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.005 1.970 1.375 ;
        RECT  1.600 1.145 1.850 1.375 ;
        RECT  1.480 1.025 1.600 1.375 ;
        RECT  1.230 1.145 1.480 1.375 ;
        RECT  1.110 1.005 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 1.005 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 1.005 0.510 1.375 ;
        RECT  0.125 1.145 0.390 1.375 ;
        RECT  0.055 0.780 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.775 0.780 2.845 1.075 ;
        RECT  2.485 0.780 2.775 0.935 ;
        RECT  2.415 0.780 2.485 1.075 ;
        RECT  2.125 0.780 2.415 0.935 ;
        RECT  2.055 0.780 2.125 1.075 ;
        RECT  1.765 0.780 2.055 0.935 ;
        RECT  1.695 0.780 1.765 1.075 ;
        RECT  1.385 0.780 1.695 0.935 ;
        RECT  1.365 0.335 1.410 0.425 ;
        RECT  1.365 0.780 1.385 1.075 ;
        RECT  0.210 0.335 1.015 0.425 ;
        RECT  0.955 0.780 1.015 1.075 ;
        RECT  0.665 0.780 0.955 0.935 ;
        RECT  0.595 0.780 0.665 1.075 ;
        RECT  0.305 0.780 0.595 0.935 ;
        RECT  0.235 0.780 0.305 1.075 ;
        RECT  2.955 0.235 3.025 0.415 ;
        RECT  1.580 0.345 2.955 0.415 ;
        RECT  1.500 0.195 1.580 0.415 ;
        RECT  0.125 0.195 1.500 0.265 ;
        RECT  0.055 0.195 0.125 0.375 ;
    END
END ND2D8BWP

MACRO ND3D0BWP
    CLASS CORE ;
    FOREIGN ND3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0899 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.205 0.805 0.915 ;
        RECT  0.630 0.205 0.735 0.275 ;
        RECT  0.725 0.845 0.735 0.915 ;
        RECT  0.655 0.845 0.725 1.060 ;
        RECT  0.380 0.845 0.655 0.915 ;
        RECT  0.295 0.845 0.380 1.060 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.435 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.665 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.210 -0.115 0.840 0.115 ;
        RECT  0.090 -0.115 0.210 0.270 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.145 0.840 1.375 ;
        RECT  0.450 0.995 0.570 1.375 ;
        RECT  0.185 1.145 0.450 1.375 ;
        RECT  0.115 0.920 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
END ND3D0BWP

MACRO ND3D1BWP
    CLASS CORE ;
    FOREIGN ND3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1612 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.185 0.805 1.070 ;
        RECT  0.385 0.730 0.715 0.800 ;
        RECT  0.260 0.730 0.385 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.520 0.390 0.650 ;
        RECT  0.315 0.325 0.385 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.565 0.380 0.645 0.650 ;
        RECT  0.525 0.380 0.565 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.130 0.410 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.145 0.840 1.375 ;
        RECT  0.500 0.895 0.580 1.375 ;
        RECT  0.140 1.145 0.500 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND3D1BWP

MACRO ND3D2BWP
    CLASS CORE ;
    FOREIGN ND3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2876 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.290 1.365 1.045 ;
        RECT  1.085 0.290 1.280 0.360 ;
        RECT  0.940 0.835 1.280 0.905 ;
        RECT  1.015 0.195 1.085 0.360 ;
        RECT  0.595 0.195 1.015 0.265 ;
        RECT  0.860 0.835 0.940 1.070 ;
        RECT  0.540 0.835 0.860 0.905 ;
        RECT  0.460 0.835 0.540 1.070 ;
        RECT  0.140 0.835 0.460 0.905 ;
        RECT  0.035 0.735 0.140 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.430 1.205 0.640 ;
        RECT  0.945 0.430 1.135 0.500 ;
        RECT  0.875 0.335 0.945 0.500 ;
        RECT  0.245 0.335 0.875 0.405 ;
        RECT  0.175 0.335 0.245 0.625 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.570 1.040 0.640 ;
        RECT  0.875 0.570 0.945 0.765 ;
        RECT  0.525 0.695 0.875 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.315 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.230 -0.115 1.350 0.220 ;
        RECT  0.140 -0.115 1.230 0.115 ;
        RECT  0.070 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.145 1.400 1.375 ;
        RECT  1.060 0.975 1.140 1.375 ;
        RECT  0.740 1.145 1.060 1.375 ;
        RECT  0.660 0.975 0.740 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.260 0.975 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
END ND3D2BWP

MACRO ND3D3BWP
    CLASS CORE ;
    FOREIGN ND3D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3522 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.510 0.845 1.590 1.055 ;
        RECT  1.210 0.845 1.510 0.935 ;
        RECT  1.130 0.845 1.210 1.055 ;
        RECT  0.850 0.845 1.130 0.935 ;
        RECT  0.770 0.845 0.850 1.055 ;
        RECT  0.595 0.845 0.770 0.935 ;
        RECT  0.490 0.350 0.595 0.935 ;
        RECT  0.410 0.350 0.490 1.055 ;
        RECT  0.385 0.350 0.410 0.935 ;
        RECT  0.130 0.350 0.385 0.420 ;
        RECT  0.130 0.845 0.385 0.935 ;
        RECT  0.050 0.215 0.130 0.420 ;
        RECT  0.050 0.845 0.130 1.055 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.645 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.085 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.280 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.440 ;
        RECT  1.420 -0.115 1.690 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.000 -0.115 1.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.680 1.770 1.375 ;
        RECT  1.420 1.145 1.690 1.375 ;
        RECT  1.300 1.010 1.420 1.375 ;
        RECT  1.050 1.145 1.300 1.375 ;
        RECT  0.930 1.010 1.050 1.375 ;
        RECT  0.690 1.145 0.930 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.330 1.145 0.570 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.510 0.845 1.590 1.055 ;
        RECT  1.210 0.845 1.510 0.935 ;
        RECT  1.130 0.845 1.210 1.055 ;
        RECT  0.850 0.845 1.130 0.935 ;
        RECT  0.770 0.845 0.850 1.055 ;
        RECT  0.665 0.845 0.770 0.935 ;
        RECT  0.130 0.350 0.315 0.420 ;
        RECT  0.130 0.845 0.315 0.935 ;
        RECT  0.050 0.215 0.130 0.420 ;
        RECT  0.050 0.845 0.130 1.055 ;
        RECT  1.490 0.210 1.610 0.415 ;
        RECT  1.210 0.345 1.490 0.415 ;
        RECT  1.130 0.185 1.210 0.415 ;
        RECT  0.730 0.345 1.130 0.415 ;
        RECT  0.210 0.205 1.050 0.275 ;
    END
END ND3D3BWP

MACRO ND3D4BWP
    CLASS CORE ;
    FOREIGN ND3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4312 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.345 2.310 0.465 ;
        RECT  2.215 0.695 2.285 1.035 ;
        RECT  1.995 0.695 2.215 0.800 ;
        RECT  1.925 0.345 1.995 0.800 ;
        RECT  1.855 0.345 1.925 1.035 ;
        RECT  1.785 0.345 1.855 0.800 ;
        RECT  1.565 0.695 1.785 0.800 ;
        RECT  1.495 0.695 1.565 1.035 ;
        RECT  1.205 0.695 1.495 0.800 ;
        RECT  1.135 0.695 1.205 1.035 ;
        RECT  0.665 0.695 1.135 0.800 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.695 0.595 0.800 ;
        RECT  0.235 0.695 0.305 1.035 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.495 0.755 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 0.495 1.595 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.395 0.355 2.485 0.625 ;
        RECT  2.085 0.545 2.395 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.850 -0.115 2.520 0.115 ;
        RECT  0.770 -0.115 0.850 0.285 ;
        RECT  0.485 -0.115 0.770 0.115 ;
        RECT  0.415 -0.115 0.485 0.285 ;
        RECT  0.130 -0.115 0.415 0.115 ;
        RECT  0.050 -0.115 0.130 0.465 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.710 2.480 1.375 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.020 0.870 2.120 1.375 ;
        RECT  1.760 1.145 2.020 1.375 ;
        RECT  1.660 0.870 1.760 1.375 ;
        RECT  1.400 1.145 1.660 1.375 ;
        RECT  1.300 0.870 1.400 1.375 ;
        RECT  1.040 1.145 1.300 1.375 ;
        RECT  0.940 0.870 1.040 1.375 ;
        RECT  0.860 1.145 0.940 1.375 ;
        RECT  0.760 0.870 0.860 1.375 ;
        RECT  0.500 1.145 0.760 1.375 ;
        RECT  0.400 0.870 0.500 1.375 ;
        RECT  0.130 1.145 0.400 1.375 ;
        RECT  0.050 0.680 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.065 0.695 2.215 0.800 ;
        RECT  1.565 0.695 1.715 0.800 ;
        RECT  1.495 0.695 1.565 1.035 ;
        RECT  1.205 0.695 1.495 0.800 ;
        RECT  1.135 0.695 1.205 1.035 ;
        RECT  0.665 0.695 1.135 0.800 ;
        RECT  0.595 0.695 0.665 1.035 ;
        RECT  0.305 0.695 0.595 0.800 ;
        RECT  0.235 0.695 0.305 1.035 ;
        RECT  2.380 0.185 2.480 0.285 ;
        RECT  0.930 0.205 2.380 0.275 ;
        RECT  0.665 0.355 1.590 0.425 ;
        RECT  0.595 0.185 0.665 0.425 ;
        RECT  0.320 0.355 0.595 0.425 ;
        RECT  0.220 0.185 0.320 0.425 ;
        RECT  2.065 0.345 2.310 0.465 ;
        RECT  2.215 0.695 2.285 1.035 ;
    END
END ND3D4BWP

MACRO ND3D8BWP
    CLASS CORE ;
    FOREIGN ND3D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8624 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.355 4.490 0.425 ;
        RECT  4.380 0.705 4.480 0.970 ;
        RECT  4.110 0.705 4.380 0.815 ;
        RECT  4.095 0.705 4.110 0.990 ;
        RECT  4.030 0.355 4.095 0.990 ;
        RECT  3.885 0.355 4.030 0.815 ;
        RECT  3.290 0.355 3.885 0.425 ;
        RECT  3.750 0.705 3.885 0.815 ;
        RECT  3.670 0.705 3.750 0.990 ;
        RECT  3.390 0.705 3.670 0.815 ;
        RECT  3.310 0.705 3.390 0.990 ;
        RECT  2.850 0.705 3.310 0.815 ;
        RECT  2.770 0.705 2.850 0.990 ;
        RECT  2.490 0.705 2.770 0.815 ;
        RECT  2.410 0.705 2.490 0.990 ;
        RECT  2.130 0.705 2.410 0.815 ;
        RECT  2.050 0.705 2.130 0.990 ;
        RECT  1.770 0.705 2.050 0.815 ;
        RECT  1.690 0.705 1.770 0.990 ;
        RECT  1.410 0.705 1.690 0.815 ;
        RECT  1.330 0.705 1.410 0.990 ;
        RECT  1.050 0.705 1.330 0.815 ;
        RECT  0.970 0.705 1.050 0.990 ;
        RECT  0.690 0.705 0.970 0.815 ;
        RECT  0.610 0.705 0.690 0.990 ;
        RECT  0.340 0.705 0.610 0.815 ;
        RECT  0.240 0.705 0.340 0.970 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 1.365 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 2.905 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.495 3.745 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 -0.115 4.760 0.115 ;
        RECT  1.330 -0.115 1.410 0.285 ;
        RECT  1.050 -0.115 1.330 0.115 ;
        RECT  0.970 -0.115 1.050 0.285 ;
        RECT  0.690 -0.115 0.970 0.115 ;
        RECT  0.610 -0.115 0.690 0.285 ;
        RECT  0.330 -0.115 0.610 0.115 ;
        RECT  0.250 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 1.145 4.760 1.375 ;
        RECT  4.575 0.695 4.645 1.375 ;
        RECT  4.310 1.145 4.575 1.375 ;
        RECT  4.190 0.885 4.310 1.375 ;
        RECT  3.950 1.145 4.190 1.375 ;
        RECT  3.830 0.885 3.950 1.375 ;
        RECT  3.590 1.145 3.830 1.375 ;
        RECT  3.470 0.885 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.130 0.885 3.210 1.375 ;
        RECT  3.030 1.145 3.130 1.375 ;
        RECT  2.950 0.885 3.030 1.375 ;
        RECT  2.690 1.145 2.950 1.375 ;
        RECT  2.570 0.885 2.690 1.375 ;
        RECT  2.330 1.145 2.570 1.375 ;
        RECT  2.210 0.885 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 0.885 1.970 1.375 ;
        RECT  1.610 1.145 1.850 1.375 ;
        RECT  1.490 0.885 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 0.885 1.250 1.375 ;
        RECT  0.890 1.145 1.130 1.375 ;
        RECT  0.770 0.885 0.890 1.375 ;
        RECT  0.530 1.145 0.770 1.375 ;
        RECT  0.410 0.885 0.530 1.375 ;
        RECT  0.150 1.145 0.410 1.375 ;
        RECT  0.070 0.695 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.355 4.490 0.425 ;
        RECT  4.380 0.705 4.480 0.970 ;
        RECT  4.165 0.705 4.380 0.815 ;
        RECT  3.290 0.355 3.815 0.425 ;
        RECT  3.750 0.705 3.815 0.815 ;
        RECT  3.670 0.705 3.750 0.990 ;
        RECT  3.390 0.705 3.670 0.815 ;
        RECT  3.310 0.705 3.390 0.990 ;
        RECT  2.850 0.705 3.310 0.815 ;
        RECT  2.770 0.705 2.850 0.990 ;
        RECT  2.490 0.705 2.770 0.815 ;
        RECT  2.410 0.705 2.490 0.990 ;
        RECT  2.130 0.705 2.410 0.815 ;
        RECT  2.050 0.705 2.130 0.990 ;
        RECT  1.770 0.705 2.050 0.815 ;
        RECT  1.690 0.705 1.770 0.990 ;
        RECT  1.410 0.705 1.690 0.815 ;
        RECT  1.330 0.705 1.410 0.990 ;
        RECT  1.050 0.705 1.330 0.815 ;
        RECT  0.970 0.705 1.050 0.990 ;
        RECT  0.690 0.705 0.970 0.815 ;
        RECT  0.610 0.705 0.690 0.990 ;
        RECT  0.340 0.705 0.610 0.815 ;
        RECT  0.240 0.705 0.340 0.970 ;
        RECT  4.575 0.215 4.645 0.475 ;
        RECT  1.670 0.215 4.575 0.285 ;
        RECT  4.230 0.550 4.540 0.625 ;
        RECT  1.585 0.355 3.050 0.425 ;
        RECT  1.515 0.185 1.585 0.425 ;
        RECT  1.225 0.355 1.515 0.425 ;
        RECT  1.155 0.185 1.225 0.425 ;
        RECT  0.865 0.355 1.155 0.425 ;
        RECT  0.795 0.185 0.865 0.425 ;
        RECT  0.505 0.355 0.795 0.425 ;
        RECT  0.435 0.185 0.505 0.425 ;
        RECT  0.160 0.355 0.435 0.425 ;
        RECT  0.060 0.185 0.160 0.425 ;
    END
END ND3D8BWP

MACRO ND4D0BWP
    CLASS CORE ;
    FOREIGN ND4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0775 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.205 0.945 0.855 ;
        RECT  0.810 0.205 0.875 0.275 ;
        RECT  0.725 0.785 0.875 0.855 ;
        RECT  0.655 0.785 0.725 1.065 ;
        RECT  0.305 0.785 0.655 0.855 ;
        RECT  0.235 0.785 0.305 1.065 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.670 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.640 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.670 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.980 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.925 0.910 1.375 ;
        RECT  0.530 1.145 0.830 1.375 ;
        RECT  0.430 0.925 0.530 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.925 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END ND4D0BWP

MACRO ND4D1BWP
    CLASS CORE ;
    FOREIGN ND4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1551 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 0.810 ;
        RECT  0.810 0.195 0.875 0.265 ;
        RECT  0.730 0.740 0.875 0.810 ;
        RECT  0.650 0.740 0.730 1.035 ;
        RECT  0.310 0.740 0.650 0.810 ;
        RECT  0.235 0.740 0.310 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.640 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.980 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.810 0.880 0.930 1.375 ;
        RECT  0.535 1.145 0.810 1.375 ;
        RECT  0.415 0.880 0.535 1.375 ;
        RECT  0.140 1.145 0.415 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND4D1BWP

MACRO ND4D2BWP
    CLASS CORE ;
    FOREIGN ND4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2730 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.835 1.590 1.075 ;
        RECT  1.220 0.835 1.490 0.905 ;
        RECT  1.140 0.835 1.220 1.075 ;
        RECT  0.680 0.835 1.140 0.905 ;
        RECT  0.600 0.835 0.680 1.075 ;
        RECT  0.385 0.835 0.600 0.905 ;
        RECT  0.315 0.345 0.385 0.905 ;
        RECT  0.220 0.345 0.315 0.415 ;
        RECT  0.245 0.735 0.315 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.545 1.645 0.625 ;
        RECT  1.430 0.495 1.505 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.495 1.225 0.765 ;
        RECT  1.105 0.495 1.145 0.615 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.545 0.715 0.615 ;
        RECT  0.525 0.545 0.545 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 -0.115 1.820 0.115 ;
        RECT  1.500 -0.115 1.580 0.285 ;
        RECT  0.000 -0.115 1.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.670 0.705 1.770 1.375 ;
        RECT  1.400 1.145 1.670 1.375 ;
        RECT  1.320 0.975 1.400 1.375 ;
        RECT  1.040 1.145 1.320 1.375 ;
        RECT  0.960 0.975 1.040 1.375 ;
        RECT  0.860 1.145 0.960 1.375 ;
        RECT  0.780 0.975 0.860 1.375 ;
        RECT  0.500 1.145 0.780 1.375 ;
        RECT  0.420 0.975 0.500 1.375 ;
        RECT  0.150 1.145 0.420 1.375 ;
        RECT  0.050 0.705 0.150 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 0.185 1.770 0.430 ;
        RECT  1.400 0.355 1.670 0.425 ;
        RECT  1.320 0.205 1.400 0.425 ;
        RECT  0.940 0.205 1.320 0.275 ;
        RECT  1.040 0.355 1.240 0.425 ;
        RECT  0.970 0.355 1.040 0.445 ;
        RECT  0.690 0.375 0.970 0.445 ;
        RECT  0.770 0.195 0.870 0.295 ;
        RECT  0.040 0.195 0.770 0.265 ;
        RECT  0.590 0.345 0.690 0.445 ;
    END
END ND4D2BWP

MACRO ND4D3BWP
    CLASS CORE ;
    FOREIGN ND4D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4773 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.230 0.700 2.310 1.035 ;
        RECT  1.950 0.700 2.230 0.815 ;
        RECT  1.870 0.700 1.950 1.035 ;
        RECT  1.590 0.700 1.870 0.815 ;
        RECT  1.510 0.700 1.590 1.035 ;
        RECT  1.230 0.700 1.510 0.815 ;
        RECT  1.150 0.700 1.230 1.035 ;
        RECT  0.870 0.700 1.150 0.815 ;
        RECT  0.790 0.700 0.870 1.035 ;
        RECT  0.785 0.700 0.790 0.960 ;
        RECT  0.595 0.845 0.785 0.960 ;
        RECT  0.510 0.355 0.595 0.960 ;
        RECT  0.430 0.355 0.510 1.035 ;
        RECT  0.385 0.355 0.430 0.960 ;
        RECT  0.160 0.355 0.385 0.425 ;
        RECT  0.150 0.845 0.385 0.960 ;
        RECT  0.060 0.185 0.160 0.425 ;
        RECT  0.070 0.845 0.150 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.205 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.645 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.090 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.295 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 -0.115 2.380 0.115 ;
        RECT  2.230 -0.115 2.310 0.425 ;
        RECT  1.970 -0.115 2.230 0.115 ;
        RECT  1.850 -0.115 1.970 0.285 ;
        RECT  0.000 -0.115 1.850 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.150 1.145 2.380 1.375 ;
        RECT  2.030 0.885 2.150 1.375 ;
        RECT  1.790 1.145 2.030 1.375 ;
        RECT  1.670 0.885 1.790 1.375 ;
        RECT  1.430 1.145 1.670 1.375 ;
        RECT  1.310 0.885 1.430 1.375 ;
        RECT  1.070 1.145 1.310 1.375 ;
        RECT  0.950 0.885 1.070 1.375 ;
        RECT  0.710 1.145 0.950 1.375 ;
        RECT  0.590 1.030 0.710 1.375 ;
        RECT  0.350 1.145 0.590 1.375 ;
        RECT  0.230 1.030 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.230 0.700 2.310 1.035 ;
        RECT  1.950 0.700 2.230 0.815 ;
        RECT  1.870 0.700 1.950 1.035 ;
        RECT  1.590 0.700 1.870 0.815 ;
        RECT  1.510 0.700 1.590 1.035 ;
        RECT  1.230 0.700 1.510 0.815 ;
        RECT  1.150 0.700 1.230 1.035 ;
        RECT  0.870 0.700 1.150 0.815 ;
        RECT  0.790 0.700 0.870 1.035 ;
        RECT  0.785 0.700 0.790 0.960 ;
        RECT  0.665 0.845 0.785 0.960 ;
        RECT  0.160 0.355 0.315 0.425 ;
        RECT  0.150 0.845 0.315 0.960 ;
        RECT  0.060 0.185 0.160 0.425 ;
        RECT  0.070 0.845 0.150 1.035 ;
        RECT  2.040 0.185 2.140 0.425 ;
        RECT  1.770 0.355 2.040 0.425 ;
        RECT  1.690 0.215 1.770 0.425 ;
        RECT  1.310 0.215 1.690 0.285 ;
        RECT  1.230 0.355 1.610 0.425 ;
        RECT  1.150 0.190 1.230 0.425 ;
        RECT  0.750 0.355 1.150 0.425 ;
        RECT  0.230 0.205 1.070 0.275 ;
    END
END ND4D3BWP

MACRO ND4D4BWP
    CLASS CORE ;
    FOREIGN ND4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.055 0.700 3.125 1.020 ;
        RECT  2.705 0.700 3.055 0.815 ;
        RECT  2.635 0.700 2.705 1.020 ;
        RECT  2.285 0.700 2.635 0.815 ;
        RECT  2.215 0.700 2.285 1.020 ;
        RECT  1.925 0.700 2.215 0.815 ;
        RECT  1.855 0.700 1.925 1.020 ;
        RECT  1.385 0.700 1.855 0.815 ;
        RECT  1.315 0.700 1.385 1.020 ;
        RECT  1.025 0.700 1.315 0.815 ;
        RECT  0.955 0.700 1.025 1.020 ;
        RECT  0.665 0.700 0.955 0.815 ;
        RECT  0.595 0.345 0.690 0.430 ;
        RECT  0.595 0.700 0.665 1.020 ;
        RECT  0.385 0.345 0.595 0.815 ;
        RECT  0.210 0.345 0.385 0.430 ;
        RECT  0.305 0.700 0.385 0.815 ;
        RECT  0.235 0.700 0.305 1.020 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.495 3.070 0.630 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.495 2.345 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.390 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.120 -0.115 3.360 0.115 ;
        RECT  3.000 -0.115 3.120 0.275 ;
        RECT  2.700 -0.115 3.000 0.115 ;
        RECT  2.580 -0.115 2.700 0.275 ;
        RECT  0.000 -0.115 2.580 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.145 3.360 1.375 ;
        RECT  3.235 0.680 3.305 1.375 ;
        RECT  2.940 1.145 3.235 1.375 ;
        RECT  2.820 0.885 2.940 1.375 ;
        RECT  2.520 1.145 2.820 1.375 ;
        RECT  2.400 0.885 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 0.885 2.130 1.375 ;
        RECT  1.750 1.145 2.010 1.375 ;
        RECT  1.670 0.885 1.750 1.375 ;
        RECT  1.570 1.145 1.670 1.375 ;
        RECT  1.490 0.885 1.570 1.375 ;
        RECT  1.230 1.145 1.490 1.375 ;
        RECT  1.110 0.885 1.230 1.375 ;
        RECT  0.870 1.145 1.110 1.375 ;
        RECT  0.750 0.885 0.870 1.375 ;
        RECT  0.510 1.145 0.750 1.375 ;
        RECT  0.390 0.885 0.510 1.375 ;
        RECT  0.140 1.145 0.390 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.055 0.700 3.125 1.020 ;
        RECT  2.705 0.700 3.055 0.815 ;
        RECT  2.635 0.700 2.705 1.020 ;
        RECT  2.285 0.700 2.635 0.815 ;
        RECT  2.215 0.700 2.285 1.020 ;
        RECT  1.925 0.700 2.215 0.815 ;
        RECT  1.855 0.700 1.925 1.020 ;
        RECT  1.385 0.700 1.855 0.815 ;
        RECT  1.315 0.700 1.385 1.020 ;
        RECT  1.025 0.700 1.315 0.815 ;
        RECT  0.955 0.700 1.025 1.020 ;
        RECT  0.665 0.700 0.955 0.815 ;
        RECT  0.665 0.345 0.690 0.430 ;
        RECT  0.210 0.345 0.315 0.430 ;
        RECT  0.305 0.700 0.315 0.815 ;
        RECT  0.235 0.700 0.305 1.020 ;
        RECT  3.220 0.185 3.320 0.430 ;
        RECT  2.890 0.355 3.220 0.425 ;
        RECT  2.810 0.190 2.890 0.425 ;
        RECT  2.470 0.355 2.810 0.425 ;
        RECT  2.390 0.190 2.470 0.425 ;
        RECT  1.650 0.355 2.390 0.425 ;
        RECT  0.930 0.205 2.310 0.275 ;
        RECT  1.490 0.345 1.570 0.470 ;
        RECT  0.845 0.345 1.490 0.415 ;
        RECT  0.775 0.205 0.845 0.415 ;
        RECT  0.130 0.205 0.775 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END ND4D4BWP

MACRO ND4D8BWP
    CLASS CORE ;
    FOREIGN ND4D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.690 2.190 0.810 ;
        RECT  2.095 0.185 2.165 0.465 ;
        RECT  1.805 0.345 2.095 0.465 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.575 0.345 1.735 0.465 ;
        RECT  1.445 0.345 1.575 0.810 ;
        RECT  1.375 0.185 1.445 0.810 ;
        RECT  1.365 0.345 1.375 0.810 ;
        RECT  1.085 0.345 1.365 0.465 ;
        RECT  1.015 0.690 1.365 0.810 ;
        RECT  1.015 0.185 1.085 0.465 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.805 0.790 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.475 0.385 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.940 0.115 ;
        RECT  2.630 -0.115 2.710 0.315 ;
        RECT  2.350 -0.115 2.630 0.115 ;
        RECT  2.270 -0.115 2.350 0.315 ;
        RECT  2.010 -0.115 2.270 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  1.650 -0.115 1.890 0.115 ;
        RECT  1.530 -0.115 1.650 0.275 ;
        RECT  1.290 -0.115 1.530 0.115 ;
        RECT  1.170 -0.115 1.290 0.265 ;
        RECT  0.900 -0.115 1.170 0.115 ;
        RECT  0.780 -0.115 0.900 0.245 ;
        RECT  0.000 -0.115 0.780 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.145 2.940 1.375 ;
        RECT  2.610 0.980 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.020 2.370 1.375 ;
        RECT  2.010 1.145 2.250 1.375 ;
        RECT  1.890 1.020 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.020 1.650 1.375 ;
        RECT  1.290 1.145 1.530 1.375 ;
        RECT  1.170 1.020 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 1.020 0.910 1.375 ;
        RECT  0.510 1.145 0.790 1.375 ;
        RECT  0.390 1.020 0.510 1.375 ;
        RECT  0.120 1.145 0.390 1.375 ;
        RECT  0.050 0.800 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.690 2.190 0.810 ;
        RECT  2.095 0.185 2.165 0.465 ;
        RECT  1.805 0.345 2.095 0.465 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.645 0.345 1.735 0.465 ;
        RECT  1.085 0.345 1.295 0.465 ;
        RECT  1.015 0.690 1.295 0.810 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  2.810 0.185 2.890 1.070 ;
        RECT  2.530 0.395 2.810 0.465 ;
        RECT  2.540 0.830 2.810 0.900 ;
        RECT  2.480 0.540 2.620 0.620 ;
        RECT  2.440 0.830 2.540 1.070 ;
        RECT  2.450 0.185 2.530 0.465 ;
        RECT  2.410 0.540 2.480 0.760 ;
        RECT  2.325 0.395 2.450 0.465 ;
        RECT  2.335 0.690 2.410 0.760 ;
        RECT  2.265 0.690 2.335 0.950 ;
        RECT  2.255 0.395 2.325 0.610 ;
        RECT  0.945 0.880 2.265 0.950 ;
        RECT  1.685 0.540 2.255 0.610 ;
        RECT  0.875 0.315 0.945 0.950 ;
        RECT  0.295 0.315 0.875 0.395 ;
        RECT  0.200 0.880 0.875 0.950 ;
        RECT  0.215 0.185 0.295 0.395 ;
        RECT  0.040 0.185 0.215 0.285 ;
    END
END ND4D8BWP

MACRO NR2D0BWP
    CLASS CORE ;
    FOREIGN NR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0474 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.345 0.525 1.065 ;
        RECT  0.315 0.345 0.455 0.415 ;
        RECT  0.435 0.925 0.455 1.065 ;
        RECT  0.245 0.185 0.315 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.115 0.560 0.115 ;
        RECT  0.420 -0.115 0.520 0.275 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.145 0.560 1.375 ;
        RECT  0.050 0.925 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END NR2D0BWP

MACRO NR2D1BWP
    CLASS CORE ;
    FOREIGN NR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0947 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.355 0.525 1.045 ;
        RECT  0.315 0.355 0.455 0.425 ;
        RECT  0.435 0.915 0.455 1.045 ;
        RECT  0.245 0.210 0.315 0.425 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.195 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.280 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.145 0.560 1.375 ;
        RECT  0.050 0.820 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END NR2D1BWP

MACRO NR2D2BWP
    CLASS CORE ;
    FOREIGN NR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1442 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.660 0.185 0.760 0.425 ;
        RECT  0.385 0.355 0.660 0.425 ;
        RECT  0.340 0.355 0.385 0.920 ;
        RECT  0.315 0.185 0.340 0.920 ;
        RECT  0.240 0.185 0.315 0.430 ;
        RECT  0.230 0.710 0.315 0.920 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.670 0.495 0.735 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.940 0.415 ;
        RECT  0.540 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.540 0.285 ;
        RECT  0.160 -0.115 0.460 0.115 ;
        RECT  0.055 -0.115 0.160 0.275 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.640 0.975 0.720 1.375 ;
        RECT  0.000 1.145 0.640 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.835 0.930 0.955 ;
        RECT  0.560 0.835 0.850 0.905 ;
        RECT  0.490 0.835 0.560 1.065 ;
        RECT  0.150 0.995 0.490 1.065 ;
        RECT  0.070 0.735 0.150 1.065 ;
    END
END NR2D2BWP

MACRO NR2D3BWP
    CLASS CORE ;
    FOREIGN NR2D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2327 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.215 1.050 0.425 ;
        RECT  0.680 0.355 0.930 0.425 ;
        RECT  0.580 0.190 0.680 0.425 ;
        RECT  0.525 0.355 0.580 0.425 ;
        RECT  0.455 0.355 0.525 0.905 ;
        RECT  0.330 0.355 0.455 0.425 ;
        RECT  0.125 0.835 0.455 0.905 ;
        RECT  0.210 0.215 0.330 0.425 ;
        RECT  0.055 0.835 0.125 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.545 1.040 0.625 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.470 ;
        RECT  0.850 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.850 0.285 ;
        RECT  0.490 -0.115 0.770 0.115 ;
        RECT  0.410 -0.115 0.490 0.285 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.680 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.975 0.850 1.375 ;
        RECT  0.000 1.145 0.770 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.835 1.030 0.995 ;
        RECT  0.665 0.835 0.950 0.905 ;
        RECT  0.595 0.835 0.665 1.065 ;
        RECT  0.210 0.995 0.595 1.065 ;
    END
END NR2D3BWP

MACRO NR2D4BWP
    CLASS CORE ;
    FOREIGN NR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2884 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.765 1.460 0.895 ;
        RECT  1.355 0.235 1.425 0.415 ;
        RECT  1.295 0.345 1.355 0.415 ;
        RECT  1.085 0.345 1.295 0.895 ;
        RECT  1.070 0.345 1.085 0.415 ;
        RECT  0.970 0.765 1.085 0.895 ;
        RECT  0.990 0.185 1.070 0.415 ;
        RECT  0.690 0.345 0.990 0.415 ;
        RECT  0.610 0.185 0.690 0.415 ;
        RECT  0.325 0.345 0.610 0.415 ;
        RECT  0.255 0.235 0.325 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 0.495 0.665 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.390 0.495 1.575 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 -0.115 1.680 0.115 ;
        RECT  1.530 -0.115 1.610 0.395 ;
        RECT  1.260 -0.115 1.530 0.115 ;
        RECT  1.160 -0.115 1.260 0.275 ;
        RECT  0.890 -0.115 1.160 0.115 ;
        RECT  0.790 -0.115 0.890 0.275 ;
        RECT  0.520 -0.115 0.790 0.115 ;
        RECT  0.420 -0.115 0.520 0.275 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.070 -0.115 0.150 0.395 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.145 1.680 1.375 ;
        RECT  0.610 0.845 0.690 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.250 0.845 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.765 1.460 0.895 ;
        RECT  1.365 0.235 1.425 0.415 ;
        RECT  0.990 0.185 1.015 0.415 ;
        RECT  0.970 0.765 1.015 0.895 ;
        RECT  0.690 0.345 0.990 0.415 ;
        RECT  0.610 0.185 0.690 0.415 ;
        RECT  0.325 0.345 0.610 0.415 ;
        RECT  0.255 0.235 0.325 0.415 ;
        RECT  1.530 0.865 1.610 1.045 ;
        RECT  0.880 0.975 1.530 1.045 ;
        RECT  0.800 0.705 0.880 1.045 ;
        RECT  0.510 0.705 0.800 0.775 ;
        RECT  0.430 0.705 0.510 1.035 ;
        RECT  0.150 0.705 0.430 0.775 ;
        RECT  0.070 0.705 0.150 1.035 ;
    END
END NR2D4BWP

MACRO NR2D8BWP
    CLASS CORE ;
    FOREIGN NR2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5768 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.750 0.210 2.870 0.415 ;
        RECT  2.415 0.775 2.870 0.905 ;
        RECT  2.490 0.345 2.750 0.415 ;
        RECT  2.415 0.185 2.490 0.415 ;
        RECT  2.410 0.185 2.415 0.905 ;
        RECT  2.205 0.345 2.410 0.905 ;
        RECT  2.130 0.345 2.205 0.415 ;
        RECT  1.670 0.775 2.205 0.905 ;
        RECT  2.050 0.185 2.130 0.415 ;
        RECT  1.770 0.345 2.050 0.415 ;
        RECT  1.690 0.185 1.770 0.415 ;
        RECT  1.410 0.345 1.690 0.415 ;
        RECT  1.330 0.185 1.410 0.415 ;
        RECT  1.050 0.345 1.330 0.415 ;
        RECT  0.970 0.185 1.050 0.415 ;
        RECT  0.690 0.345 0.970 0.415 ;
        RECT  0.610 0.185 0.690 0.415 ;
        RECT  0.350 0.345 0.610 0.415 ;
        RECT  0.230 0.210 0.350 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 1.385 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 0.495 2.100 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.465 ;
        RECT  2.680 -0.115 2.950 0.115 ;
        RECT  2.580 -0.115 2.680 0.275 ;
        RECT  2.320 -0.115 2.580 0.115 ;
        RECT  2.220 -0.115 2.320 0.275 ;
        RECT  1.960 -0.115 2.220 0.115 ;
        RECT  1.860 -0.115 1.960 0.275 ;
        RECT  1.600 -0.115 1.860 0.115 ;
        RECT  1.500 -0.115 1.600 0.275 ;
        RECT  1.240 -0.115 1.500 0.115 ;
        RECT  1.140 -0.115 1.240 0.275 ;
        RECT  0.880 -0.115 1.140 0.115 ;
        RECT  0.780 -0.115 0.880 0.275 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.420 -0.115 0.520 0.275 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.070 -0.115 0.150 0.465 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.145 3.080 1.375 ;
        RECT  1.330 0.845 1.410 1.375 ;
        RECT  1.050 1.145 1.330 1.375 ;
        RECT  0.970 0.845 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.845 0.690 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.250 0.845 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.210 2.870 0.415 ;
        RECT  2.485 0.775 2.870 0.905 ;
        RECT  2.490 0.345 2.750 0.415 ;
        RECT  2.485 0.185 2.490 0.415 ;
        RECT  2.130 0.345 2.135 0.415 ;
        RECT  1.670 0.775 2.135 0.905 ;
        RECT  2.050 0.185 2.130 0.415 ;
        RECT  1.770 0.345 2.050 0.415 ;
        RECT  1.690 0.185 1.770 0.415 ;
        RECT  1.410 0.345 1.690 0.415 ;
        RECT  1.330 0.185 1.410 0.415 ;
        RECT  1.050 0.345 1.330 0.415 ;
        RECT  0.970 0.185 1.050 0.415 ;
        RECT  0.690 0.345 0.970 0.415 ;
        RECT  0.610 0.185 0.690 0.415 ;
        RECT  0.350 0.345 0.610 0.415 ;
        RECT  0.230 0.210 0.350 0.415 ;
        RECT  2.950 0.735 3.030 1.045 ;
        RECT  1.590 0.975 2.950 1.045 ;
        RECT  2.640 0.540 2.920 0.625 ;
        RECT  1.510 0.705 1.590 1.045 ;
        RECT  1.230 0.705 1.510 0.775 ;
        RECT  1.150 0.705 1.230 1.035 ;
        RECT  0.870 0.705 1.150 0.775 ;
        RECT  0.790 0.705 0.870 1.035 ;
        RECT  0.510 0.705 0.790 0.775 ;
        RECT  0.430 0.705 0.510 1.035 ;
        RECT  0.150 0.705 0.430 0.775 ;
        RECT  0.070 0.705 0.150 1.035 ;
    END
END NR2D8BWP

MACRO NR2XD0BWP
    CLASS CORE ;
    FOREIGN NR2XD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0699 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.340 0.525 1.075 ;
        RECT  0.315 0.340 0.455 0.410 ;
        RECT  0.420 0.835 0.455 1.075 ;
        RECT  0.245 0.185 0.315 0.410 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 -0.115 0.560 0.115 ;
        RECT  0.420 -0.115 0.520 0.270 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.145 0.560 1.375 ;
        RECT  0.050 0.815 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END NR2XD0BWP

MACRO NR2XD1BWP
    CLASS CORE ;
    FOREIGN NR2XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.715 0.710 0.925 ;
        RECT  0.590 0.355 0.665 0.925 ;
        RECT  0.540 0.355 0.590 0.425 ;
        RECT  0.440 0.185 0.540 0.425 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.385 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.625 ;
        RECT  0.735 0.545 0.875 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 -0.115 0.980 0.115 ;
        RECT  0.630 -0.115 0.710 0.285 ;
        RECT  0.350 -0.115 0.630 0.115 ;
        RECT  0.260 -0.115 0.350 0.440 ;
        RECT  0.000 -0.115 0.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.250 0.845 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.795 0.735 0.865 1.065 ;
        RECT  0.505 0.995 0.795 1.065 ;
        RECT  0.435 0.705 0.505 1.065 ;
        RECT  0.150 0.705 0.435 0.775 ;
        RECT  0.070 0.705 0.150 1.035 ;
    END
END NR2XD1BWP

MACRO NR2XD2BWP
    CLASS CORE ;
    FOREIGN NR2XD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.845 1.450 0.915 ;
        RECT  1.355 0.200 1.435 0.415 ;
        RECT  1.085 0.325 1.355 0.415 ;
        RECT  1.065 0.325 1.085 0.915 ;
        RECT  1.015 0.200 1.065 0.915 ;
        RECT  0.995 0.200 1.015 0.415 ;
        RECT  0.970 0.845 1.015 0.915 ;
        RECT  0.705 0.325 0.995 0.415 ;
        RECT  0.635 0.200 0.705 0.415 ;
        RECT  0.325 0.325 0.635 0.415 ;
        RECT  0.255 0.200 0.325 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.700 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.495 1.515 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 -0.115 1.680 0.115 ;
        RECT  1.530 -0.115 1.610 0.330 ;
        RECT  1.270 -0.115 1.530 0.115 ;
        RECT  1.150 -0.115 1.270 0.255 ;
        RECT  0.910 -0.115 1.150 0.115 ;
        RECT  0.790 -0.115 0.910 0.255 ;
        RECT  0.540 -0.115 0.790 0.115 ;
        RECT  0.420 -0.115 0.540 0.255 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.070 -0.115 0.150 0.320 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.145 1.680 1.375 ;
        RECT  0.630 0.845 0.710 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.260 0.845 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.895 1.605 1.055 ;
        RECT  0.885 0.985 1.535 1.055 ;
        RECT  0.815 0.705 0.885 1.055 ;
        RECT  0.525 0.705 0.815 0.775 ;
        RECT  0.455 0.705 0.525 1.055 ;
        RECT  0.145 0.705 0.455 0.775 ;
        RECT  0.075 0.705 0.145 1.035 ;
    END
END NR2XD2BWP

MACRO NR2XD3BWP
    CLASS CORE ;
    FOREIGN NR2XD3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3024 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.695 2.170 0.815 ;
        RECT  2.070 0.190 2.150 0.415 ;
        RECT  1.785 0.335 2.070 0.415 ;
        RECT  1.715 0.190 1.785 0.415 ;
        RECT  1.435 0.335 1.715 0.415 ;
        RECT  1.425 0.335 1.435 0.815 ;
        RECT  1.355 0.190 1.425 0.815 ;
        RECT  1.225 0.335 1.355 0.815 ;
        RECT  1.065 0.335 1.225 0.415 ;
        RECT  0.995 0.190 1.065 0.415 ;
        RECT  0.685 0.335 0.995 0.415 ;
        RECT  0.615 0.190 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.190 0.305 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 1.085 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 2.345 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.330 ;
        RECT  1.990 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.990 0.265 ;
        RECT  1.630 -0.115 1.870 0.115 ;
        RECT  1.510 -0.115 1.630 0.265 ;
        RECT  1.270 -0.115 1.510 0.115 ;
        RECT  1.150 -0.115 1.270 0.265 ;
        RECT  0.900 -0.115 1.150 0.115 ;
        RECT  0.780 -0.115 0.900 0.265 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.265 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.330 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.145 2.380 1.375 ;
        RECT  0.960 1.025 1.080 1.375 ;
        RECT  0.685 1.145 0.960 1.375 ;
        RECT  0.615 0.860 0.685 1.375 ;
        RECT  0.315 1.145 0.615 1.375 ;
        RECT  0.245 0.860 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.695 2.170 0.815 ;
        RECT  2.070 0.190 2.150 0.415 ;
        RECT  1.785 0.335 2.070 0.415 ;
        RECT  1.715 0.190 1.785 0.415 ;
        RECT  1.505 0.335 1.715 0.415 ;
        RECT  1.065 0.335 1.155 0.415 ;
        RECT  0.995 0.190 1.065 0.415 ;
        RECT  0.685 0.335 0.995 0.415 ;
        RECT  0.615 0.190 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.190 0.305 0.415 ;
        RECT  2.255 0.885 2.325 1.005 ;
        RECT  0.865 0.885 2.255 0.955 ;
        RECT  0.795 0.715 0.865 1.035 ;
        RECT  0.505 0.715 0.795 0.785 ;
        RECT  0.435 0.715 0.505 1.035 ;
        RECT  0.125 0.715 0.435 0.790 ;
        RECT  0.055 0.715 0.125 1.055 ;
    END
END NR2XD3BWP

MACRO NR2XD4BWP
    CLASS CORE ;
    FOREIGN NR2XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.775 2.850 0.905 ;
        RECT  2.775 0.195 2.845 0.415 ;
        RECT  2.485 0.335 2.775 0.415 ;
        RECT  2.415 0.195 2.485 0.415 ;
        RECT  2.125 0.335 2.415 0.415 ;
        RECT  2.055 0.195 2.125 0.415 ;
        RECT  1.995 0.335 2.055 0.415 ;
        RECT  1.785 0.335 1.995 0.905 ;
        RECT  1.765 0.335 1.785 0.415 ;
        RECT  1.690 0.775 1.785 0.905 ;
        RECT  1.695 0.195 1.765 0.415 ;
        RECT  1.405 0.335 1.695 0.415 ;
        RECT  1.335 0.190 1.405 0.415 ;
        RECT  1.045 0.335 1.335 0.415 ;
        RECT  0.975 0.190 1.045 0.415 ;
        RECT  0.685 0.335 0.975 0.415 ;
        RECT  0.615 0.195 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.195 0.305 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 1.400 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 3.045 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.305 ;
        RECT  2.690 -0.115 2.950 0.115 ;
        RECT  2.570 -0.115 2.690 0.265 ;
        RECT  2.330 -0.115 2.570 0.115 ;
        RECT  2.210 -0.115 2.330 0.265 ;
        RECT  1.970 -0.115 2.210 0.115 ;
        RECT  1.850 -0.115 1.970 0.265 ;
        RECT  1.610 -0.115 1.850 0.115 ;
        RECT  1.490 -0.115 1.610 0.265 ;
        RECT  1.250 -0.115 1.490 0.115 ;
        RECT  1.130 -0.115 1.250 0.265 ;
        RECT  0.890 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.890 0.265 ;
        RECT  0.520 -0.115 0.770 0.115 ;
        RECT  0.400 -0.115 0.520 0.265 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.145 3.080 1.375 ;
        RECT  1.330 0.855 1.410 1.375 ;
        RECT  1.050 1.145 1.330 1.375 ;
        RECT  0.970 0.855 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.855 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.855 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.065 0.775 2.850 0.905 ;
        RECT  2.775 0.195 2.845 0.415 ;
        RECT  2.485 0.335 2.775 0.415 ;
        RECT  2.415 0.195 2.485 0.415 ;
        RECT  2.125 0.335 2.415 0.415 ;
        RECT  2.065 0.195 2.125 0.415 ;
        RECT  1.695 0.195 1.715 0.415 ;
        RECT  1.690 0.775 1.715 0.905 ;
        RECT  1.405 0.335 1.695 0.415 ;
        RECT  1.335 0.190 1.405 0.415 ;
        RECT  1.045 0.335 1.335 0.415 ;
        RECT  0.975 0.190 1.045 0.415 ;
        RECT  0.685 0.335 0.975 0.415 ;
        RECT  0.615 0.195 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.195 0.305 0.415 ;
        RECT  2.955 0.735 3.025 1.055 ;
        RECT  1.585 0.985 2.955 1.055 ;
        RECT  1.515 0.715 1.585 1.055 ;
        RECT  1.225 0.715 1.515 0.785 ;
        RECT  1.155 0.715 1.225 1.035 ;
        RECT  0.865 0.715 1.155 0.785 ;
        RECT  0.795 0.715 0.865 1.035 ;
        RECT  0.505 0.715 0.795 0.785 ;
        RECT  0.435 0.715 0.505 1.035 ;
        RECT  0.125 0.715 0.435 0.785 ;
        RECT  0.055 0.715 0.125 1.035 ;
    END
END NR2XD4BWP

MACRO NR2XD8BWP
    CLASS CORE ;
    FOREIGN NR2XD8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.8064 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.745 5.790 0.865 ;
        RECT  5.715 0.195 5.785 0.415 ;
        RECT  5.425 0.335 5.715 0.415 ;
        RECT  5.355 0.195 5.425 0.415 ;
        RECT  5.065 0.335 5.355 0.415 ;
        RECT  4.995 0.195 5.065 0.415 ;
        RECT  4.705 0.335 4.995 0.415 ;
        RECT  4.635 0.195 4.705 0.415 ;
        RECT  4.345 0.335 4.635 0.415 ;
        RECT  4.275 0.195 4.345 0.415 ;
        RECT  3.985 0.335 4.275 0.415 ;
        RECT  3.915 0.195 3.985 0.415 ;
        RECT  3.675 0.335 3.915 0.415 ;
        RECT  3.625 0.335 3.675 0.865 ;
        RECT  3.555 0.195 3.625 0.865 ;
        RECT  3.465 0.335 3.555 0.865 ;
        RECT  3.265 0.335 3.465 0.415 ;
        RECT  3.190 0.745 3.465 0.865 ;
        RECT  3.195 0.195 3.265 0.415 ;
        RECT  2.905 0.335 3.195 0.415 ;
        RECT  2.835 0.195 2.905 0.415 ;
        RECT  2.525 0.335 2.835 0.415 ;
        RECT  2.455 0.195 2.525 0.415 ;
        RECT  2.145 0.335 2.455 0.415 ;
        RECT  2.075 0.195 2.145 0.415 ;
        RECT  1.785 0.335 2.075 0.415 ;
        RECT  1.715 0.195 1.785 0.415 ;
        RECT  1.405 0.335 1.715 0.415 ;
        RECT  1.335 0.195 1.405 0.415 ;
        RECT  1.045 0.335 1.335 0.415 ;
        RECT  0.975 0.195 1.045 0.415 ;
        RECT  0.685 0.335 0.975 0.415 ;
        RECT  0.615 0.195 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.195 0.305 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.3616 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 2.850 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3616 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.900 0.495 5.985 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 -0.115 6.020 0.115 ;
        RECT  5.890 -0.115 5.970 0.325 ;
        RECT  5.630 -0.115 5.890 0.115 ;
        RECT  5.510 -0.115 5.630 0.265 ;
        RECT  5.270 -0.115 5.510 0.115 ;
        RECT  5.150 -0.115 5.270 0.265 ;
        RECT  4.910 -0.115 5.150 0.115 ;
        RECT  4.790 -0.115 4.910 0.265 ;
        RECT  4.550 -0.115 4.790 0.115 ;
        RECT  4.430 -0.115 4.550 0.265 ;
        RECT  4.190 -0.115 4.430 0.115 ;
        RECT  4.070 -0.115 4.190 0.265 ;
        RECT  3.830 -0.115 4.070 0.115 ;
        RECT  3.710 -0.115 3.830 0.265 ;
        RECT  3.470 -0.115 3.710 0.115 ;
        RECT  3.350 -0.115 3.470 0.265 ;
        RECT  3.110 -0.115 3.350 0.115 ;
        RECT  2.990 -0.115 3.110 0.265 ;
        RECT  2.740 -0.115 2.990 0.115 ;
        RECT  2.620 -0.115 2.740 0.265 ;
        RECT  2.360 -0.115 2.620 0.115 ;
        RECT  2.240 -0.115 2.360 0.265 ;
        RECT  1.990 -0.115 2.240 0.115 ;
        RECT  1.870 -0.115 1.990 0.265 ;
        RECT  1.620 -0.115 1.870 0.115 ;
        RECT  1.500 -0.115 1.620 0.265 ;
        RECT  1.250 -0.115 1.500 0.115 ;
        RECT  1.130 -0.115 1.250 0.265 ;
        RECT  0.890 -0.115 1.130 0.115 ;
        RECT  0.770 -0.115 0.890 0.265 ;
        RECT  0.520 -0.115 0.770 0.115 ;
        RECT  0.400 -0.115 0.520 0.265 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.325 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 6.020 1.375 ;
        RECT  2.820 0.845 2.900 1.375 ;
        RECT  2.520 1.145 2.820 1.375 ;
        RECT  2.440 0.845 2.520 1.375 ;
        RECT  2.140 1.145 2.440 1.375 ;
        RECT  2.060 0.845 2.140 1.375 ;
        RECT  1.770 1.145 2.060 1.375 ;
        RECT  1.690 0.845 1.770 1.375 ;
        RECT  1.410 1.145 1.690 1.375 ;
        RECT  1.330 0.845 1.410 1.375 ;
        RECT  1.050 1.145 1.330 1.375 ;
        RECT  0.970 0.845 1.050 1.375 ;
        RECT  0.690 1.145 0.970 1.375 ;
        RECT  0.610 0.845 0.690 1.375 ;
        RECT  0.320 1.145 0.610 1.375 ;
        RECT  0.240 0.845 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.745 5.790 0.865 ;
        RECT  5.715 0.195 5.785 0.415 ;
        RECT  5.425 0.335 5.715 0.415 ;
        RECT  5.355 0.195 5.425 0.415 ;
        RECT  5.065 0.335 5.355 0.415 ;
        RECT  4.995 0.195 5.065 0.415 ;
        RECT  4.705 0.335 4.995 0.415 ;
        RECT  4.635 0.195 4.705 0.415 ;
        RECT  4.345 0.335 4.635 0.415 ;
        RECT  4.275 0.195 4.345 0.415 ;
        RECT  3.985 0.335 4.275 0.415 ;
        RECT  3.915 0.195 3.985 0.415 ;
        RECT  3.745 0.335 3.915 0.415 ;
        RECT  3.265 0.335 3.395 0.415 ;
        RECT  3.190 0.745 3.395 0.865 ;
        RECT  3.195 0.195 3.265 0.415 ;
        RECT  2.905 0.335 3.195 0.415 ;
        RECT  2.835 0.195 2.905 0.415 ;
        RECT  2.525 0.335 2.835 0.415 ;
        RECT  2.455 0.195 2.525 0.415 ;
        RECT  2.145 0.335 2.455 0.415 ;
        RECT  2.075 0.195 2.145 0.415 ;
        RECT  1.785 0.335 2.075 0.415 ;
        RECT  1.715 0.195 1.785 0.415 ;
        RECT  1.405 0.335 1.715 0.415 ;
        RECT  1.335 0.195 1.405 0.415 ;
        RECT  1.045 0.335 1.335 0.415 ;
        RECT  0.975 0.195 1.045 0.415 ;
        RECT  0.685 0.335 0.975 0.415 ;
        RECT  0.615 0.195 0.685 0.415 ;
        RECT  0.305 0.335 0.615 0.415 ;
        RECT  0.235 0.195 0.305 0.415 ;
        RECT  5.895 0.735 5.965 1.055 ;
        RECT  3.085 0.985 5.895 1.055 ;
        RECT  3.015 0.705 3.085 1.055 ;
        RECT  2.705 0.705 3.015 0.775 ;
        RECT  2.635 0.705 2.705 1.035 ;
        RECT  2.330 0.705 2.635 0.775 ;
        RECT  2.255 0.705 2.330 1.035 ;
        RECT  1.950 0.705 2.255 0.775 ;
        RECT  1.875 0.705 1.950 1.035 ;
        RECT  1.590 0.705 1.875 0.775 ;
        RECT  1.510 0.705 1.590 1.035 ;
        RECT  1.225 0.705 1.510 0.775 ;
        RECT  1.155 0.705 1.225 1.035 ;
        RECT  0.865 0.705 1.155 0.775 ;
        RECT  0.795 0.705 0.865 1.035 ;
        RECT  0.505 0.705 0.795 0.775 ;
        RECT  0.435 0.705 0.505 1.035 ;
        RECT  0.125 0.705 0.435 0.775 ;
        RECT  0.055 0.705 0.125 1.035 ;
    END
END NR2XD8BWP

MACRO NR3D0BWP
    CLASS CORE ;
    FOREIGN NR3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0838 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.205 0.805 1.075 ;
        RECT  0.715 0.205 0.735 0.415 ;
        RECT  0.700 0.835 0.735 1.075 ;
        RECT  0.385 0.345 0.715 0.415 ;
        RECT  0.295 0.205 0.385 0.415 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 -0.115 0.840 0.115 ;
        RECT  0.470 -0.115 0.610 0.275 ;
        RECT  0.200 -0.115 0.470 0.115 ;
        RECT  0.100 -0.115 0.200 0.280 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.145 0.840 1.375 ;
        RECT  0.040 0.705 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END NR3D0BWP

MACRO NR3D1BWP
    CLASS CORE ;
    FOREIGN NR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1677 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.205 1.225 1.070 ;
        RECT  0.120 0.205 1.155 0.275 ;
        RECT  1.135 0.670 1.155 1.070 ;
        RECT  0.125 0.890 1.135 0.960 ;
        RECT  0.035 0.890 0.125 1.055 ;
        RECT  0.035 0.205 0.120 0.345 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.355 0.900 0.425 ;
        RECT  0.455 0.355 0.525 0.640 ;
        RECT  0.315 0.520 0.455 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.355 1.085 0.510 ;
        RECT  0.985 0.355 1.055 0.820 ;
        RECT  0.245 0.750 0.985 0.820 ;
        RECT  0.170 0.495 0.245 0.820 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.145 1.260 1.375 ;
        RECT  0.570 1.030 0.690 1.375 ;
        RECT  0.000 1.145 0.570 1.375 ;
        END
    END VDD
END NR3D1BWP

MACRO NR3D2BWP
    CLASS CORE ;
    FOREIGN NR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2530 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.210 2.205 0.370 ;
        RECT  1.925 0.300 2.115 0.370 ;
        RECT  1.925 0.855 2.030 0.925 ;
        RECT  1.855 0.300 1.925 0.925 ;
        RECT  1.605 0.300 1.855 0.370 ;
        RECT  1.550 0.855 1.855 0.925 ;
        RECT  1.535 0.215 1.605 0.370 ;
        RECT  1.245 0.300 1.535 0.370 ;
        RECT  1.175 0.215 1.245 0.370 ;
        RECT  0.885 0.300 1.175 0.370 ;
        RECT  0.815 0.215 0.885 0.370 ;
        RECT  0.305 0.300 0.815 0.370 ;
        RECT  0.235 0.210 0.305 0.370 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.450 0.665 0.520 ;
        RECT  0.315 0.450 0.385 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.450 1.225 0.625 ;
        RECT  0.875 0.450 1.015 0.520 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.450 1.785 0.765 ;
        RECT  1.435 0.450 1.715 0.520 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 -0.115 2.240 0.115 ;
        RECT  1.910 -0.115 2.030 0.220 ;
        RECT  0.510 -0.115 1.910 0.115 ;
        RECT  0.390 -0.115 0.510 0.220 ;
        RECT  0.130 -0.115 0.390 0.115 ;
        RECT  0.050 -0.115 0.130 0.365 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.145 2.240 1.375 ;
        RECT  0.610 0.845 0.690 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.110 0.910 2.190 1.065 ;
        RECT  1.440 0.995 2.110 1.065 ;
        RECT  1.360 0.680 1.440 1.065 ;
        RECT  1.070 0.995 1.360 1.065 ;
        RECT  1.140 0.705 1.250 0.925 ;
        RECT  0.870 0.705 1.140 0.775 ;
        RECT  0.950 0.855 1.070 1.065 ;
        RECT  0.790 0.705 0.870 1.000 ;
        RECT  0.530 0.705 0.790 0.775 ;
        RECT  0.455 0.705 0.530 1.050 ;
        RECT  0.430 0.845 0.455 1.050 ;
        RECT  0.130 0.845 0.430 0.915 ;
        RECT  0.050 0.845 0.130 1.050 ;
    END
END NR3D2BWP

MACRO NR3D3BWP
    CLASS CORE ;
    FOREIGN NR3D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3743 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.775 3.160 0.905 ;
        RECT  2.555 0.205 3.105 0.325 ;
        RECT  2.335 0.205 2.555 0.905 ;
        RECT  0.275 0.205 2.335 0.325 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.435 1.090 0.625 ;
        RECT  0.290 0.435 0.875 0.530 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.435 2.065 0.625 ;
        RECT  1.435 0.435 1.855 0.530 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.435 3.325 0.625 ;
        RECT  2.695 0.435 3.115 0.530 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 -0.115 3.360 0.115 ;
        RECT  3.210 -0.115 3.290 0.340 ;
        RECT  0.000 -0.115 3.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.145 3.360 1.375 ;
        RECT  1.040 0.845 1.120 1.375 ;
        RECT  0.700 1.145 1.040 1.375 ;
        RECT  0.620 0.845 0.700 1.375 ;
        RECT  0.310 1.145 0.620 1.375 ;
        RECT  0.230 0.905 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.625 0.775 3.160 0.905 ;
        RECT  2.625 0.205 3.105 0.325 ;
        RECT  0.275 0.205 2.275 0.325 ;
        RECT  3.230 0.885 3.310 1.065 ;
        RECT  2.230 0.995 3.230 1.065 ;
        RECT  2.150 0.640 2.230 1.065 ;
        RECT  1.880 0.995 2.150 1.065 ;
        RECT  1.950 0.705 2.070 0.915 ;
        RECT  1.710 0.705 1.950 0.775 ;
        RECT  1.780 0.845 1.880 1.065 ;
        RECT  1.400 0.995 1.780 1.065 ;
        RECT  1.590 0.705 1.710 0.915 ;
        RECT  1.330 0.705 1.590 0.775 ;
        RECT  1.250 0.705 1.330 1.010 ;
        RECT  0.910 0.705 1.250 0.775 ;
        RECT  0.830 0.705 0.910 1.010 ;
        RECT  0.490 0.705 0.830 0.775 ;
        RECT  0.410 0.705 0.490 1.010 ;
        RECT  0.130 0.705 0.410 0.775 ;
        RECT  0.050 0.705 0.130 1.045 ;
    END
END NR3D3BWP

MACRO NR3D4BWP
    CLASS CORE ;
    FOREIGN NR3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5277 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.875 0.785 3.945 1.040 ;
        RECT  3.255 0.785 3.875 0.905 ;
        RECT  3.255 0.215 3.825 0.335 ;
        RECT  3.045 0.215 3.255 0.905 ;
        RECT  0.435 0.215 3.045 0.335 ;
        RECT  2.790 0.785 3.045 0.905 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.445 1.225 0.625 ;
        RECT  0.285 0.445 1.015 0.515 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.445 2.350 0.625 ;
        RECT  1.430 0.445 2.135 0.515 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.445 3.885 0.625 ;
        RECT  3.340 0.445 3.675 0.525 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.345 ;
        RECT  0.325 -0.115 3.930 0.115 ;
        RECT  0.255 -0.115 0.325 0.345 ;
        RECT  0.000 -0.115 0.255 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 4.060 1.375 ;
        RECT  1.130 0.845 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.845 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.915 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.915 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.875 0.785 3.945 1.040 ;
        RECT  3.325 0.785 3.875 0.905 ;
        RECT  3.325 0.215 3.825 0.335 ;
        RECT  0.435 0.215 2.975 0.335 ;
        RECT  2.790 0.785 2.975 0.905 ;
        RECT  2.690 0.995 3.790 1.065 ;
        RECT  2.695 0.445 2.955 0.530 ;
        RECT  2.610 0.640 2.690 1.065 ;
        RECT  2.300 0.995 2.610 1.065 ;
        RECT  2.370 0.705 2.490 0.915 ;
        RECT  2.130 0.705 2.370 0.775 ;
        RECT  2.200 0.845 2.300 1.065 ;
        RECT  1.940 0.995 2.200 1.065 ;
        RECT  2.010 0.705 2.130 0.915 ;
        RECT  1.770 0.705 2.010 0.775 ;
        RECT  1.840 0.845 1.940 1.065 ;
        RECT  1.460 0.995 1.840 1.065 ;
        RECT  1.650 0.705 1.770 0.915 ;
        RECT  1.390 0.705 1.650 0.775 ;
        RECT  1.310 0.705 1.390 1.010 ;
        RECT  1.030 0.705 1.310 0.775 ;
        RECT  0.950 0.705 1.030 1.010 ;
        RECT  0.670 0.705 0.950 0.775 ;
        RECT  0.590 0.705 0.670 1.010 ;
        RECT  0.310 0.705 0.590 0.775 ;
        RECT  0.230 0.705 0.310 1.010 ;
    END
END NR3D4BWP

MACRO NR3D8BWP
    CLASS CORE ;
    FOREIGN NR3D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.0040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.150 0.720 7.230 1.070 ;
        RECT  5.495 0.720 7.150 0.895 ;
        RECT  5.495 0.225 7.045 0.345 ;
        RECT  5.285 0.225 5.495 0.895 ;
        RECT  0.255 0.225 5.285 0.345 ;
        RECT  4.970 0.720 5.285 0.895 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.3616 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.445 2.345 0.625 ;
        RECT  0.420 0.445 2.135 0.525 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3584 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.445 4.585 0.625 ;
        RECT  2.660 0.445 4.375 0.525 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3616 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.895 0.445 7.105 0.625 ;
        RECT  5.720 0.445 6.895 0.525 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.230 -0.115 7.280 0.115 ;
        RECT  7.150 -0.115 7.230 0.345 ;
        RECT  0.150 -0.115 7.150 0.115 ;
        RECT  0.070 -0.115 0.150 0.320 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.145 7.280 1.375 ;
        RECT  2.240 0.845 2.320 1.375 ;
        RECT  1.930 1.145 2.240 1.375 ;
        RECT  1.850 0.845 1.930 1.375 ;
        RECT  1.570 1.145 1.850 1.375 ;
        RECT  1.490 0.845 1.570 1.375 ;
        RECT  1.210 1.145 1.490 1.375 ;
        RECT  1.130 0.845 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.845 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.845 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.770 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.150 0.720 7.230 1.070 ;
        RECT  5.565 0.720 7.150 0.895 ;
        RECT  5.565 0.225 7.045 0.345 ;
        RECT  0.255 0.225 5.215 0.345 ;
        RECT  4.970 0.720 5.215 0.895 ;
        RECT  4.890 0.985 7.070 1.065 ;
        RECT  4.810 0.700 4.890 1.065 ;
        RECT  4.520 0.985 4.810 1.065 ;
        RECT  4.590 0.705 4.710 0.915 ;
        RECT  4.350 0.705 4.590 0.775 ;
        RECT  4.420 0.845 4.520 1.065 ;
        RECT  4.160 0.985 4.420 1.065 ;
        RECT  4.230 0.705 4.350 0.915 ;
        RECT  3.990 0.705 4.230 0.775 ;
        RECT  4.060 0.845 4.160 1.065 ;
        RECT  3.800 0.985 4.060 1.065 ;
        RECT  3.870 0.705 3.990 0.915 ;
        RECT  3.630 0.705 3.870 0.775 ;
        RECT  3.700 0.845 3.800 1.065 ;
        RECT  3.440 0.985 3.700 1.065 ;
        RECT  3.510 0.705 3.630 0.915 ;
        RECT  3.270 0.705 3.510 0.775 ;
        RECT  3.340 0.845 3.440 1.065 ;
        RECT  3.080 0.985 3.340 1.065 ;
        RECT  3.150 0.705 3.270 0.915 ;
        RECT  2.910 0.705 3.150 0.775 ;
        RECT  2.980 0.845 3.080 1.065 ;
        RECT  2.600 0.985 2.980 1.065 ;
        RECT  2.790 0.705 2.910 0.915 ;
        RECT  2.530 0.705 2.790 0.775 ;
        RECT  2.450 0.705 2.530 1.020 ;
        RECT  2.110 0.705 2.450 0.775 ;
        RECT  2.030 0.705 2.110 1.020 ;
        RECT  1.750 0.705 2.030 0.775 ;
        RECT  1.670 0.705 1.750 1.020 ;
        RECT  1.390 0.705 1.670 0.775 ;
        RECT  1.310 0.705 1.390 1.020 ;
        RECT  1.030 0.705 1.310 0.775 ;
        RECT  0.950 0.705 1.030 1.020 ;
        RECT  0.670 0.705 0.950 0.775 ;
        RECT  0.590 0.705 0.670 1.020 ;
        RECT  0.310 0.705 0.590 0.775 ;
        RECT  0.230 0.705 0.310 1.070 ;
    END
END NR3D8BWP

MACRO NR4D0BWP
    CLASS CORE ;
    FOREIGN NR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0967 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.945 1.075 ;
        RECT  0.725 0.345 0.875 0.415 ;
        RECT  0.840 0.835 0.875 1.075 ;
        RECT  0.655 0.185 0.725 0.415 ;
        RECT  0.305 0.345 0.655 0.415 ;
        RECT  0.235 0.185 0.305 0.415 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.610 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.115 0.980 0.115 ;
        RECT  0.820 -0.115 0.920 0.275 ;
        RECT  0.530 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.145 0.980 1.375 ;
        RECT  0.055 0.695 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
END NR4D0BWP

MACRO NR4D1BWP
    CLASS CORE ;
    FOREIGN NR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1312 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.340 1.440 0.415 ;
        RECT  0.735 0.340 0.805 0.880 ;
        RECT  0.385 0.800 0.735 0.880 ;
        RECT  0.310 0.340 0.385 0.880 ;
        RECT  0.240 0.340 0.310 0.415 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.130 0.495 1.155 0.640 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.530 0.640 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.530 0.235 0.630 ;
        RECT  0.035 0.355 0.105 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 0.520 0.550 0.640 ;
        RECT  0.455 0.355 0.530 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 -0.115 1.680 0.115 ;
        RECT  1.520 -0.115 1.600 0.425 ;
        RECT  1.180 -0.115 1.520 0.115 ;
        RECT  1.100 -0.115 1.180 0.270 ;
        RECT  0.580 -0.115 1.100 0.115 ;
        RECT  0.500 -0.115 0.580 0.270 ;
        RECT  0.170 -0.115 0.500 0.115 ;
        RECT  0.070 -0.115 0.170 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.145 1.680 1.375 ;
        RECT  1.160 0.985 1.240 1.375 ;
        RECT  0.000 1.145 1.160 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.520 0.845 1.600 0.985 ;
        RECT  0.980 0.845 1.520 0.915 ;
        RECT  0.900 0.845 0.980 1.030 ;
        RECT  0.160 0.955 0.900 1.030 ;
        RECT  0.080 0.735 0.160 1.030 ;
    END
END NR4D1BWP

MACRO NR4D2BWP
    CLASS CORE ;
    FOREIGN NR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.855 2.590 0.925 ;
        RECT  2.415 0.215 2.485 0.925 ;
        RECT  0.455 0.215 2.415 0.335 ;
        RECT  2.110 0.855 2.415 0.925 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.445 0.820 0.515 ;
        RECT  0.175 0.355 0.245 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.445 1.390 0.765 ;
        RECT  0.920 0.445 1.295 0.515 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0896 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.445 1.925 0.765 ;
        RECT  1.480 0.445 1.855 0.515 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0904 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.445 2.345 0.765 ;
        RECT  1.995 0.445 2.275 0.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 2.800 1.375 ;
        RECT  0.660 0.845 0.740 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.260 0.880 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.670 0.910 2.750 1.065 ;
        RECT  2.030 0.995 2.670 1.065 ;
        RECT  1.950 0.845 2.030 1.065 ;
        RECT  1.665 0.845 1.950 0.915 ;
        RECT  1.490 0.995 1.870 1.065 ;
        RECT  1.590 0.635 1.665 0.915 ;
        RECT  1.410 0.880 1.490 1.065 ;
        RECT  1.030 0.995 1.410 1.065 ;
        RECT  0.950 0.845 1.330 0.915 ;
        RECT  0.870 0.705 0.950 1.020 ;
        RECT  0.530 0.705 0.870 0.775 ;
        RECT  0.450 0.705 0.530 1.020 ;
        RECT  0.150 0.705 0.450 0.775 ;
        RECT  0.070 0.705 0.150 1.020 ;
    END
END NR4D2BWP

MACRO NR4D3BWP
    CLASS CORE ;
    FOREIGN NR4D3BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4496 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.215 4.145 0.335 ;
        RECT  3.395 0.770 3.990 0.915 ;
        RECT  3.175 0.215 3.395 0.915 ;
        RECT  0.075 0.215 3.175 0.335 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.435 1.085 0.505 ;
        RECT  0.300 0.435 0.525 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.435 1.990 0.505 ;
        RECT  1.295 0.435 1.505 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.435 2.930 0.625 ;
        RECT  2.270 0.435 2.695 0.505 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1356 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.435 4.025 0.625 ;
        RECT  3.535 0.435 3.815 0.505 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.145 4.200 1.375 ;
        RECT  0.980 0.845 1.060 1.375 ;
        RECT  0.670 1.145 0.980 1.375 ;
        RECT  0.590 0.845 0.670 1.375 ;
        RECT  0.310 1.145 0.590 1.375 ;
        RECT  0.230 0.895 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.215 4.145 0.335 ;
        RECT  3.465 0.770 3.990 0.915 ;
        RECT  0.075 0.215 3.115 0.335 ;
        RECT  4.070 0.895 4.150 1.065 ;
        RECT  3.070 0.995 4.070 1.065 ;
        RECT  2.990 0.705 3.070 1.065 ;
        RECT  2.730 0.705 2.990 0.775 ;
        RECT  2.540 0.990 2.910 1.065 ;
        RECT  2.610 0.705 2.730 0.915 ;
        RECT  2.370 0.705 2.610 0.775 ;
        RECT  2.440 0.845 2.540 1.065 ;
        RECT  2.170 0.990 2.440 1.065 ;
        RECT  2.250 0.705 2.370 0.915 ;
        RECT  2.090 0.640 2.170 1.065 ;
        RECT  1.820 0.990 2.090 1.065 ;
        RECT  1.890 0.705 2.010 0.915 ;
        RECT  1.650 0.705 1.890 0.775 ;
        RECT  1.720 0.845 1.820 1.065 ;
        RECT  1.350 0.990 1.720 1.065 ;
        RECT  1.530 0.705 1.650 0.915 ;
        RECT  1.270 0.705 1.530 0.775 ;
        RECT  1.190 0.705 1.270 1.000 ;
        RECT  0.850 0.705 1.190 0.775 ;
        RECT  0.770 0.705 0.850 1.000 ;
        RECT  0.490 0.705 0.770 0.775 ;
        RECT  0.410 0.705 0.490 1.000 ;
        RECT  0.130 0.705 0.410 0.775 ;
        RECT  0.050 0.705 0.130 1.035 ;
    END
END NR4D3BWP

MACRO NR4D4BWP
    CLASS CORE ;
    FOREIGN NR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.6000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.910 0.775 4.990 1.030 ;
        RECT  4.235 0.775 4.910 0.915 ;
        RECT  4.235 0.215 4.745 0.335 ;
        RECT  4.025 0.215 4.235 0.915 ;
        RECT  0.435 0.215 4.025 0.335 ;
        RECT  3.810 0.775 4.025 0.915 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.445 1.225 0.625 ;
        RECT  0.315 0.445 1.015 0.515 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.445 2.485 0.625 ;
        RECT  1.435 0.445 2.275 0.515 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.445 3.580 0.515 ;
        RECT  2.660 0.445 2.905 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1808 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.445 4.865 0.625 ;
        RECT  4.375 0.445 4.655 0.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.925 -0.115 5.040 0.115 ;
        RECT  4.855 -0.115 4.925 0.320 ;
        RECT  0.325 -0.115 4.855 0.115 ;
        RECT  0.255 -0.115 0.325 0.320 ;
        RECT  0.000 -0.115 0.255 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 5.040 1.375 ;
        RECT  1.130 0.845 1.210 1.375 ;
        RECT  0.850 1.145 1.130 1.375 ;
        RECT  0.770 0.845 0.850 1.375 ;
        RECT  0.490 1.145 0.770 1.375 ;
        RECT  0.410 0.845 0.490 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.795 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.910 0.775 4.990 1.030 ;
        RECT  4.305 0.775 4.910 0.915 ;
        RECT  4.305 0.215 4.745 0.335 ;
        RECT  0.435 0.215 3.955 0.335 ;
        RECT  3.810 0.775 3.955 0.915 ;
        RECT  3.725 0.995 4.830 1.065 ;
        RECT  3.655 0.640 3.725 1.065 ;
        RECT  3.380 0.995 3.655 1.065 ;
        RECT  3.450 0.705 3.570 0.915 ;
        RECT  3.210 0.705 3.450 0.775 ;
        RECT  3.280 0.845 3.380 1.065 ;
        RECT  3.020 0.995 3.280 1.065 ;
        RECT  3.090 0.705 3.210 0.915 ;
        RECT  2.850 0.705 3.090 0.775 ;
        RECT  2.920 0.845 3.020 1.065 ;
        RECT  2.650 0.995 2.920 1.065 ;
        RECT  2.730 0.705 2.850 0.915 ;
        RECT  2.310 0.705 2.730 0.775 ;
        RECT  2.570 0.925 2.650 1.065 ;
        RECT  2.390 0.925 2.470 1.065 ;
        RECT  2.120 0.990 2.390 1.065 ;
        RECT  2.190 0.705 2.310 0.915 ;
        RECT  1.950 0.705 2.190 0.775 ;
        RECT  2.020 0.845 2.120 1.065 ;
        RECT  1.760 0.990 2.020 1.065 ;
        RECT  1.830 0.705 1.950 0.915 ;
        RECT  1.590 0.705 1.830 0.775 ;
        RECT  1.660 0.845 1.760 1.065 ;
        RECT  1.390 0.990 1.660 1.065 ;
        RECT  1.470 0.705 1.590 0.915 ;
        RECT  1.310 0.705 1.390 1.065 ;
        RECT  1.030 0.705 1.310 0.775 ;
        RECT  0.950 0.705 1.030 1.020 ;
        RECT  0.670 0.705 0.950 0.775 ;
        RECT  0.590 0.705 0.670 1.020 ;
        RECT  0.310 0.705 0.590 0.775 ;
        RECT  0.230 0.705 0.310 1.075 ;
    END
END NR4D4BWP

MACRO NR4D8BWP
    CLASS CORE ;
    FOREIGN NR4D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.680 2.190 0.800 ;
        RECT  2.095 0.185 2.170 0.465 ;
        RECT  1.805 0.355 2.095 0.465 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.575 0.355 1.735 0.465 ;
        RECT  1.445 0.355 1.575 0.800 ;
        RECT  1.375 0.185 1.445 0.800 ;
        RECT  1.365 0.355 1.375 0.800 ;
        RECT  1.090 0.355 1.365 0.465 ;
        RECT  1.020 0.680 1.365 0.800 ;
        RECT  1.020 0.185 1.090 0.465 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.465 0.805 0.780 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.590 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.465 0.385 0.780 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.940 0.115 ;
        RECT  2.630 -0.115 2.710 0.305 ;
        RECT  2.345 -0.115 2.630 0.115 ;
        RECT  2.275 -0.115 2.345 0.305 ;
        RECT  2.010 -0.115 2.275 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  1.650 -0.115 1.890 0.115 ;
        RECT  1.530 -0.115 1.650 0.275 ;
        RECT  1.290 -0.115 1.530 0.115 ;
        RECT  1.170 -0.115 1.290 0.275 ;
        RECT  0.900 -0.115 1.170 0.115 ;
        RECT  0.780 -0.115 0.900 0.245 ;
        RECT  0.510 -0.115 0.780 0.115 ;
        RECT  0.390 -0.115 0.510 0.245 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.145 2.940 1.375 ;
        RECT  2.610 0.970 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.010 2.370 1.375 ;
        RECT  2.010 1.145 2.250 1.375 ;
        RECT  1.890 1.010 2.010 1.375 ;
        RECT  1.650 1.145 1.890 1.375 ;
        RECT  1.530 1.010 1.650 1.375 ;
        RECT  1.290 1.145 1.530 1.375 ;
        RECT  1.170 1.010 1.290 1.375 ;
        RECT  0.900 1.145 1.170 1.375 ;
        RECT  0.780 1.010 0.900 1.375 ;
        RECT  0.000 1.145 0.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.680 2.190 0.800 ;
        RECT  2.095 0.185 2.170 0.465 ;
        RECT  1.805 0.355 2.095 0.465 ;
        RECT  1.735 0.185 1.805 0.465 ;
        RECT  1.645 0.355 1.735 0.465 ;
        RECT  1.090 0.355 1.295 0.465 ;
        RECT  1.020 0.680 1.295 0.800 ;
        RECT  1.020 0.185 1.090 0.465 ;
        RECT  2.810 0.185 2.890 1.070 ;
        RECT  2.800 0.185 2.810 0.465 ;
        RECT  2.540 0.830 2.810 0.900 ;
        RECT  2.530 0.395 2.800 0.465 ;
        RECT  2.500 0.540 2.730 0.620 ;
        RECT  2.440 0.830 2.540 1.070 ;
        RECT  2.450 0.185 2.530 0.465 ;
        RECT  2.430 0.540 2.500 0.760 ;
        RECT  2.315 0.395 2.450 0.465 ;
        RECT  2.335 0.690 2.430 0.760 ;
        RECT  2.265 0.690 2.335 0.940 ;
        RECT  2.245 0.395 2.315 0.610 ;
        RECT  0.950 0.870 2.265 0.940 ;
        RECT  1.775 0.540 2.245 0.610 ;
        RECT  0.875 0.315 0.950 0.940 ;
        RECT  0.210 0.315 0.875 0.385 ;
        RECT  0.125 0.870 0.875 0.940 ;
        RECT  0.055 0.735 0.125 1.035 ;
    END
END NR4D8BWP

MACRO OA211D0BWP
    CLASS CORE ;
    FOREIGN OA211D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.195 1.085 1.055 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.355 0.755 0.800 ;
        RECT  0.595 0.355 0.685 0.485 ;
        RECT  0.665 0.730 0.685 0.800 ;
        RECT  0.595 0.730 0.665 0.905 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.555 0.600 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.000 -0.115 0.780 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.145 1.120 1.375 ;
        RECT  0.780 1.130 0.900 1.375 ;
        RECT  0.520 1.145 0.780 1.375 ;
        RECT  0.400 1.130 0.520 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 0.930 0.640 ;
        RECT  0.850 0.205 0.920 1.055 ;
        RECT  0.665 0.205 0.850 0.275 ;
        RECT  0.130 0.985 0.850 1.055 ;
        RECT  0.595 0.195 0.665 0.275 ;
        RECT  0.210 0.195 0.595 0.265 ;
        RECT  0.130 0.345 0.520 0.415 ;
        RECT  0.050 0.195 0.130 0.415 ;
        RECT  0.050 0.915 0.130 1.055 ;
    END
END OA211D0BWP

MACRO OA211D1BWP
    CLASS CORE ;
    FOREIGN OA211D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.215 1.085 1.065 ;
        RECT  0.950 0.215 1.015 0.285 ;
        RECT  0.950 0.985 1.015 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.690 0.495 0.735 0.640 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.575 0.640 ;
        RECT  0.455 0.495 0.525 0.905 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.195 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.860 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.860 0.285 ;
        RECT  0.000 -0.115 0.780 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 1.145 1.120 1.375 ;
        RECT  0.790 0.985 0.870 1.375 ;
        RECT  0.520 1.145 0.790 1.375 ;
        RECT  0.400 1.130 0.520 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.915 ;
        RECT  0.210 0.355 0.875 0.425 ;
        RECT  0.685 0.845 0.875 0.915 ;
        RECT  0.615 0.845 0.685 1.055 ;
        RECT  0.130 0.985 0.615 1.055 ;
        RECT  0.145 0.215 0.510 0.285 ;
        RECT  0.035 0.185 0.145 0.285 ;
        RECT  0.050 0.735 0.130 1.055 ;
    END
END OA211D1BWP

MACRO OA211D2BWP
    CLASS CORE ;
    FOREIGN OA211D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.815 ;
        RECT  1.135 0.355 1.155 0.465 ;
        RECT  1.135 0.735 1.155 0.815 ;
        RECT  1.065 0.185 1.135 0.465 ;
        RECT  1.065 0.735 1.135 1.035 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.495 0.665 0.905 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.400 0.115 ;
        RECT  1.240 -0.115 1.320 0.285 ;
        RECT  0.950 -0.115 1.240 0.115 ;
        RECT  0.830 -0.115 0.950 0.275 ;
        RECT  0.000 -0.115 0.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.400 1.375 ;
        RECT  1.240 0.895 1.320 1.375 ;
        RECT  0.950 1.145 1.240 1.375 ;
        RECT  0.830 1.115 0.950 1.375 ;
        RECT  0.550 1.145 0.830 1.375 ;
        RECT  0.430 1.115 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.520 1.020 0.640 ;
        RECT  0.925 0.345 0.995 1.045 ;
        RECT  0.240 0.345 0.925 0.415 ;
        RECT  0.160 0.975 0.925 1.045 ;
        RECT  0.060 0.205 0.540 0.275 ;
        RECT  0.080 0.735 0.160 1.045 ;
    END
END OA211D2BWP

MACRO OA211D4BWP
    CLASS CORE ;
    FOREIGN OA211D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.465 ;
        RECT  2.275 0.695 2.285 1.035 ;
        RECT  2.215 0.185 2.275 1.035 ;
        RECT  2.065 0.355 2.215 0.790 ;
        RECT  1.925 0.355 2.065 0.465 ;
        RECT  1.925 0.695 2.065 0.790 ;
        RECT  1.855 0.185 1.925 0.465 ;
        RECT  1.855 0.695 1.925 1.035 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.765 ;
        RECT  0.245 0.695 0.705 0.765 ;
        RECT  0.165 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.765 ;
        RECT  0.955 0.695 1.435 0.765 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.760 -0.115 2.010 0.115 ;
        RECT  1.660 -0.115 1.760 0.275 ;
        RECT  0.510 -0.115 1.660 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.885 2.130 1.375 ;
        RECT  1.760 1.145 2.010 1.375 ;
        RECT  1.660 0.975 1.760 1.375 ;
        RECT  1.580 1.145 1.660 1.375 ;
        RECT  1.480 0.975 1.580 1.375 ;
        RECT  0.860 1.145 1.480 1.375 ;
        RECT  0.760 0.975 0.860 1.375 ;
        RECT  0.500 1.145 0.760 1.375 ;
        RECT  0.400 0.975 0.500 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.835 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.355 1.995 0.465 ;
        RECT  1.925 0.695 1.995 0.790 ;
        RECT  1.855 0.185 1.925 0.465 ;
        RECT  1.855 0.695 1.925 1.035 ;
        RECT  1.775 0.545 1.970 0.615 ;
        RECT  1.705 0.345 1.775 0.905 ;
        RECT  0.930 0.345 1.705 0.415 ;
        RECT  1.220 0.835 1.705 0.905 ;
        RECT  0.845 0.195 1.590 0.265 ;
        RECT  1.120 0.835 1.220 1.075 ;
        RECT  0.680 0.835 1.120 0.905 ;
        RECT  0.775 0.195 0.845 0.415 ;
        RECT  0.130 0.345 0.775 0.415 ;
        RECT  0.580 0.835 0.680 1.075 ;
        RECT  0.320 0.835 0.580 0.905 ;
        RECT  0.220 0.835 0.320 1.075 ;
        RECT  0.050 0.265 0.130 0.415 ;
    END
END OA211D4BWP

MACRO OA21D0BWP
    CLASS CORE ;
    FOREIGN OA21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0437 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.185 0.945 1.065 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.275 ;
        RECT  0.000 -0.115 0.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 1.125 0.720 1.375 ;
        RECT  0.130 1.145 0.600 1.375 ;
        RECT  0.050 0.925 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.715 0.355 0.785 1.055 ;
        RECT  0.210 0.355 0.715 0.425 ;
        RECT  0.390 0.985 0.715 1.055 ;
        RECT  0.145 0.215 0.530 0.285 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA21D0BWP

MACRO OA21D1BWP
    CLASS CORE ;
    FOREIGN OA21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0874 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.195 0.945 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.275 ;
        RECT  0.000 -0.115 0.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 0.985 0.720 1.375 ;
        RECT  0.140 1.145 0.600 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.715 0.355 0.785 0.915 ;
        RECT  0.210 0.355 0.715 0.425 ;
        RECT  0.525 0.845 0.715 0.915 ;
        RECT  0.145 0.215 0.530 0.285 ;
        RECT  0.455 0.845 0.525 1.055 ;
        RECT  0.390 0.985 0.455 1.055 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA21D1BWP

MACRO OA21D2BWP
    CLASS CORE ;
    FOREIGN OA21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.765 ;
        RECT  0.870 0.355 0.875 0.465 ;
        RECT  0.870 0.675 0.875 0.765 ;
        RECT  0.800 0.185 0.870 0.465 ;
        RECT  0.800 0.675 0.870 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.115 1.120 0.115 ;
        RECT  0.970 -0.115 1.050 0.285 ;
        RECT  0.680 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.680 0.285 ;
        RECT  0.000 -0.115 0.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.145 1.120 1.375 ;
        RECT  0.970 0.955 1.050 1.375 ;
        RECT  0.675 1.145 0.970 1.375 ;
        RECT  0.605 0.975 0.675 1.375 ;
        RECT  0.140 1.145 0.605 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.660 0.355 0.730 0.905 ;
        RECT  0.210 0.355 0.660 0.425 ;
        RECT  0.525 0.835 0.660 0.905 ;
        RECT  0.455 0.835 0.525 1.060 ;
        RECT  0.145 0.215 0.510 0.285 ;
        RECT  0.390 0.985 0.455 1.060 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA21D2BWP

MACRO OA21D4BWP
    CLASS CORE ;
    FOREIGN OA21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 0.185 1.855 1.010 ;
        RECT  1.645 0.355 1.775 0.810 ;
        RECT  1.465 0.355 1.645 0.465 ;
        RECT  1.465 0.695 1.645 0.810 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.695 1.465 1.010 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.115 0.915 ;
        RECT  0.245 0.845 1.015 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.775 ;
        RECT  0.385 0.705 0.855 0.775 ;
        RECT  0.315 0.495 0.385 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 -0.115 2.100 0.115 ;
        RECT  1.950 -0.115 2.030 0.475 ;
        RECT  1.680 -0.115 1.950 0.115 ;
        RECT  1.560 -0.115 1.680 0.275 ;
        RECT  1.280 -0.115 1.560 0.115 ;
        RECT  1.160 -0.115 1.280 0.275 ;
        RECT  0.130 -0.115 1.160 0.115 ;
        RECT  0.050 -0.115 0.130 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.145 2.100 1.375 ;
        RECT  1.950 0.675 2.030 1.375 ;
        RECT  1.680 1.145 1.950 1.375 ;
        RECT  1.560 0.880 1.680 1.375 ;
        RECT  1.280 1.145 1.560 1.375 ;
        RECT  1.160 1.125 1.280 1.375 ;
        RECT  0.700 1.145 1.160 1.375 ;
        RECT  0.580 1.125 0.700 1.375 ;
        RECT  0.120 1.145 0.580 1.375 ;
        RECT  0.050 0.960 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.465 0.355 1.575 0.465 ;
        RECT  1.465 0.695 1.575 0.810 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.695 1.465 1.010 ;
        RECT  1.315 0.545 1.555 0.615 ;
        RECT  1.245 0.345 1.315 1.055 ;
        RECT  0.390 0.345 1.245 0.415 ;
        RECT  0.210 0.985 1.245 1.055 ;
        RECT  0.210 0.205 1.070 0.275 ;
    END
END OA21D4BWP

MACRO OA221D0BWP
    CLASS CORE ;
    FOREIGN OA221D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.345 1.505 1.060 ;
        RECT  1.370 0.345 1.435 0.415 ;
        RECT  1.370 0.985 1.435 1.060 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.120 0.495 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.355 0.525 0.640 ;
        RECT  0.420 0.520 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.280 0.420 ;
        RECT  0.000 -0.115 1.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.145 1.540 1.375 ;
        RECT  1.190 0.985 1.290 1.375 ;
        RECT  0.710 1.145 1.190 1.375 ;
        RECT  0.590 1.115 0.710 1.375 ;
        RECT  0.130 1.145 0.590 1.375 ;
        RECT  0.050 0.945 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.510 1.365 0.915 ;
        RECT  1.110 0.845 1.295 0.915 ;
        RECT  0.610 0.345 1.110 0.415 ;
        RECT  1.040 0.845 1.110 1.045 ;
        RECT  0.340 0.975 1.040 1.045 ;
        RECT  0.130 0.195 0.920 0.275 ;
        RECT  0.270 0.345 0.340 1.045 ;
        RECT  0.220 0.345 0.270 0.415 ;
        RECT  0.050 0.195 0.130 0.315 ;
    END
END OA221D0BWP

MACRO OA221D1BWP
    CLASS CORE ;
    FOREIGN OA221D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 1.075 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.110 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.540 0.780 0.620 ;
        RECT  0.595 0.540 0.685 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.355 0.525 0.640 ;
        RECT  0.400 0.520 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 -0.115 1.540 0.115 ;
        RECT  1.180 -0.115 1.260 0.435 ;
        RECT  0.000 -0.115 1.180 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.160 0.975 1.280 1.375 ;
        RECT  0.690 1.145 1.160 1.375 ;
        RECT  0.570 1.115 0.690 1.375 ;
        RECT  0.140 1.145 0.570 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.265 0.520 1.335 0.905 ;
        RECT  1.085 0.835 1.265 0.905 ;
        RECT  1.015 0.835 1.085 1.045 ;
        RECT  0.960 0.185 1.060 0.425 ;
        RECT  0.490 0.975 1.015 1.045 ;
        RECT  0.700 0.355 0.960 0.425 ;
        RECT  0.130 0.205 0.890 0.275 ;
        RECT  0.600 0.355 0.700 0.455 ;
        RECT  0.410 0.730 0.490 1.045 ;
        RECT  0.330 0.730 0.410 0.800 ;
        RECT  0.260 0.350 0.330 0.800 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA221D1BWP

MACRO OA221D2BWP
    CLASS CORE ;
    FOREIGN OA221D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.765 ;
        RECT  1.425 0.355 1.435 0.470 ;
        RECT  1.430 0.695 1.435 0.765 ;
        RECT  1.360 0.695 1.430 1.045 ;
        RECT  1.355 0.185 1.425 0.470 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.110 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.945 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.755 0.640 ;
        RECT  0.595 0.495 0.665 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.400 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.620 -0.115 1.680 0.115 ;
        RECT  1.520 -0.115 1.620 0.275 ;
        RECT  1.240 -0.115 1.520 0.115 ;
        RECT  1.160 -0.115 1.240 0.435 ;
        RECT  0.000 -0.115 1.160 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.145 1.680 1.375 ;
        RECT  1.530 0.845 1.610 1.375 ;
        RECT  1.240 1.145 1.530 1.375 ;
        RECT  1.160 0.985 1.240 1.375 ;
        RECT  0.690 1.145 1.160 1.375 ;
        RECT  0.570 1.115 0.690 1.375 ;
        RECT  0.140 1.145 0.570 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.220 0.520 1.290 0.905 ;
        RECT  1.085 0.835 1.220 0.905 ;
        RECT  1.015 0.835 1.085 1.045 ;
        RECT  0.960 0.185 1.060 0.425 ;
        RECT  0.330 0.975 1.015 1.045 ;
        RECT  0.590 0.355 0.960 0.425 ;
        RECT  0.140 0.205 0.890 0.275 ;
        RECT  0.260 0.345 0.330 1.045 ;
        RECT  0.230 0.345 0.260 0.445 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END OA221D2BWP

MACRO OA221D4BWP
    CLASS CORE ;
    FOREIGN OA221D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.705 0.465 ;
        RECT  2.695 0.695 2.705 1.035 ;
        RECT  2.635 0.185 2.695 1.035 ;
        RECT  2.485 0.355 2.635 0.815 ;
        RECT  2.345 0.355 2.485 0.465 ;
        RECT  2.345 0.695 2.485 0.815 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.695 2.345 1.035 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.945 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.495 1.365 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.525 0.775 ;
        RECT  1.020 0.705 1.435 0.775 ;
        RECT  0.950 0.520 1.020 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.730 0.640 ;
        RECT  0.595 0.495 0.665 0.905 ;
        RECT  0.245 0.835 0.595 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.475 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.280 ;
        RECT  2.170 -0.115 2.430 0.115 ;
        RECT  2.090 -0.115 2.170 0.435 ;
        RECT  1.820 -0.115 2.090 0.115 ;
        RECT  1.720 -0.115 1.820 0.275 ;
        RECT  0.000 -0.115 1.720 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.675 2.890 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 0.885 2.550 1.375 ;
        RECT  2.190 1.145 2.430 1.375 ;
        RECT  2.070 0.985 2.190 1.375 ;
        RECT  1.820 1.145 2.070 1.375 ;
        RECT  1.720 0.985 1.820 1.375 ;
        RECT  1.640 1.145 1.720 1.375 ;
        RECT  1.540 0.985 1.640 1.375 ;
        RECT  0.900 1.145 1.540 1.375 ;
        RECT  0.780 1.115 0.900 1.375 ;
        RECT  0.145 1.145 0.780 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.465 ;
        RECT  2.345 0.695 2.415 0.815 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.695 2.345 1.035 ;
        RECT  2.200 0.545 2.320 0.615 ;
        RECT  2.130 0.545 2.200 0.915 ;
        RECT  1.990 0.845 2.130 0.915 ;
        RECT  1.900 0.185 2.000 0.425 ;
        RECT  1.910 0.845 1.990 1.075 ;
        RECT  1.270 0.845 1.910 0.915 ;
        RECT  0.990 0.355 1.900 0.425 ;
        RECT  0.130 0.205 1.650 0.275 ;
        RECT  1.190 0.845 1.270 1.045 ;
        RECT  0.870 0.975 1.190 1.045 ;
        RECT  0.800 0.345 0.870 1.045 ;
        RECT  0.210 0.345 0.800 0.415 ;
        RECT  0.390 0.975 0.800 1.045 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA221D4BWP

MACRO OA222D0BWP
    CLASS CORE ;
    FOREIGN OA222D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.045 ;
        RECT  1.535 0.185 1.575 0.285 ;
        RECT  1.540 0.940 1.575 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.635 1.085 0.905 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.640 ;
        RECT  1.260 0.520 1.295 0.640 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.635 0.665 0.905 ;
        RECT  0.545 0.635 0.595 0.780 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.435 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.450 -0.115 1.680 0.115 ;
        RECT  1.370 -0.115 1.450 0.270 ;
        RECT  1.085 -0.115 1.370 0.115 ;
        RECT  1.015 -0.115 1.085 0.270 ;
        RECT  0.000 -0.115 1.015 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.145 1.680 1.375 ;
        RECT  1.360 0.920 1.440 1.375 ;
        RECT  0.910 1.145 1.360 1.375 ;
        RECT  0.790 1.115 0.910 1.375 ;
        RECT  0.170 1.145 0.790 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.435 0.675 1.505 0.840 ;
        RECT  1.285 0.770 1.435 0.840 ;
        RECT  1.225 0.185 1.290 0.255 ;
        RECT  1.215 0.770 1.285 1.045 ;
        RECT  1.155 0.185 1.225 0.420 ;
        RECT  0.320 0.975 1.215 1.045 ;
        RECT  0.610 0.350 1.155 0.420 ;
        RECT  0.050 0.195 0.930 0.265 ;
        RECT  0.105 0.345 0.370 0.415 ;
        RECT  0.250 0.890 0.320 1.045 ;
        RECT  0.105 0.890 0.250 0.960 ;
        RECT  0.035 0.345 0.105 0.960 ;
    END
END OA222D0BWP

MACRO OA222D1BWP
    CLASS CORE ;
    FOREIGN OA222D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.195 1.645 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.495 1.085 0.905 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.540 1.340 0.625 ;
        RECT  1.155 0.355 1.225 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.905 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.435 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 -0.115 1.680 0.115 ;
        RECT  1.360 -0.115 1.440 0.440 ;
        RECT  1.070 -0.115 1.360 0.115 ;
        RECT  0.950 -0.115 1.070 0.145 ;
        RECT  0.000 -0.115 0.950 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 0.985 1.460 1.375 ;
        RECT  0.910 1.145 1.340 1.375 ;
        RECT  0.790 1.115 0.910 1.375 ;
        RECT  0.170 1.145 0.790 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.420 0.520 1.490 0.915 ;
        RECT  1.235 0.845 1.420 0.915 ;
        RECT  0.590 0.215 1.270 0.285 ;
        RECT  1.165 0.845 1.235 1.045 ;
        RECT  0.385 0.975 1.165 1.045 ;
        RECT  0.510 0.355 0.890 0.425 ;
        RECT  0.430 0.195 0.510 0.425 ;
        RECT  0.050 0.195 0.430 0.265 ;
        RECT  0.315 0.890 0.385 1.045 ;
        RECT  0.105 0.345 0.350 0.415 ;
        RECT  0.105 0.890 0.315 0.960 ;
        RECT  0.035 0.345 0.105 0.960 ;
    END
END OA222D1BWP

MACRO OA222D2BWP
    CLASS CORE ;
    FOREIGN OA222D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.355 1.645 0.780 ;
        RECT  1.575 0.185 1.590 1.045 ;
        RECT  1.520 0.185 1.575 0.465 ;
        RECT  1.520 0.710 1.575 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.290 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.810 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 -0.115 1.820 0.115 ;
        RECT  1.675 -0.115 1.785 0.280 ;
        RECT  1.410 -0.115 1.675 0.115 ;
        RECT  1.330 -0.115 1.410 0.435 ;
        RECT  1.060 -0.115 1.330 0.115 ;
        RECT  0.960 -0.115 1.060 0.275 ;
        RECT  0.000 -0.115 0.960 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.860 1.770 1.375 ;
        RECT  1.430 1.145 1.690 1.375 ;
        RECT  1.310 1.030 1.430 1.375 ;
        RECT  0.890 1.145 1.310 1.375 ;
        RECT  0.770 1.030 0.890 1.375 ;
        RECT  0.170 1.145 0.770 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.440 0.545 1.500 0.615 ;
        RECT  1.370 0.545 1.440 0.960 ;
        RECT  0.105 0.890 1.370 0.960 ;
        RECT  1.130 0.205 1.250 0.415 ;
        RECT  0.590 0.345 1.130 0.415 ;
        RECT  0.510 0.195 0.890 0.265 ;
        RECT  0.430 0.195 0.510 0.425 ;
        RECT  0.050 0.195 0.430 0.265 ;
        RECT  0.105 0.345 0.350 0.415 ;
        RECT  0.035 0.345 0.105 0.960 ;
    END
END OA222D2BWP

MACRO OA222D4BWP
    CLASS CORE ;
    FOREIGN OA222D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.695 3.125 1.035 ;
        RECT  3.055 0.185 3.115 1.035 ;
        RECT  2.905 0.355 3.055 0.815 ;
        RECT  2.765 0.355 2.905 0.465 ;
        RECT  2.765 0.695 2.905 0.815 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.695 2.765 1.035 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.215 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.495 2.485 0.905 ;
        RECT  2.055 0.835 2.385 0.905 ;
        RECT  1.985 0.545 2.055 0.905 ;
        RECT  1.820 0.545 1.985 0.615 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.515 0.765 ;
        RECT  1.415 0.695 1.435 0.765 ;
        RECT  1.345 0.695 1.415 0.905 ;
        RECT  1.085 0.835 1.345 0.905 ;
        RECT  1.015 0.495 1.085 0.905 ;
        RECT  0.950 0.495 1.015 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.730 0.640 ;
        RECT  0.595 0.495 0.665 0.905 ;
        RECT  0.245 0.835 0.595 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.475 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.280 ;
        RECT  2.580 -0.115 2.850 0.115 ;
        RECT  2.500 -0.115 2.580 0.425 ;
        RECT  2.210 -0.115 2.500 0.115 ;
        RECT  2.130 -0.115 2.210 0.285 ;
        RECT  0.000 -0.115 2.130 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.675 3.310 1.375 ;
        RECT  2.970 1.145 3.230 1.375 ;
        RECT  2.850 0.885 2.970 1.375 ;
        RECT  2.600 1.145 2.850 1.375 ;
        RECT  2.480 1.115 2.600 1.375 ;
        RECT  1.665 1.145 2.480 1.375 ;
        RECT  1.545 1.115 1.665 1.375 ;
        RECT  0.900 1.145 1.545 1.375 ;
        RECT  0.780 1.115 0.900 1.375 ;
        RECT  0.145 1.145 0.780 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.355 2.835 0.465 ;
        RECT  2.765 0.695 2.835 0.815 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.695 0.695 2.765 1.035 ;
        RECT  2.625 0.545 2.740 0.615 ;
        RECT  2.555 0.545 2.625 1.045 ;
        RECT  0.870 0.975 2.555 1.045 ;
        RECT  2.290 0.215 2.410 0.425 ;
        RECT  2.025 0.355 2.290 0.425 ;
        RECT  1.955 0.190 2.025 0.425 ;
        RECT  0.990 0.355 1.955 0.425 ;
        RECT  1.520 0.835 1.880 0.905 ;
        RECT  0.130 0.205 1.650 0.275 ;
        RECT  0.800 0.345 0.870 1.045 ;
        RECT  0.210 0.345 0.800 0.415 ;
        RECT  0.390 0.975 0.800 1.045 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA222D4BWP

MACRO OA22D0BWP
    CLASS CORE ;
    FOREIGN OA22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0468 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.195 1.365 1.060 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.635 0.825 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.140 -0.115 1.400 0.115 ;
        RECT  1.020 -0.115 1.140 0.285 ;
        RECT  0.340 -0.115 1.020 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.165 1.145 1.400 1.375 ;
        RECT  1.045 1.115 1.165 1.375 ;
        RECT  0.915 1.145 1.045 1.375 ;
        RECT  0.795 1.115 0.915 1.375 ;
        RECT  0.130 1.145 0.795 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.130 0.355 1.200 1.045 ;
        RECT  0.600 0.355 1.130 0.425 ;
        RECT  0.410 0.975 1.130 1.045 ;
        RECT  0.140 0.215 0.930 0.285 ;
        RECT  0.040 0.215 0.140 0.315 ;
    END
END OA22D0BWP

MACRO OA22D1BWP
    CLASS CORE ;
    FOREIGN OA22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.185 1.225 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 -0.115 1.260 0.115 ;
        RECT  0.940 -0.115 1.040 0.275 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.145 1.260 1.375 ;
        RECT  0.950 0.980 1.030 1.375 ;
        RECT  0.850 1.145 0.950 1.375 ;
        RECT  0.770 0.980 0.850 1.375 ;
        RECT  0.140 1.145 0.770 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.345 1.065 0.905 ;
        RECT  0.570 0.345 0.995 0.415 ;
        RECT  0.675 0.835 0.995 0.905 ;
        RECT  0.490 0.195 0.870 0.265 ;
        RECT  0.605 0.835 0.675 1.045 ;
        RECT  0.390 0.975 0.605 1.045 ;
        RECT  0.410 0.195 0.490 0.415 ;
        RECT  0.130 0.345 0.410 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OA22D1BWP

MACRO OA22D2BWP
    CLASS CORE ;
    FOREIGN OA22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.185 1.245 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.575 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 -0.115 1.540 0.115 ;
        RECT  1.355 -0.115 1.425 0.475 ;
        RECT  1.070 -0.115 1.355 0.115 ;
        RECT  0.990 -0.115 1.070 0.275 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.135 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 1.145 1.540 1.375 ;
        RECT  1.355 0.675 1.425 1.375 ;
        RECT  1.070 1.145 1.355 1.375 ;
        RECT  0.990 0.980 1.070 1.375 ;
        RECT  0.890 1.145 0.990 1.375 ;
        RECT  0.810 0.980 0.890 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.010 0.355 1.085 0.905 ;
        RECT  0.605 0.355 1.010 0.425 ;
        RECT  0.730 0.835 1.010 0.905 ;
        RECT  0.130 0.205 0.920 0.275 ;
        RECT  0.660 0.835 0.730 1.045 ;
        RECT  0.410 0.975 0.660 1.045 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA22D2BWP

MACRO OA22D4BWP
    CLASS CORE ;
    FOREIGN OA22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.185 2.285 0.465 ;
        RECT  2.275 0.770 2.285 1.050 ;
        RECT  2.215 0.185 2.275 1.050 ;
        RECT  2.065 0.355 2.215 0.905 ;
        RECT  1.925 0.355 2.065 0.465 ;
        RECT  1.925 0.770 2.065 0.905 ;
        RECT  1.855 0.185 1.925 0.465 ;
        RECT  1.855 0.770 1.925 1.050 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.775 ;
        RECT  0.525 0.705 0.665 0.775 ;
        RECT  0.455 0.705 0.525 0.915 ;
        RECT  0.105 0.845 0.455 0.915 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.915 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.420 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.775 ;
        RECT  0.945 0.705 1.435 0.775 ;
        RECT  0.875 0.495 0.945 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.225 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.465 ;
        RECT  2.130 -0.115 2.390 0.115 ;
        RECT  2.010 -0.115 2.130 0.280 ;
        RECT  1.760 -0.115 2.010 0.115 ;
        RECT  1.660 -0.115 1.760 0.275 ;
        RECT  0.670 -0.115 1.660 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.310 -0.115 0.590 0.115 ;
        RECT  0.230 -0.115 0.310 0.275 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.675 2.470 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.980 2.130 1.375 ;
        RECT  1.760 1.145 2.010 1.375 ;
        RECT  1.660 0.985 1.760 1.375 ;
        RECT  1.580 1.145 1.660 1.375 ;
        RECT  1.480 0.985 1.580 1.375 ;
        RECT  0.870 1.145 1.480 1.375 ;
        RECT  0.750 0.990 0.870 1.375 ;
        RECT  0.140 1.145 0.750 1.375 ;
        RECT  0.040 0.985 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.355 1.995 0.465 ;
        RECT  1.925 0.770 1.995 0.905 ;
        RECT  1.855 0.185 1.925 0.465 ;
        RECT  1.855 0.770 1.925 1.050 ;
        RECT  1.775 0.545 1.970 0.615 ;
        RECT  1.705 0.345 1.775 0.915 ;
        RECT  0.930 0.345 1.705 0.415 ;
        RECT  1.210 0.845 1.705 0.915 ;
        RECT  0.845 0.195 1.590 0.265 ;
        RECT  1.130 0.845 1.210 1.075 ;
        RECT  0.680 0.845 1.130 0.915 ;
        RECT  0.775 0.195 0.845 0.415 ;
        RECT  0.500 0.345 0.775 0.415 ;
        RECT  0.610 0.845 0.680 1.055 ;
        RECT  0.390 0.985 0.610 1.055 ;
        RECT  0.400 0.190 0.500 0.415 ;
        RECT  0.130 0.345 0.400 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OA22D4BWP

MACRO OA31D0BWP
    CLASS CORE ;
    FOREIGN OA31D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0437 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.085 1.060 ;
        RECT  0.995 0.185 1.015 0.305 ;
        RECT  0.995 0.925 1.015 1.060 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.520 0.755 0.705 ;
        RECT  0.665 0.635 0.685 0.705 ;
        RECT  0.595 0.635 0.665 0.905 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.580 0.565 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.735 0.385 1.045 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.890 -0.115 1.120 0.115 ;
        RECT  0.790 -0.115 0.890 0.265 ;
        RECT  0.000 -0.115 0.790 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 1.115 0.880 1.375 ;
        RECT  0.130 1.145 0.760 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.925 0.520 0.945 0.640 ;
        RECT  0.855 0.335 0.925 1.045 ;
        RECT  0.130 0.335 0.855 0.405 ;
        RECT  0.570 0.975 0.855 1.045 ;
        RECT  0.210 0.195 0.710 0.265 ;
        RECT  0.050 0.185 0.130 0.405 ;
    END
END OA31D0BWP

MACRO OA31D1BWP
    CLASS CORE ;
    FOREIGN OA31D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.195 1.085 1.070 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.905 ;
        RECT  0.595 0.775 0.665 0.905 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.560 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 1.120 0.115 ;
        RECT  0.760 -0.115 0.880 0.145 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 1.115 0.880 1.375 ;
        RECT  0.140 1.145 0.760 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.855 0.215 0.925 1.045 ;
        RECT  0.145 0.215 0.855 0.285 ;
        RECT  0.570 0.975 0.855 1.045 ;
        RECT  0.210 0.355 0.690 0.425 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA31D1BWP

MACRO OA31D2BWP
    CLASS CORE ;
    FOREIGN OA31D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.775 ;
        RECT  1.145 0.355 1.155 0.465 ;
        RECT  1.145 0.705 1.155 0.775 ;
        RECT  1.075 0.195 1.145 0.465 ;
        RECT  1.075 0.705 1.145 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.905 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.245 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.115 1.400 0.115 ;
        RECT  1.250 -0.115 1.330 0.285 ;
        RECT  0.960 -0.115 1.250 0.115 ;
        RECT  0.840 -0.115 0.960 0.145 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.145 1.400 1.375 ;
        RECT  1.240 0.845 1.340 1.375 ;
        RECT  0.960 1.145 1.240 1.375 ;
        RECT  0.840 1.115 0.960 1.375 ;
        RECT  0.185 1.145 0.840 1.375 ;
        RECT  0.115 0.705 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.935 0.215 1.005 1.045 ;
        RECT  0.200 0.215 0.935 0.285 ;
        RECT  0.630 0.975 0.935 1.045 ;
        RECT  0.270 0.355 0.750 0.425 ;
        RECT  0.100 0.185 0.200 0.285 ;
    END
END OA31D2BWP

MACRO OA31D4BWP
    CLASS CORE ;
    FOREIGN OA31D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.335 0.185 2.415 1.035 ;
        RECT  2.205 0.355 2.335 0.815 ;
        RECT  2.045 0.355 2.205 0.465 ;
        RECT  2.045 0.695 2.205 0.815 ;
        RECT  1.975 0.185 2.045 0.465 ;
        RECT  1.975 0.695 2.045 1.035 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.355 1.505 0.640 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.810 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.905 0.520 0.975 0.775 ;
        RECT  0.405 0.705 0.905 0.775 ;
        RECT  0.315 0.495 0.405 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 0.520 1.150 0.915 ;
        RECT  0.245 0.845 1.080 0.915 ;
        RECT  0.145 0.495 0.245 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.480 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.280 ;
        RECT  1.870 -0.115 2.130 0.115 ;
        RECT  1.790 -0.115 1.870 0.465 ;
        RECT  1.500 -0.115 1.790 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  0.000 -0.115 1.380 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.675 2.590 1.375 ;
        RECT  2.250 1.145 2.510 1.375 ;
        RECT  2.130 0.885 2.250 1.375 ;
        RECT  1.870 1.145 2.130 1.375 ;
        RECT  1.790 0.685 1.870 1.375 ;
        RECT  1.650 1.145 1.790 1.375 ;
        RECT  1.570 0.850 1.650 1.375 ;
        RECT  1.300 1.145 1.570 1.375 ;
        RECT  1.180 1.125 1.300 1.375 ;
        RECT  0.160 1.145 1.180 1.375 ;
        RECT  0.060 0.985 0.160 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.045 0.355 2.135 0.465 ;
        RECT  2.045 0.695 2.135 0.815 ;
        RECT  1.975 0.185 2.045 0.465 ;
        RECT  1.975 0.695 2.045 1.035 ;
        RECT  1.680 0.545 2.125 0.615 ;
        RECT  1.610 0.210 1.690 0.470 ;
        RECT  1.610 0.545 1.680 0.780 ;
        RECT  0.150 0.210 1.610 0.280 ;
        RECT  1.490 0.710 1.610 0.780 ;
        RECT  1.370 0.710 1.490 1.070 ;
        RECT  1.290 0.710 1.370 0.780 ;
        RECT  1.220 0.350 1.290 1.055 ;
        RECT  0.230 0.350 1.220 0.420 ;
        RECT  0.630 0.985 1.220 1.055 ;
        RECT  0.070 0.210 0.150 0.385 ;
    END
END OA31D4BWP

MACRO OA32D0BWP
    CLASS CORE ;
    FOREIGN OA32D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 1.055 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.635 0.810 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.610 0.835 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.195 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.540 0.115 ;
        RECT  1.190 -0.115 1.310 0.145 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.800 -0.115 0.920 0.145 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.540 1.375 ;
        RECT  1.210 0.990 1.330 1.375 ;
        RECT  0.130 1.145 1.210 1.375 ;
        RECT  0.050 0.915 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.215 1.345 0.915 ;
        RECT  0.145 0.215 1.275 0.285 ;
        RECT  0.950 0.845 1.275 0.915 ;
        RECT  0.220 0.355 1.130 0.425 ;
        RECT  0.880 0.845 0.950 1.055 ;
        RECT  0.610 0.985 0.880 1.055 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA32D0BWP

MACRO OA32D1BWP
    CLASS CORE ;
    FOREIGN OA32D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.585 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.540 0.115 ;
        RECT  1.190 -0.115 1.310 0.140 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.800 -0.115 0.920 0.140 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.540 1.375 ;
        RECT  1.210 0.990 1.330 1.375 ;
        RECT  1.085 1.145 1.210 1.375 ;
        RECT  1.015 0.995 1.085 1.375 ;
        RECT  0.140 1.145 1.015 1.375 ;
        RECT  0.040 0.705 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.215 1.345 0.915 ;
        RECT  0.145 0.215 1.275 0.285 ;
        RECT  0.945 0.845 1.275 0.915 ;
        RECT  0.220 0.355 1.110 0.425 ;
        RECT  0.875 0.845 0.945 1.045 ;
        RECT  0.610 0.975 0.875 1.045 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA32D1BWP

MACRO OA32D2BWP
    CLASS CORE ;
    FOREIGN OA32D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.355 1.505 0.765 ;
        RECT  1.435 0.195 1.445 1.045 ;
        RECT  1.375 0.195 1.435 0.465 ;
        RECT  1.375 0.695 1.435 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.540 1.010 0.615 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 -0.115 1.680 0.115 ;
        RECT  1.535 -0.115 1.645 0.285 ;
        RECT  1.270 -0.115 1.535 0.115 ;
        RECT  1.150 -0.115 1.270 0.140 ;
        RECT  0.880 -0.115 1.150 0.115 ;
        RECT  0.760 -0.115 0.880 0.140 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.835 1.630 1.375 ;
        RECT  1.280 1.145 1.550 1.375 ;
        RECT  1.180 0.985 1.280 1.375 ;
        RECT  0.140 1.145 1.180 1.375 ;
        RECT  0.040 0.705 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.235 0.215 1.305 0.915 ;
        RECT  0.145 0.215 1.235 0.285 ;
        RECT  1.005 0.845 1.235 0.915 ;
        RECT  0.210 0.355 1.070 0.425 ;
        RECT  0.935 0.845 1.005 1.045 ;
        RECT  0.570 0.975 0.935 1.045 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA32D2BWP

MACRO OA32D4BWP
    CLASS CORE ;
    FOREIGN OA32D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.705 0.465 ;
        RECT  2.695 0.695 2.705 1.035 ;
        RECT  2.635 0.185 2.695 1.035 ;
        RECT  2.485 0.355 2.635 0.815 ;
        RECT  2.345 0.355 2.485 0.465 ;
        RECT  2.345 0.695 2.485 0.815 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.695 2.345 1.035 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.645 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.495 1.925 0.765 ;
        RECT  1.785 0.690 1.830 0.765 ;
        RECT  1.715 0.690 1.785 0.905 ;
        RECT  1.365 0.835 1.715 0.905 ;
        RECT  1.265 0.495 1.365 0.905 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.775 ;
        RECT  0.410 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.410 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.120 0.915 ;
        RECT  0.245 0.845 1.015 0.915 ;
        RECT  0.155 0.495 0.245 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.475 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.280 ;
        RECT  2.180 -0.115 2.430 0.115 ;
        RECT  2.080 -0.115 2.180 0.275 ;
        RECT  1.800 -0.115 2.080 0.115 ;
        RECT  1.680 -0.115 1.800 0.135 ;
        RECT  1.420 -0.115 1.680 0.115 ;
        RECT  1.300 -0.115 1.420 0.135 ;
        RECT  0.000 -0.115 1.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.675 2.890 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 0.885 2.550 1.375 ;
        RECT  2.150 1.145 2.430 1.375 ;
        RECT  2.070 0.975 2.150 1.375 ;
        RECT  1.980 1.145 2.070 1.375 ;
        RECT  1.860 1.125 1.980 1.375 ;
        RECT  1.240 1.145 1.860 1.375 ;
        RECT  1.120 1.125 1.240 1.375 ;
        RECT  0.145 1.145 1.120 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.465 ;
        RECT  2.345 0.695 2.415 0.815 ;
        RECT  2.275 0.185 2.345 0.465 ;
        RECT  2.275 0.695 2.345 1.035 ;
        RECT  2.195 0.540 2.320 0.620 ;
        RECT  2.125 0.345 2.195 0.905 ;
        RECT  0.210 0.345 2.125 0.415 ;
        RECT  1.945 0.835 2.125 0.905 ;
        RECT  0.130 0.205 1.990 0.275 ;
        RECT  1.875 0.835 1.945 1.055 ;
        RECT  0.570 0.985 1.875 1.055 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA32D4BWP

MACRO OA33D0BWP
    CLASS CORE ;
    FOREIGN OA33D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.190 1.505 1.070 ;
        RECT  1.400 0.190 1.435 0.290 ;
        RECT  1.400 0.970 1.435 1.070 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.495 0.805 0.765 ;
        RECT  0.685 0.495 0.730 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.965 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.225 0.765 ;
        RECT  1.110 0.495 1.135 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.760 0.610 0.830 ;
        RECT  0.455 0.760 0.525 1.045 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.320 0.140 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.140 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.540 1.375 ;
        RECT  1.200 1.120 1.320 1.375 ;
        RECT  0.130 1.145 1.200 1.375 ;
        RECT  0.050 0.925 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.355 1.365 0.905 ;
        RECT  1.295 0.355 1.330 1.050 ;
        RECT  1.275 0.355 1.295 0.425 ;
        RECT  1.255 0.835 1.295 1.050 ;
        RECT  1.200 0.215 1.275 0.425 ;
        RECT  0.610 0.980 1.255 1.050 ;
        RECT  0.145 0.215 1.200 0.285 ;
        RECT  0.220 0.355 1.120 0.425 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OA33D0BWP

MACRO OA33D1BWP
    CLASS CORE ;
    FOREIGN OA33D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.495 0.805 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.130 0.640 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.905 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.540 0.115 ;
        RECT  1.180 -0.115 1.300 0.135 ;
        RECT  0.880 -0.115 1.180 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 1.125 1.300 1.375 ;
        RECT  0.140 1.145 1.180 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.205 1.345 1.055 ;
        RECT  0.140 0.205 1.275 0.275 ;
        RECT  0.570 0.985 1.275 1.055 ;
        RECT  0.210 0.345 1.080 0.415 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END OA33D1BWP

MACRO OA33D2BWP
    CLASS CORE ;
    FOREIGN OA33D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.355 1.505 0.765 ;
        RECT  1.435 0.195 1.450 1.045 ;
        RECT  1.380 0.195 1.435 0.470 ;
        RECT  1.380 0.695 1.435 1.045 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.640 0.545 0.735 0.615 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.130 0.640 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.905 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.520 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 -0.115 1.680 0.115 ;
        RECT  1.535 -0.115 1.645 0.285 ;
        RECT  1.280 -0.115 1.535 0.115 ;
        RECT  1.160 -0.115 1.280 0.135 ;
        RECT  0.880 -0.115 1.160 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.145 1.680 1.375 ;
        RECT  1.540 0.850 1.640 1.375 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.160 1.125 1.280 1.375 ;
        RECT  0.140 1.145 1.160 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.240 0.205 1.310 1.055 ;
        RECT  0.140 0.205 1.240 0.275 ;
        RECT  0.570 0.985 1.240 1.055 ;
        RECT  0.210 0.345 1.080 0.415 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END OA33D2BWP

MACRO OA33D4BWP
    CLASS CORE ;
    FOREIGN OA33D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.125 0.465 ;
        RECT  3.115 0.695 3.125 1.045 ;
        RECT  3.055 0.185 3.115 1.045 ;
        RECT  2.905 0.350 3.055 0.815 ;
        RECT  2.765 0.350 2.905 0.465 ;
        RECT  2.745 0.695 2.905 0.815 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.675 0.695 2.745 1.045 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.095 0.655 ;
        RECT  1.995 0.495 2.065 0.775 ;
        RECT  1.530 0.705 1.995 0.775 ;
        RECT  1.435 0.495 1.530 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.495 2.345 0.785 ;
        RECT  2.205 0.715 2.270 0.785 ;
        RECT  2.135 0.715 2.205 0.915 ;
        RECT  1.365 0.845 2.135 0.915 ;
        RECT  1.285 0.495 1.365 0.915 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.670 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.775 ;
        RECT  0.385 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.385 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 0.520 1.140 0.915 ;
        RECT  0.245 0.845 1.060 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.130 0.495 0.175 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.475 ;
        RECT  2.970 -0.115 3.230 0.115 ;
        RECT  2.850 -0.115 2.970 0.280 ;
        RECT  2.590 -0.115 2.850 0.115 ;
        RECT  2.510 -0.115 2.590 0.275 ;
        RECT  2.240 -0.115 2.510 0.115 ;
        RECT  2.120 -0.115 2.240 0.135 ;
        RECT  1.860 -0.115 2.120 0.115 ;
        RECT  1.740 -0.115 1.860 0.135 ;
        RECT  1.480 -0.115 1.740 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  0.000 -0.115 1.360 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.675 3.310 1.375 ;
        RECT  2.960 1.145 3.230 1.375 ;
        RECT  2.840 0.885 2.960 1.375 ;
        RECT  2.585 1.145 2.840 1.375 ;
        RECT  2.475 0.995 2.585 1.375 ;
        RECT  2.380 1.145 2.475 1.375 ;
        RECT  2.260 1.125 2.380 1.375 ;
        RECT  1.280 1.145 2.260 1.375 ;
        RECT  1.160 1.125 1.280 1.375 ;
        RECT  0.145 1.145 1.160 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.350 2.835 0.465 ;
        RECT  2.745 0.695 2.835 0.815 ;
        RECT  2.695 0.185 2.765 0.465 ;
        RECT  2.675 0.695 2.745 1.045 ;
        RECT  2.605 0.545 2.805 0.615 ;
        RECT  2.535 0.345 2.605 0.925 ;
        RECT  0.220 0.345 2.535 0.415 ;
        RECT  2.345 0.855 2.535 0.925 ;
        RECT  0.130 0.205 2.430 0.275 ;
        RECT  2.275 0.855 2.345 1.055 ;
        RECT  0.610 0.985 2.275 1.055 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA33D4BWP

MACRO OAI211D0BWP
    CLASS CORE ;
    FOREIGN OAI211D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0844 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.915 0.745 1.045 ;
        RECT  0.525 0.975 0.675 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.125 0.975 0.455 1.045 ;
        RECT  0.055 0.915 0.125 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.760 0.545 0.875 0.615 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.310 ;
        RECT  0.000 -0.115 0.850 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.920 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 1.115 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.205 0.530 0.275 ;
        RECT  0.050 0.205 0.130 0.335 ;
    END
END OAI211D0BWP

MACRO OAI211D1BWP
    CLASS CORE ;
    FOREIGN OAI211D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1521 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.765 0.745 1.045 ;
        RECT  0.525 0.975 0.675 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.125 0.975 0.455 1.045 ;
        RECT  0.055 0.915 0.125 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.760 0.545 0.875 0.615 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.940 0.415 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.840 0.845 0.940 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.115 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.205 0.530 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OAI211D1BWP

MACRO OAI211D2BWP
    CLASS CORE ;
    FOREIGN OAI211D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 1.470 0.415 ;
        RECT  0.945 0.985 1.290 1.055 ;
        RECT  0.875 0.715 0.945 1.055 ;
        RECT  0.805 0.345 0.875 0.785 ;
        RECT  0.670 0.985 0.875 1.055 ;
        RECT  0.590 0.835 0.670 1.055 ;
        RECT  0.320 0.835 0.590 0.905 ;
        RECT  0.220 0.835 0.320 1.075 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.735 0.640 ;
        RECT  0.595 0.520 0.665 0.765 ;
        RECT  0.245 0.695 0.595 0.765 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.525 0.905 ;
        RECT  1.085 0.835 1.435 0.905 ;
        RECT  1.015 0.520 1.085 0.905 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 1.680 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.145 1.680 1.375 ;
        RECT  1.535 0.985 1.645 1.375 ;
        RECT  0.900 1.145 1.535 1.375 ;
        RECT  0.780 1.125 0.900 1.375 ;
        RECT  0.500 1.145 0.780 1.375 ;
        RECT  0.400 0.985 0.500 1.375 ;
        RECT  0.140 1.145 0.400 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.550 0.205 1.630 0.395 ;
        RECT  0.670 0.205 1.550 0.275 ;
        RECT  0.600 0.205 0.670 0.415 ;
        RECT  0.130 0.345 0.600 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OAI211D2BWP

MACRO OAI211D4BWP
    CLASS CORE ;
    FOREIGN OAI211D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5674 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.040 0.705 3.120 1.035 ;
        RECT  2.720 0.705 3.040 0.820 ;
        RECT  2.640 0.705 2.720 1.035 ;
        RECT  2.320 0.705 2.640 0.820 ;
        RECT  2.240 0.705 2.320 1.035 ;
        RECT  1.930 0.705 2.240 0.820 ;
        RECT  1.850 0.705 1.930 1.035 ;
        RECT  0.735 0.705 1.850 0.820 ;
        RECT  0.735 0.345 1.590 0.415 ;
        RECT  0.525 0.345 0.735 0.820 ;
        RECT  0.130 0.345 0.525 0.415 ;
        RECT  0.210 0.700 0.525 0.820 ;
        RECT  0.050 0.255 0.130 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.390 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 -0.115 3.360 0.115 ;
        RECT  3.010 -0.115 3.150 0.275 ;
        RECT  2.750 -0.115 3.010 0.115 ;
        RECT  2.610 -0.115 2.750 0.275 ;
        RECT  0.000 -0.115 2.610 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.145 3.360 1.375 ;
        RECT  3.220 0.705 3.320 1.375 ;
        RECT  2.940 1.145 3.220 1.375 ;
        RECT  2.820 0.890 2.940 1.375 ;
        RECT  2.540 1.145 2.820 1.375 ;
        RECT  2.420 0.890 2.540 1.375 ;
        RECT  2.140 1.145 2.420 1.375 ;
        RECT  2.020 0.890 2.140 1.375 ;
        RECT  1.745 1.145 2.020 1.375 ;
        RECT  1.675 0.895 1.745 1.375 ;
        RECT  1.410 1.145 1.675 1.375 ;
        RECT  1.290 1.030 1.410 1.375 ;
        RECT  1.050 1.145 1.290 1.375 ;
        RECT  0.930 1.030 1.050 1.375 ;
        RECT  0.000 1.145 0.930 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.040 0.705 3.120 1.035 ;
        RECT  2.720 0.705 3.040 0.820 ;
        RECT  2.640 0.705 2.720 1.035 ;
        RECT  2.320 0.705 2.640 0.820 ;
        RECT  2.240 0.705 2.320 1.035 ;
        RECT  1.930 0.705 2.240 0.820 ;
        RECT  1.850 0.705 1.930 1.035 ;
        RECT  0.805 0.705 1.850 0.820 ;
        RECT  0.805 0.345 1.590 0.415 ;
        RECT  0.130 0.345 0.455 0.415 ;
        RECT  0.210 0.700 0.455 0.820 ;
        RECT  0.050 0.255 0.130 0.415 ;
        RECT  3.230 0.255 3.310 0.415 ;
        RECT  2.920 0.345 3.230 0.415 ;
        RECT  2.840 0.185 2.920 0.415 ;
        RECT  2.520 0.345 2.840 0.415 ;
        RECT  2.440 0.185 2.520 0.415 ;
        RECT  1.750 0.345 2.440 0.415 ;
        RECT  0.210 0.205 2.340 0.275 ;
        RECT  1.670 0.345 1.750 0.475 ;
        RECT  0.130 0.890 1.590 0.960 ;
        RECT  0.055 0.735 0.130 1.035 ;
    END
END OAI211D4BWP

MACRO OAI21D0BWP
    CLASS CORE ;
    FOREIGN OAI21D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0723 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.935 0.545 1.055 ;
        RECT  0.455 0.345 0.525 1.055 ;
        RECT  0.240 0.345 0.455 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.625 ;
        RECT  0.610 0.540 0.715 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.620 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.840 0.115 ;
        RECT  0.650 -0.115 0.730 0.280 ;
        RECT  0.000 -0.115 0.650 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 1.145 0.840 1.375 ;
        RECT  0.655 0.925 0.725 1.375 ;
        RECT  0.130 1.145 0.655 1.375 ;
        RECT  0.050 0.925 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.205 0.570 0.275 ;
        RECT  0.050 0.205 0.130 0.325 ;
    END
END OAI21D0BWP

MACRO OAI21D1BWP
    CLASS CORE ;
    FOREIGN OAI21D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1194 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.695 0.560 1.075 ;
        RECT  0.455 0.345 0.525 1.075 ;
        RECT  0.240 0.345 0.455 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.540 0.735 0.620 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.115 0.840 0.115 ;
        RECT  0.655 -0.115 0.725 0.415 ;
        RECT  0.000 -0.115 0.655 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.640 0.850 0.740 1.375 ;
        RECT  0.140 1.145 0.640 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.145 0.205 0.570 0.275 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OAI21D1BWP

MACRO OAI21D2BWP
    CLASS CORE ;
    FOREIGN OAI21D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2344 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.845 1.225 1.045 ;
        RECT  0.525 0.845 1.135 0.915 ;
        RECT  0.665 0.345 1.050 0.415 ;
        RECT  0.570 0.345 0.665 0.490 ;
        RECT  0.395 0.420 0.570 0.490 ;
        RECT  0.415 0.845 0.525 1.075 ;
        RECT  0.395 0.845 0.415 0.915 ;
        RECT  0.315 0.420 0.395 0.915 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.775 ;
        RECT  0.665 0.705 1.015 0.775 ;
        RECT  0.585 0.560 0.665 0.775 ;
        RECT  0.490 0.560 0.585 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 -0.115 1.260 0.115 ;
        RECT  0.210 -0.115 0.330 0.210 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.870 1.145 1.260 1.375 ;
        RECT  0.750 0.985 0.870 1.375 ;
        RECT  0.330 1.145 0.750 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.130 0.205 1.210 0.375 ;
        RECT  0.485 0.205 1.130 0.275 ;
        RECT  0.415 0.205 0.485 0.350 ;
        RECT  0.130 0.280 0.415 0.350 ;
        RECT  0.050 0.230 0.130 0.350 ;
    END
END OAI21D2BWP

MACRO OAI21D4BWP
    CLASS CORE ;
    FOREIGN OAI21D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.695 2.290 0.985 ;
        RECT  1.930 0.695 2.210 0.800 ;
        RECT  1.850 0.695 1.930 0.985 ;
        RECT  0.735 0.695 1.850 0.800 ;
        RECT  0.735 0.345 1.410 0.415 ;
        RECT  0.525 0.345 0.735 0.800 ;
        RECT  0.210 0.345 0.525 0.415 ;
        RECT  0.210 0.695 0.525 0.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.385 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 -0.115 2.520 0.115 ;
        RECT  2.380 -0.115 2.480 0.415 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.020 -0.115 2.120 0.275 ;
        RECT  1.760 -0.115 2.020 0.115 ;
        RECT  1.660 -0.115 1.760 0.275 ;
        RECT  0.000 -0.115 1.660 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.710 2.480 1.375 ;
        RECT  2.130 1.145 2.380 1.375 ;
        RECT  2.010 0.870 2.130 1.375 ;
        RECT  1.750 1.145 2.010 1.375 ;
        RECT  1.670 0.870 1.750 1.375 ;
        RECT  1.400 1.145 1.670 1.375 ;
        RECT  1.300 1.010 1.400 1.375 ;
        RECT  1.040 1.145 1.300 1.375 ;
        RECT  0.940 1.010 1.040 1.375 ;
        RECT  0.000 1.145 0.940 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.210 0.695 2.290 0.985 ;
        RECT  1.930 0.695 2.210 0.800 ;
        RECT  1.850 0.695 1.930 0.985 ;
        RECT  0.805 0.695 1.850 0.800 ;
        RECT  0.805 0.345 1.410 0.415 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.210 0.695 0.455 0.800 ;
        RECT  2.190 0.185 2.310 0.415 ;
        RECT  1.490 0.205 1.570 0.415 ;
        RECT  0.130 0.205 1.490 0.275 ;
        RECT  1.230 0.870 1.470 0.940 ;
        RECT  1.110 0.870 1.230 1.075 ;
        RECT  0.870 0.870 1.110 0.940 ;
        RECT  0.750 0.870 0.870 1.075 ;
        RECT  0.510 0.870 0.750 0.940 ;
        RECT  0.390 0.870 0.510 1.075 ;
        RECT  0.125 0.870 0.390 0.940 ;
        RECT  0.050 0.205 0.130 0.395 ;
        RECT  0.055 0.735 0.125 1.035 ;
        RECT  1.930 0.345 2.190 0.415 ;
        RECT  1.850 0.185 1.930 0.415 ;
        RECT  1.570 0.345 1.850 0.415 ;
        RECT  1.470 0.870 1.590 1.075 ;
    END
END OAI21D4BWP

MACRO OAI221D0BWP
    CLASS CORE ;
    FOREIGN OAI221D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0730 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.845 1.025 1.060 ;
        RECT  0.385 0.845 0.955 0.915 ;
        RECT  0.330 0.495 0.385 0.915 ;
        RECT  0.315 0.335 0.330 0.915 ;
        RECT  0.260 0.335 0.315 0.565 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.210 0.335 0.260 0.405 ;
        RECT  0.035 0.845 0.125 1.060 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.635 1.225 0.905 ;
        RECT  1.040 0.635 1.155 0.705 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.630 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.415 ;
        RECT  0.000 -0.115 1.130 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.260 1.375 ;
        RECT  1.120 0.985 1.220 1.375 ;
        RECT  0.680 1.145 1.120 1.375 ;
        RECT  0.580 0.985 0.680 1.375 ;
        RECT  0.500 1.145 0.580 1.375 ;
        RECT  0.400 0.985 0.500 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.195 1.025 0.415 ;
        RECT  0.560 0.195 0.955 0.265 ;
        RECT  0.480 0.345 0.870 0.415 ;
        RECT  0.410 0.195 0.480 0.415 ;
        RECT  0.125 0.195 0.410 0.265 ;
        RECT  0.055 0.195 0.125 0.415 ;
    END
END OAI221D0BWP

MACRO OAI221D1BWP
    CLASS CORE ;
    FOREIGN OAI221D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1459 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.940 0.835 1.040 1.075 ;
        RECT  0.385 0.835 0.940 0.905 ;
        RECT  0.315 0.355 0.385 0.905 ;
        RECT  0.210 0.355 0.315 0.425 ;
        RECT  0.140 0.835 0.315 0.905 ;
        RECT  0.035 0.695 0.140 1.075 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.905 ;
        RECT  1.070 0.495 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.260 0.115 ;
        RECT  1.120 -0.115 1.220 0.425 ;
        RECT  0.000 -0.115 1.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.260 1.375 ;
        RECT  1.120 0.985 1.220 1.375 ;
        RECT  0.680 1.145 1.120 1.375 ;
        RECT  0.580 0.975 0.680 1.375 ;
        RECT  0.500 1.145 0.580 1.375 ;
        RECT  0.400 0.975 0.500 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 0.185 1.040 0.425 ;
        RECT  0.570 0.355 0.940 0.425 ;
        RECT  0.140 0.205 0.870 0.275 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END OAI221D1BWP

MACRO OAI221D2BWP
    CLASS CORE ;
    FOREIGN OAI221D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3248 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.975 2.030 1.045 ;
        RECT  0.890 0.545 0.945 1.045 ;
        RECT  0.875 0.345 0.890 1.045 ;
        RECT  0.820 0.345 0.875 0.615 ;
        RECT  0.145 0.975 0.875 1.045 ;
        RECT  0.130 0.345 0.820 0.415 ;
        RECT  0.035 0.975 0.145 1.075 ;
        RECT  0.035 0.215 0.130 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.945 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.385 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.495 1.695 0.640 ;
        RECT  1.575 0.495 1.645 0.905 ;
        RECT  1.085 0.835 1.575 0.905 ;
        RECT  1.085 0.545 1.150 0.615 ;
        RECT  1.015 0.545 1.085 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.495 0.750 0.640 ;
        RECT  0.595 0.495 0.685 0.905 ;
        RECT  0.245 0.835 0.595 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.240 0.115 ;
        RECT  1.880 -0.115 2.000 0.275 ;
        RECT  0.000 -0.115 1.880 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.700 2.190 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.720 1.115 1.840 1.375 ;
        RECT  1.070 1.145 1.720 1.375 ;
        RECT  0.950 1.115 1.070 1.375 ;
        RECT  0.520 1.145 0.950 1.375 ;
        RECT  0.400 1.115 0.520 1.375 ;
        RECT  0.000 1.145 0.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.100 0.185 2.200 0.425 ;
        RECT  1.770 0.355 2.100 0.425 ;
        RECT  1.690 0.190 1.770 0.425 ;
        RECT  1.060 0.355 1.690 0.425 ;
        RECT  0.210 0.205 1.610 0.275 ;
        RECT  0.960 0.355 1.060 0.455 ;
    END
END OAI221D2BWP

MACRO OAI221D4BWP
    CLASS CORE ;
    FOREIGN OAI221D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2078 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.685 1.820 0.800 ;
        RECT  1.700 0.185 1.770 0.465 ;
        RECT  1.575 0.350 1.700 0.465 ;
        RECT  1.410 0.350 1.575 0.800 ;
        RECT  1.365 0.185 1.410 0.800 ;
        RECT  1.330 0.185 1.365 0.465 ;
        RECT  1.350 0.685 1.365 0.800 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.230 0.640 ;
        RECT  1.085 0.520 1.155 0.640 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.975 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.980 -0.115 2.240 0.115 ;
        RECT  1.900 -0.115 1.980 0.300 ;
        RECT  1.610 -0.115 1.900 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  1.230 -0.115 1.490 0.115 ;
        RECT  1.150 -0.115 1.230 0.275 ;
        RECT  0.000 -0.115 1.150 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 1.145 2.240 1.375 ;
        RECT  1.900 1.010 2.020 1.375 ;
        RECT  1.650 1.145 1.900 1.375 ;
        RECT  1.530 1.010 1.650 1.375 ;
        RECT  1.280 1.145 1.530 1.375 ;
        RECT  1.160 1.010 1.280 1.375 ;
        RECT  0.720 1.145 1.160 1.375 ;
        RECT  0.600 1.115 0.720 1.375 ;
        RECT  0.495 1.145 0.600 1.375 ;
        RECT  0.425 0.975 0.495 1.375 ;
        RECT  0.000 1.145 0.425 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.685 1.820 0.800 ;
        RECT  1.700 0.185 1.770 0.465 ;
        RECT  1.645 0.350 1.700 0.465 ;
        RECT  2.120 0.185 2.190 1.070 ;
        RECT  2.115 0.185 2.120 0.440 ;
        RECT  1.910 0.370 2.115 0.440 ;
        RECT  1.980 0.520 2.050 0.940 ;
        RECT  1.065 0.870 1.980 0.940 ;
        RECT  1.840 0.370 1.910 0.615 ;
        RECT  1.760 0.545 1.840 0.615 ;
        RECT  0.590 0.345 1.070 0.415 ;
        RECT  0.995 0.870 1.065 1.045 ;
        RECT  0.645 0.975 0.995 1.045 ;
        RECT  0.130 0.205 0.890 0.275 ;
        RECT  0.575 0.835 0.645 1.045 ;
        RECT  0.385 0.835 0.575 0.905 ;
        RECT  0.315 0.345 0.385 0.905 ;
        RECT  0.210 0.345 0.315 0.415 ;
        RECT  0.310 0.835 0.315 0.905 ;
        RECT  0.240 0.835 0.310 1.045 ;
        RECT  0.125 0.975 0.240 1.045 ;
        RECT  0.050 0.205 0.130 0.395 ;
        RECT  0.055 0.925 0.125 1.045 ;
    END
END OAI221D4BWP

MACRO OAI221XD4BWP
    CLASS CORE ;
    FOREIGN OAI221XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5180 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.345 3.970 0.415 ;
        RECT  2.975 0.705 3.250 0.820 ;
        RECT  2.765 0.345 2.975 0.820 ;
        RECT  0.685 0.705 2.765 0.820 ;
        RECT  0.615 0.705 0.685 1.035 ;
        RECT  0.325 0.705 0.615 0.820 ;
        RECT  0.255 0.705 0.325 1.035 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.675 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.645 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 4.025 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.325 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 -0.115 4.200 0.115 ;
        RECT  0.780 -0.115 0.880 0.275 ;
        RECT  0.510 -0.115 0.780 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.160 -0.115 0.430 0.115 ;
        RECT  0.060 -0.115 0.160 0.415 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.145 4.200 1.375 ;
        RECT  3.870 0.855 3.950 1.375 ;
        RECT  3.590 1.145 3.870 1.375 ;
        RECT  3.510 0.855 3.590 1.375 ;
        RECT  1.610 1.145 3.510 1.375 ;
        RECT  1.490 1.030 1.610 1.375 ;
        RECT  1.250 1.145 1.490 1.375 ;
        RECT  1.130 1.030 1.250 1.375 ;
        RECT  0.870 1.145 1.130 1.375 ;
        RECT  0.790 0.895 0.870 1.375 ;
        RECT  0.510 1.145 0.790 1.375 ;
        RECT  0.430 0.895 0.510 1.375 ;
        RECT  0.145 1.145 0.430 1.375 ;
        RECT  0.075 0.705 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.345 3.970 0.415 ;
        RECT  3.045 0.705 3.250 0.820 ;
        RECT  0.685 0.705 2.695 0.820 ;
        RECT  0.615 0.705 0.685 1.035 ;
        RECT  0.325 0.705 0.615 0.820 ;
        RECT  0.255 0.705 0.325 1.035 ;
        RECT  4.050 0.195 4.130 0.395 ;
        RECT  4.050 0.715 4.130 1.035 ;
        RECT  2.685 0.195 4.050 0.265 ;
        RECT  3.770 0.715 4.050 0.785 ;
        RECT  3.690 0.715 3.770 1.025 ;
        RECT  3.410 0.715 3.690 0.785 ;
        RECT  3.330 0.715 3.410 1.030 ;
        RECT  2.590 0.960 3.330 1.030 ;
        RECT  2.615 0.195 2.685 0.435 ;
        RECT  2.485 0.195 2.615 0.265 ;
        RECT  0.950 0.890 2.510 0.960 ;
        RECT  2.415 0.195 2.485 0.435 ;
        RECT  0.950 0.195 2.415 0.265 ;
        RECT  0.690 0.345 2.335 0.415 ;
        RECT  0.610 0.255 0.690 0.415 ;
        RECT  0.330 0.345 0.610 0.415 ;
        RECT  0.250 0.255 0.330 0.415 ;
    END
END OAI221XD4BWP

MACRO OAI222D0BWP
    CLASS CORE ;
    FOREIGN OAI222D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0935 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.985 1.150 1.055 ;
        RECT  0.455 0.345 0.525 1.055 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.225 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.625 ;
        RECT  1.320 0.545 1.435 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.905 ;
        RECT  0.810 0.635 0.875 0.705 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 -0.115 1.540 0.115 ;
        RECT  1.395 -0.115 1.505 0.275 ;
        RECT  1.140 -0.115 1.395 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.000 -0.115 1.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.910 1.490 1.375 ;
        RECT  0.940 1.145 1.410 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.130 1.145 0.820 1.375 ;
        RECT  0.050 0.910 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.230 0.185 1.310 0.415 ;
        RECT  0.660 0.345 1.230 0.415 ;
        RECT  0.130 0.195 0.970 0.265 ;
        RECT  0.050 0.195 0.130 0.325 ;
    END
END OAI222D0BWP

MACRO OAI222D1BWP
    CLASS CORE ;
    FOREIGN OAI222D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1767 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.840 1.150 1.055 ;
        RECT  0.525 0.985 1.030 1.055 ;
        RECT  0.455 0.345 0.525 1.075 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.225 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.625 ;
        RECT  1.320 0.545 1.435 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.545 0.945 0.905 ;
        RECT  0.790 0.545 0.875 0.615 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 -0.115 1.540 0.115 ;
        RECT  1.395 -0.115 1.505 0.275 ;
        RECT  1.140 -0.115 1.395 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.000 -0.115 1.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.705 1.500 1.375 ;
        RECT  0.970 1.145 1.400 1.375 ;
        RECT  0.850 1.125 0.970 1.375 ;
        RECT  0.140 1.145 0.850 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.205 1.325 0.415 ;
        RECT  0.650 0.345 1.210 0.415 ;
        RECT  0.130 0.195 0.950 0.265 ;
        RECT  0.050 0.195 0.130 0.395 ;
    END
END OAI222D1BWP

MACRO OAI222D2BWP
    CLASS CORE ;
    FOREIGN OAI222D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.3166 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.845 2.130 1.050 ;
        RECT  1.390 0.845 1.995 0.915 ;
        RECT  1.295 0.845 1.390 1.075 ;
        RECT  0.945 0.845 1.295 0.915 ;
        RECT  0.875 0.545 0.945 0.915 ;
        RECT  0.870 0.545 0.875 0.615 ;
        RECT  0.850 0.845 0.875 0.915 ;
        RECT  0.800 0.345 0.870 0.615 ;
        RECT  0.735 0.845 0.850 1.075 ;
        RECT  0.130 0.345 0.800 0.415 ;
        RECT  0.125 0.845 0.735 0.915 ;
        RECT  0.050 0.215 0.130 0.415 ;
        RECT  0.050 0.845 0.125 1.045 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.205 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.495 2.395 0.640 ;
        RECT  2.275 0.495 2.345 0.765 ;
        RECT  1.925 0.695 2.275 0.765 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.790 0.495 1.855 0.640 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.775 ;
        RECT  1.105 0.705 1.575 0.775 ;
        RECT  1.015 0.520 1.105 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.730 0.640 ;
        RECT  0.595 0.495 0.665 0.775 ;
        RECT  0.245 0.705 0.595 0.775 ;
        RECT  0.155 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.310 -0.115 2.520 0.115 ;
        RECT  2.190 -0.115 2.310 0.275 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.275 ;
        RECT  0.000 -0.115 1.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.145 2.520 1.375 ;
        RECT  2.380 0.845 2.480 1.375 ;
        RECT  1.770 1.145 2.380 1.375 ;
        RECT  1.650 0.985 1.770 1.375 ;
        RECT  1.050 1.145 1.650 1.375 ;
        RECT  0.930 0.985 1.050 1.375 ;
        RECT  0.510 1.145 0.930 1.375 ;
        RECT  0.390 0.985 0.510 1.375 ;
        RECT  0.000 1.145 0.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.255 2.470 0.415 ;
        RECT  2.110 0.345 2.390 0.415 ;
        RECT  2.030 0.185 2.110 0.415 ;
        RECT  1.750 0.345 2.030 0.415 ;
        RECT  1.670 0.185 1.750 0.415 ;
        RECT  1.040 0.345 1.670 0.415 ;
        RECT  0.210 0.205 1.590 0.275 ;
        RECT  0.940 0.345 1.040 0.445 ;
    END
END OAI222D2BWP

MACRO OAI222D4BWP
    CLASS CORE ;
    FOREIGN OAI222D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.785 2.090 0.905 ;
        RECT  1.995 0.185 2.065 0.465 ;
        RECT  1.855 0.350 1.995 0.465 ;
        RECT  1.685 0.350 1.855 0.905 ;
        RECT  1.645 0.185 1.685 0.905 ;
        RECT  1.615 0.185 1.645 0.465 ;
        RECT  1.590 0.785 1.645 0.905 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.225 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.510 0.625 ;
        RECT  1.320 0.545 1.435 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.810 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.540 0.880 0.615 ;
        RECT  0.735 0.540 0.805 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.350 0.525 0.640 ;
        RECT  0.400 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.180 -0.115 2.260 0.300 ;
        RECT  1.900 -0.115 2.180 0.115 ;
        RECT  1.780 -0.115 1.900 0.270 ;
        RECT  1.510 -0.115 1.780 0.115 ;
        RECT  1.410 -0.115 1.510 0.275 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.000 -0.115 1.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.160 1.125 2.280 1.375 ;
        RECT  1.900 1.145 2.160 1.375 ;
        RECT  1.780 1.125 1.900 1.375 ;
        RECT  1.520 1.145 1.780 1.375 ;
        RECT  1.400 1.125 1.520 1.375 ;
        RECT  0.970 1.145 1.400 1.375 ;
        RECT  0.850 1.125 0.970 1.375 ;
        RECT  0.150 1.145 0.850 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.785 2.090 0.905 ;
        RECT  1.995 0.185 2.065 0.465 ;
        RECT  1.925 0.350 1.995 0.465 ;
        RECT  2.460 0.370 2.485 0.915 ;
        RECT  2.450 0.370 2.460 1.075 ;
        RECT  2.415 0.255 2.450 1.075 ;
        RECT  2.370 0.255 2.415 0.440 ;
        RECT  2.360 0.835 2.415 1.075 ;
        RECT  2.205 0.370 2.370 0.440 ;
        RECT  2.275 0.520 2.345 0.765 ;
        RECT  2.260 0.695 2.275 0.765 ;
        RECT  2.190 0.695 2.260 1.055 ;
        RECT  2.135 0.370 2.205 0.615 ;
        RECT  0.330 0.985 2.190 1.055 ;
        RECT  1.990 0.545 2.135 0.615 ;
        RECT  1.210 0.205 1.330 0.415 ;
        RECT  0.640 0.345 1.210 0.415 ;
        RECT  0.150 0.195 0.950 0.265 ;
        RECT  0.260 0.335 0.330 1.055 ;
        RECT  0.070 0.195 0.150 0.395 ;
    END
END OAI222D4BWP

MACRO OAI222XD4BWP
    CLASS CORE ;
    FOREIGN OAI222XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5180 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.345 4.670 0.415 ;
        RECT  3.830 0.705 3.950 0.925 ;
        RECT  3.675 0.705 3.830 0.820 ;
        RECT  3.605 0.345 3.675 0.820 ;
        RECT  3.470 0.345 3.605 0.925 ;
        RECT  3.465 0.345 3.470 0.820 ;
        RECT  1.430 0.705 3.465 0.820 ;
        RECT  1.310 0.705 1.430 0.925 ;
        RECT  1.070 0.705 1.310 0.820 ;
        RECT  0.950 0.705 1.070 0.925 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.665 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.565 0.495 3.055 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.350 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.725 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.495 4.025 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.600 -0.115 4.900 0.115 ;
        RECT  1.500 -0.115 1.600 0.275 ;
        RECT  1.230 -0.115 1.500 0.115 ;
        RECT  1.150 -0.115 1.230 0.275 ;
        RECT  0.870 -0.115 1.150 0.115 ;
        RECT  0.790 -0.115 0.870 0.275 ;
        RECT  0.510 -0.115 0.790 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.650 1.145 4.900 1.375 ;
        RECT  4.570 0.855 4.650 1.375 ;
        RECT  4.290 1.145 4.570 1.375 ;
        RECT  4.210 0.855 4.290 1.375 ;
        RECT  2.330 1.145 4.210 1.375 ;
        RECT  2.210 1.030 2.330 1.375 ;
        RECT  1.970 1.145 2.210 1.375 ;
        RECT  1.850 1.030 1.970 1.375 ;
        RECT  0.690 1.145 1.850 1.375 ;
        RECT  0.610 0.855 0.690 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.250 0.855 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.345 4.670 0.415 ;
        RECT  3.830 0.705 3.950 0.925 ;
        RECT  3.745 0.705 3.830 0.820 ;
        RECT  1.430 0.705 3.395 0.820 ;
        RECT  1.310 0.705 1.430 0.925 ;
        RECT  1.070 0.705 1.310 0.820 ;
        RECT  0.950 0.705 1.070 0.925 ;
        RECT  4.750 0.195 4.830 0.395 ;
        RECT  4.750 0.715 4.830 1.045 ;
        RECT  3.385 0.195 4.750 0.265 ;
        RECT  4.470 0.715 4.750 0.785 ;
        RECT  4.390 0.715 4.470 1.045 ;
        RECT  4.110 0.715 4.390 0.785 ;
        RECT  4.030 0.715 4.110 1.065 ;
        RECT  3.290 0.995 4.030 1.065 ;
        RECT  3.315 0.195 3.385 0.460 ;
        RECT  3.205 0.195 3.315 0.265 ;
        RECT  3.130 0.890 3.210 1.025 ;
        RECT  3.135 0.195 3.205 0.460 ;
        RECT  1.670 0.195 3.135 0.265 ;
        RECT  1.670 0.890 3.130 0.960 ;
        RECT  1.410 0.345 3.050 0.415 ;
        RECT  1.510 0.915 1.590 1.065 ;
        RECT  0.870 0.995 1.510 1.065 ;
        RECT  1.330 0.255 1.410 0.415 ;
        RECT  1.050 0.345 1.330 0.415 ;
        RECT  0.970 0.255 1.050 0.415 ;
        RECT  0.690 0.345 0.970 0.415 ;
        RECT  0.790 0.715 0.870 1.065 ;
        RECT  0.510 0.715 0.790 0.785 ;
        RECT  0.610 0.255 0.690 0.415 ;
        RECT  0.330 0.345 0.610 0.415 ;
        RECT  0.430 0.715 0.510 1.035 ;
        RECT  0.150 0.715 0.430 0.785 ;
        RECT  0.250 0.255 0.330 0.415 ;
        RECT  0.070 0.715 0.150 1.035 ;
    END
END OAI222XD4BWP

MACRO OAI22D0BWP
    CLASS CORE ;
    FOREIGN OAI22D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0783 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.915 0.925 1.045 ;
        RECT  0.525 0.975 0.855 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.125 0.975 0.455 1.045 ;
        RECT  0.055 0.915 0.125 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.635 0.685 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.760 0.545 0.875 0.615 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.000 -0.115 0.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.145 0.980 1.375 ;
        RECT  0.440 1.115 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.205 0.940 0.305 ;
        RECT  0.145 0.205 0.840 0.275 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OAI22D0BWP

MACRO OAI22D1BWP
    CLASS CORE ;
    FOREIGN OAI22D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1398 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.915 0.925 1.045 ;
        RECT  0.525 0.975 0.855 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.210 0.345 0.455 0.415 ;
        RECT  0.125 0.975 0.455 1.045 ;
        RECT  0.055 0.915 0.125 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.685 0.670 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.760 0.545 0.875 0.615 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.135 ;
        RECT  0.000 -0.115 0.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.145 0.980 1.375 ;
        RECT  0.440 1.115 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.205 0.930 0.395 ;
        RECT  0.130 0.205 0.850 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OAI22D1BWP

MACRO OAI22D2BWP
    CLASS CORE ;
    FOREIGN OAI22D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 0.345 1.470 0.415 ;
        RECT  0.805 0.985 1.290 1.055 ;
        RECT  0.810 0.345 0.880 0.835 ;
        RECT  0.805 0.765 0.810 0.835 ;
        RECT  0.735 0.765 0.805 1.055 ;
        RECT  0.390 0.985 0.735 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.740 0.640 ;
        RECT  0.595 0.520 0.665 0.905 ;
        RECT  0.245 0.835 0.595 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.525 0.905 ;
        RECT  1.085 0.835 1.435 0.905 ;
        RECT  1.010 0.495 1.085 0.905 ;
        RECT  0.950 0.495 1.010 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.115 1.680 0.115 ;
        RECT  0.600 -0.115 0.720 0.135 ;
        RECT  0.330 -0.115 0.600 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.145 1.680 1.375 ;
        RECT  1.535 0.985 1.645 1.375 ;
        RECT  0.900 1.145 1.535 1.375 ;
        RECT  0.780 1.135 0.900 1.375 ;
        RECT  0.145 1.145 0.780 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.550 0.205 1.630 0.395 ;
        RECT  0.705 0.205 1.550 0.275 ;
        RECT  0.625 0.205 0.705 0.415 ;
        RECT  0.485 0.345 0.625 0.415 ;
        RECT  0.415 0.185 0.485 0.415 ;
        RECT  0.130 0.345 0.415 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OAI22D2BWP

MACRO OAI22D4BWP
    CLASS CORE ;
    FOREIGN OAI22D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4196 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.805 3.120 0.875 ;
        RECT  1.660 0.540 1.740 0.875 ;
        RECT  1.540 0.540 1.660 0.620 ;
        RECT  1.460 0.345 1.540 0.620 ;
        RECT  0.735 0.345 1.460 0.415 ;
        RECT  0.525 0.345 0.735 0.900 ;
        RECT  0.230 0.345 0.525 0.415 ;
        RECT  0.230 0.775 0.525 0.900 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.385 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.115 3.360 0.115 ;
        RECT  3.010 -0.115 3.110 0.275 ;
        RECT  2.730 -0.115 3.010 0.115 ;
        RECT  2.630 -0.115 2.730 0.275 ;
        RECT  2.350 -0.115 2.630 0.115 ;
        RECT  2.250 -0.115 2.350 0.275 ;
        RECT  1.970 -0.115 2.250 0.115 ;
        RECT  1.870 -0.115 1.970 0.275 ;
        RECT  0.000 -0.115 1.870 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.145 3.360 1.375 ;
        RECT  2.240 1.115 2.360 1.375 ;
        RECT  1.980 1.145 2.240 1.375 ;
        RECT  1.860 1.115 1.980 1.375 ;
        RECT  1.410 1.145 1.860 1.375 ;
        RECT  1.330 0.860 1.410 1.375 ;
        RECT  1.045 1.145 1.330 1.375 ;
        RECT  0.975 0.860 1.045 1.375 ;
        RECT  0.000 1.145 0.975 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 0.805 3.120 0.875 ;
        RECT  1.660 0.540 1.740 0.875 ;
        RECT  1.540 0.540 1.660 0.620 ;
        RECT  1.460 0.345 1.540 0.620 ;
        RECT  0.805 0.345 1.460 0.415 ;
        RECT  0.230 0.345 0.455 0.415 ;
        RECT  0.230 0.775 0.455 0.900 ;
        RECT  3.210 0.255 3.290 0.415 ;
        RECT  3.210 0.735 3.290 1.045 ;
        RECT  2.905 0.345 3.210 0.415 ;
        RECT  1.670 0.975 3.210 1.045 ;
        RECT  2.835 0.185 2.905 0.415 ;
        RECT  2.525 0.345 2.835 0.415 ;
        RECT  2.455 0.185 2.525 0.415 ;
        RECT  2.145 0.345 2.455 0.415 ;
        RECT  2.075 0.185 2.145 0.415 ;
        RECT  1.800 0.345 2.075 0.415 ;
        RECT  1.730 0.205 1.800 0.415 ;
        RECT  0.150 0.205 1.730 0.275 ;
        RECT  1.510 0.710 1.590 1.035 ;
        RECT  1.230 0.710 1.510 0.780 ;
        RECT  1.150 0.710 1.230 1.035 ;
        RECT  0.905 0.710 1.150 0.780 ;
        RECT  0.835 0.710 0.905 1.045 ;
        RECT  0.150 0.975 0.835 1.045 ;
        RECT  0.070 0.205 0.150 0.395 ;
        RECT  0.070 0.735 0.150 1.045 ;
    END
END OAI22D4BWP

MACRO OAI31D0BWP
    CLASS CORE ;
    FOREIGN OAI31D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0851 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.970 0.750 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.135 0.345 0.455 0.415 ;
        RECT  0.035 0.185 0.135 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.625 ;
        RECT  0.750 0.545 0.875 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.680 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.635 0.385 0.950 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 -0.115 0.980 0.115 ;
        RECT  0.825 -0.115 0.935 0.275 ;
        RECT  0.000 -0.115 0.825 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.145 0.980 1.375 ;
        RECT  0.845 0.940 0.915 1.375 ;
        RECT  0.135 1.145 0.845 1.375 ;
        RECT  0.065 0.940 0.135 1.375 ;
        RECT  0.000 1.145 0.065 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.230 0.205 0.750 0.275 ;
    END
END OAI31D0BWP

MACRO OAI31D1BWP
    CLASS CORE ;
    FOREIGN OAI31D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1493 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.970 0.750 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.135 0.345 0.455 0.415 ;
        RECT  0.065 0.215 0.135 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.625 ;
        RECT  0.750 0.545 0.875 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 -0.115 0.980 0.115 ;
        RECT  0.825 -0.115 0.935 0.275 ;
        RECT  0.000 -0.115 0.825 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.830 0.705 0.930 1.375 ;
        RECT  0.150 1.145 0.830 1.375 ;
        RECT  0.050 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.630 0.205 0.750 0.415 ;
        RECT  0.230 0.205 0.630 0.275 ;
    END
END OAI31D1BWP

MACRO OAI31D2BWP
    CLASS CORE ;
    FOREIGN OAI31D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.735 1.450 1.055 ;
        RECT  1.295 0.345 1.365 1.055 ;
        RECT  0.210 0.345 1.295 0.415 ;
        RECT  0.570 0.985 1.295 1.055 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.355 1.645 0.625 ;
        RECT  1.440 0.545 1.555 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.775 ;
        RECT  0.410 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.410 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.135 0.640 ;
        RECT  1.015 0.495 1.085 0.915 ;
        RECT  0.245 0.845 1.015 0.915 ;
        RECT  0.155 0.495 0.245 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.440 -0.115 1.680 0.115 ;
        RECT  1.320 -0.115 1.440 0.135 ;
        RECT  0.000 -0.115 1.320 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.145 1.680 1.375 ;
        RECT  1.540 0.705 1.640 1.375 ;
        RECT  1.260 1.145 1.540 1.375 ;
        RECT  1.140 1.125 1.260 1.375 ;
        RECT  0.145 1.145 1.140 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.185 1.645 0.285 ;
        RECT  0.130 0.205 1.535 0.275 ;
        RECT  0.050 0.205 0.130 0.385 ;
    END
END OAI31D2BWP

MACRO OAI31D4BWP
    CLASS CORE ;
    FOREIGN OAI31D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.5374 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.045 0.695 3.115 1.035 ;
        RECT  2.715 0.695 3.045 0.765 ;
        RECT  2.645 0.695 2.715 1.035 ;
        RECT  0.735 0.695 2.645 0.765 ;
        RECT  0.735 0.345 2.350 0.415 ;
        RECT  0.690 0.345 0.735 0.765 ;
        RECT  0.570 0.345 0.690 0.925 ;
        RECT  0.525 0.345 0.570 0.765 ;
        RECT  0.125 0.345 0.525 0.415 ;
        RECT  0.330 0.695 0.525 0.765 ;
        RECT  0.210 0.695 0.330 0.925 ;
        RECT  0.055 0.255 0.125 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.185 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.385 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.140 -0.115 3.360 0.115 ;
        RECT  3.020 -0.115 3.140 0.275 ;
        RECT  2.740 -0.115 3.020 0.115 ;
        RECT  2.620 -0.115 2.740 0.275 ;
        RECT  0.000 -0.115 2.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.145 3.360 1.375 ;
        RECT  3.220 0.705 3.320 1.375 ;
        RECT  2.915 1.145 3.220 1.375 ;
        RECT  2.845 0.845 2.915 1.375 ;
        RECT  2.515 1.145 2.845 1.375 ;
        RECT  2.445 0.845 2.515 1.375 ;
        RECT  2.140 1.145 2.445 1.375 ;
        RECT  2.020 0.990 2.140 1.375 ;
        RECT  0.000 1.145 2.020 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.695 3.115 1.035 ;
        RECT  2.715 0.695 3.045 0.765 ;
        RECT  2.645 0.695 2.715 1.035 ;
        RECT  0.805 0.695 2.645 0.765 ;
        RECT  0.805 0.345 2.350 0.415 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.330 0.695 0.455 0.765 ;
        RECT  0.210 0.695 0.330 0.925 ;
        RECT  0.055 0.255 0.125 0.415 ;
        RECT  3.235 0.255 3.305 0.415 ;
        RECT  2.915 0.345 3.235 0.415 ;
        RECT  2.845 0.185 2.915 0.415 ;
        RECT  2.515 0.345 2.845 0.415 ;
        RECT  2.445 0.205 2.515 0.415 ;
        RECT  0.210 0.205 2.445 0.275 ;
        RECT  2.220 0.845 2.340 1.045 ;
        RECT  1.925 0.845 2.220 0.915 ;
        RECT  1.855 0.845 1.925 1.075 ;
        RECT  0.930 0.845 1.855 0.915 ;
        RECT  0.845 0.995 1.590 1.065 ;
        RECT  0.775 0.835 0.845 1.065 ;
        RECT  0.485 0.995 0.775 1.065 ;
        RECT  0.415 0.835 0.485 1.065 ;
        RECT  0.130 0.995 0.415 1.065 ;
        RECT  0.050 0.735 0.130 1.065 ;
    END
END OAI31D4BWP

MACRO OAI32D0BWP
    CLASS CORE ;
    FOREIGN OAI32D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0790 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.985 0.710 1.055 ;
        RECT  0.130 0.345 0.540 0.415 ;
        RECT  0.240 0.890 0.310 1.055 ;
        RECT  0.105 0.890 0.240 0.960 ;
        RECT  0.105 0.185 0.130 0.415 ;
        RECT  0.035 0.185 0.105 0.960 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.900 0.545 1.015 0.615 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.635 0.665 0.905 ;
        RECT  0.550 0.635 0.595 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.800 -0.115 0.900 0.275 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.940 1.070 1.375 ;
        RECT  0.170 1.145 0.990 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.185 1.065 0.415 ;
        RECT  0.705 0.345 0.995 0.415 ;
        RECT  0.635 0.205 0.705 0.415 ;
        RECT  0.220 0.205 0.635 0.275 ;
    END
END OAI32D0BWP

MACRO OAI32D1BWP
    CLASS CORE ;
    FOREIGN OAI32D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1411 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.985 0.710 1.055 ;
        RECT  0.130 0.345 0.540 0.415 ;
        RECT  0.315 0.890 0.390 1.055 ;
        RECT  0.105 0.890 0.315 0.960 ;
        RECT  0.105 0.215 0.130 0.415 ;
        RECT  0.035 0.215 0.105 0.960 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.900 0.545 1.015 0.615 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.905 ;
        RECT  0.550 0.495 0.595 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.430 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.800 -0.115 0.900 0.275 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.845 1.070 1.375 ;
        RECT  0.170 1.145 0.990 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.255 1.065 0.415 ;
        RECT  0.705 0.345 0.995 0.415 ;
        RECT  0.635 0.205 0.705 0.415 ;
        RECT  0.220 0.205 0.635 0.275 ;
    END
END OAI32D1BWP

MACRO OAI32D2BWP
    CLASS CORE ;
    FOREIGN OAI32D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.845 1.670 1.055 ;
        RECT  1.230 0.985 1.550 1.055 ;
        RECT  1.160 0.345 1.230 1.055 ;
        RECT  0.210 0.345 1.160 0.415 ;
        RECT  1.155 0.775 1.160 1.055 ;
        RECT  0.570 0.985 1.155 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.775 ;
        RECT  1.370 0.705 1.855 0.775 ;
        RECT  1.300 0.520 1.370 0.775 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.495 0.945 0.765 ;
        RECT  0.385 0.695 0.845 0.765 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.090 0.640 ;
        RECT  1.015 0.495 1.085 0.905 ;
        RECT  0.245 0.835 1.015 0.905 ;
        RECT  0.175 0.495 0.245 0.905 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.860 -0.115 2.100 0.115 ;
        RECT  1.740 -0.115 1.860 0.135 ;
        RECT  1.440 -0.115 1.740 0.115 ;
        RECT  1.320 -0.115 1.440 0.135 ;
        RECT  0.000 -0.115 1.320 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.145 2.100 1.375 ;
        RECT  1.940 0.845 2.040 1.375 ;
        RECT  1.260 1.145 1.940 1.375 ;
        RECT  1.140 1.125 1.260 1.375 ;
        RECT  0.145 1.145 1.140 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 0.205 2.050 0.395 ;
        RECT  0.130 0.205 1.970 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OAI32D2BWP

MACRO OAI32D4BWP
    CLASS CORE ;
    FOREIGN OAI32D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.185 2.005 0.465 ;
        RECT  1.995 0.695 2.005 1.035 ;
        RECT  1.935 0.185 1.995 1.035 ;
        RECT  1.785 0.355 1.935 0.815 ;
        RECT  1.645 0.355 1.785 0.465 ;
        RECT  1.645 0.695 1.785 0.815 ;
        RECT  1.575 0.185 1.645 0.465 ;
        RECT  1.575 0.695 1.645 1.035 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.905 ;
        RECT  0.700 0.495 0.735 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.950 0.790 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.565 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.475 ;
        RECT  1.850 -0.115 2.110 0.115 ;
        RECT  1.730 -0.115 1.850 0.280 ;
        RECT  1.440 -0.115 1.730 0.115 ;
        RECT  1.360 -0.115 1.440 0.315 ;
        RECT  0.880 -0.115 1.360 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.675 2.190 1.375 ;
        RECT  1.850 1.145 2.110 1.375 ;
        RECT  1.730 0.885 1.850 1.375 ;
        RECT  1.440 1.145 1.730 1.375 ;
        RECT  1.360 0.845 1.440 1.375 ;
        RECT  1.070 1.145 1.360 1.375 ;
        RECT  0.950 1.125 1.070 1.375 ;
        RECT  0.140 1.145 0.950 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.355 1.715 0.465 ;
        RECT  1.645 0.695 1.715 0.815 ;
        RECT  1.575 0.185 1.645 0.465 ;
        RECT  1.575 0.695 1.645 1.035 ;
        RECT  1.495 0.545 1.670 0.615 ;
        RECT  1.425 0.395 1.495 0.775 ;
        RECT  1.230 0.395 1.425 0.465 ;
        RECT  1.230 0.705 1.425 0.775 ;
        RECT  1.090 0.545 1.320 0.615 ;
        RECT  1.160 0.185 1.230 0.465 ;
        RECT  1.160 0.705 1.230 1.035 ;
        RECT  1.020 0.345 1.090 1.055 ;
        RECT  0.210 0.205 1.070 0.275 ;
        RECT  0.130 0.345 1.020 0.415 ;
        RECT  0.570 0.985 1.020 1.055 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OAI32D4BWP

MACRO OAI32XD4BWP
    CLASS CORE ;
    FOREIGN OAI32XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.345 3.850 0.415 ;
        RECT  3.730 0.695 3.850 0.915 ;
        RECT  3.490 0.695 3.730 0.765 ;
        RECT  3.370 0.695 3.490 0.915 ;
        RECT  2.695 0.695 3.370 0.765 ;
        RECT  2.485 0.345 2.695 0.765 ;
        RECT  1.730 0.345 2.485 0.415 ;
        RECT  1.655 0.695 2.485 0.765 ;
        RECT  1.585 0.695 1.655 0.915 ;
        RECT  1.250 0.845 1.585 0.915 ;
        RECT  1.170 0.845 1.250 1.075 ;
        RECT  0.530 0.845 1.170 0.915 ;
        RECT  0.410 0.845 0.530 1.050 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.420 1.255 0.625 ;
        RECT  0.665 0.420 1.130 0.490 ;
        RECT  0.595 0.420 0.665 0.625 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.505 0.775 ;
        RECT  0.980 0.705 1.430 0.775 ;
        RECT  0.850 0.560 0.980 0.775 ;
        RECT  0.245 0.705 0.850 0.775 ;
        RECT  0.155 0.495 0.245 0.775 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.885 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 3.185 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 2.205 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 4.060 0.115 ;
        RECT  1.340 -0.115 1.460 0.210 ;
        RECT  1.090 -0.115 1.340 0.115 ;
        RECT  0.970 -0.115 1.090 0.210 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.210 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.210 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.145 4.060 1.375 ;
        RECT  2.290 0.995 2.370 1.375 ;
        RECT  2.030 1.145 2.290 1.375 ;
        RECT  1.910 1.000 2.030 1.375 ;
        RECT  1.620 1.145 1.910 1.375 ;
        RECT  1.540 0.985 1.620 1.375 ;
        RECT  0.880 1.145 1.540 1.375 ;
        RECT  0.800 0.985 0.880 1.375 ;
        RECT  0.130 1.145 0.800 1.375 ;
        RECT  0.050 0.855 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.345 3.850 0.415 ;
        RECT  3.730 0.695 3.850 0.915 ;
        RECT  3.490 0.695 3.730 0.765 ;
        RECT  3.370 0.695 3.490 0.915 ;
        RECT  2.765 0.695 3.370 0.765 ;
        RECT  1.730 0.345 2.415 0.415 ;
        RECT  1.655 0.695 2.415 0.765 ;
        RECT  1.585 0.695 1.655 0.915 ;
        RECT  1.250 0.845 1.585 0.915 ;
        RECT  1.170 0.845 1.250 1.075 ;
        RECT  0.530 0.845 1.170 0.915 ;
        RECT  0.410 0.845 0.530 1.050 ;
        RECT  3.930 0.205 4.010 0.375 ;
        RECT  3.930 0.755 4.010 1.065 ;
        RECT  1.640 0.205 3.930 0.275 ;
        RECT  3.660 0.995 3.930 1.065 ;
        RECT  3.560 0.845 3.660 1.070 ;
        RECT  3.300 0.995 3.560 1.065 ;
        RECT  3.200 0.845 3.300 1.065 ;
        RECT  2.470 0.995 3.200 1.065 ;
        RECT  2.185 0.845 3.130 0.915 ;
        RECT  2.115 0.845 2.185 1.075 ;
        RECT  1.810 0.845 2.115 0.915 ;
        RECT  1.730 0.845 1.810 0.985 ;
        RECT  1.560 0.205 1.640 0.350 ;
        RECT  0.130 0.280 1.560 0.350 ;
        RECT  0.050 0.230 0.130 0.350 ;
    END
END OAI32XD4BWP

MACRO OAI33D0BWP
    CLASS CORE ;
    FOREIGN OAI33D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0912 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.975 0.770 1.045 ;
        RECT  0.525 0.345 0.550 0.415 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.035 0.185 0.125 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.905 ;
        RECT  0.780 0.635 0.875 0.705 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.625 ;
        RECT  1.180 0.545 1.295 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.635 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.365 -0.115 1.400 0.115 ;
        RECT  1.255 -0.115 1.365 0.275 ;
        RECT  0.980 -0.115 1.255 0.115 ;
        RECT  0.860 -0.115 0.980 0.270 ;
        RECT  0.000 -0.115 0.860 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.270 0.920 1.350 1.375 ;
        RECT  0.130 1.145 1.270 1.375 ;
        RECT  0.050 0.920 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 0.195 1.160 0.410 ;
        RECT  0.735 0.340 1.080 0.410 ;
        RECT  0.665 0.195 0.735 0.410 ;
        RECT  0.220 0.195 0.665 0.265 ;
    END
END OAI33D0BWP

MACRO OAI33D1BWP
    CLASS CORE ;
    FOREIGN OAI33D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1657 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.975 0.760 1.045 ;
        RECT  0.525 0.345 0.550 0.415 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.905 ;
        RECT  0.805 0.495 0.875 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.625 ;
        RECT  1.180 0.545 1.295 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.365 -0.115 1.400 0.115 ;
        RECT  1.255 -0.115 1.365 0.275 ;
        RECT  0.980 -0.115 1.255 0.115 ;
        RECT  0.860 -0.115 0.980 0.270 ;
        RECT  0.000 -0.115 0.860 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.705 1.360 1.375 ;
        RECT  0.140 1.145 1.260 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.060 0.200 1.180 0.410 ;
        RECT  0.735 0.340 1.060 0.410 ;
        RECT  0.665 0.195 0.735 0.410 ;
        RECT  0.220 0.195 0.665 0.265 ;
    END
END OAI33D1BWP

MACRO OAI33D2BWP
    CLASS CORE ;
    FOREIGN OAI33D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2408 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.335 2.345 0.910 ;
        RECT  1.310 0.335 2.275 0.405 ;
        RECT  2.140 0.840 2.275 0.910 ;
        RECT  2.070 0.840 2.140 1.055 ;
        RECT  0.570 0.985 2.070 1.055 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.570 0.665 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 0.430 0.945 0.625 ;
        RECT  0.385 0.430 0.820 0.500 ;
        RECT  0.315 0.430 0.385 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.135 0.640 ;
        RECT  1.015 0.495 1.085 0.915 ;
        RECT  0.245 0.845 1.015 0.915 ;
        RECT  0.170 0.495 0.245 0.915 ;
        RECT  0.035 0.495 0.170 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0552 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.615 1.785 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.535 2.040 0.625 ;
        RECT  1.855 0.475 1.925 0.625 ;
        RECT  1.505 0.475 1.855 0.545 ;
        RECT  1.435 0.475 1.505 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.000 0.695 2.115 0.765 ;
        RECT  1.930 0.695 2.000 0.915 ;
        RECT  1.365 0.845 1.930 0.915 ;
        RECT  1.295 0.495 1.365 0.915 ;
        RECT  1.255 0.495 1.295 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.060 -0.115 2.380 0.115 ;
        RECT  0.940 -0.115 1.060 0.220 ;
        RECT  0.690 -0.115 0.940 0.115 ;
        RECT  0.570 -0.115 0.690 0.220 ;
        RECT  0.330 -0.115 0.570 0.115 ;
        RECT  0.210 -0.115 0.330 0.220 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.145 2.380 1.375 ;
        RECT  2.220 0.990 2.320 1.375 ;
        RECT  1.240 1.145 2.220 1.375 ;
        RECT  1.120 1.125 1.240 1.375 ;
        RECT  0.130 1.145 1.120 1.375 ;
        RECT  0.050 0.980 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.195 2.330 0.265 ;
        RECT  1.155 0.195 1.225 0.360 ;
        RECT  0.130 0.290 1.155 0.360 ;
        RECT  0.050 0.230 0.130 0.360 ;
    END
END OAI33D2BWP

MACRO OAI33D4BWP
    CLASS CORE ;
    FOREIGN OAI33D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.785 1.785 0.905 ;
        RECT  1.710 0.185 1.780 0.465 ;
        RECT  1.575 0.355 1.710 0.465 ;
        RECT  1.430 0.355 1.575 0.905 ;
        RECT  1.365 0.185 1.430 0.905 ;
        RECT  1.360 0.185 1.365 0.465 ;
        RECT  1.340 0.785 1.365 0.905 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.660 0.495 0.735 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.125 0.640 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.550 0.905 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.125 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.240 0.115 ;
        RECT  1.880 -0.115 2.000 0.280 ;
        RECT  1.630 -0.115 1.880 0.115 ;
        RECT  1.510 -0.115 1.630 0.275 ;
        RECT  1.260 -0.115 1.510 0.115 ;
        RECT  1.140 -0.115 1.260 0.135 ;
        RECT  0.880 -0.115 1.140 0.115 ;
        RECT  0.760 -0.115 0.880 0.135 ;
        RECT  0.000 -0.115 0.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.145 2.240 1.375 ;
        RECT  1.880 1.115 2.000 1.375 ;
        RECT  1.620 1.145 1.880 1.375 ;
        RECT  1.500 1.115 1.620 1.375 ;
        RECT  1.240 1.145 1.500 1.375 ;
        RECT  1.120 1.115 1.240 1.375 ;
        RECT  0.140 1.145 1.120 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.785 1.785 0.905 ;
        RECT  1.710 0.185 1.780 0.465 ;
        RECT  1.645 0.355 1.710 0.465 ;
        RECT  2.180 0.370 2.200 0.905 ;
        RECT  2.130 0.195 2.180 1.075 ;
        RECT  2.080 0.195 2.130 0.440 ;
        RECT  2.080 0.835 2.130 1.075 ;
        RECT  1.920 0.370 2.080 0.440 ;
        RECT  1.990 0.520 2.060 0.765 ;
        RECT  1.925 0.695 1.990 0.765 ;
        RECT  1.855 0.695 1.925 1.045 ;
        RECT  1.850 0.370 1.920 0.615 ;
        RECT  1.265 0.975 1.855 1.045 ;
        RECT  1.730 0.545 1.850 0.615 ;
        RECT  1.195 0.205 1.265 1.045 ;
        RECT  0.145 0.205 1.195 0.275 ;
        RECT  0.570 0.975 1.195 1.045 ;
        RECT  0.210 0.345 1.070 0.415 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OAI33D4BWP

MACRO OAI33XD4BWP
    CLASS CORE ;
    FOREIGN OAI33XD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.4900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.345 4.690 0.415 ;
        RECT  4.570 0.695 4.690 0.925 ;
        RECT  4.330 0.695 4.570 0.765 ;
        RECT  4.210 0.695 4.330 0.925 ;
        RECT  3.535 0.695 4.210 0.765 ;
        RECT  3.325 0.345 3.535 0.765 ;
        RECT  2.590 0.345 3.325 0.415 ;
        RECT  0.690 0.695 3.325 0.765 ;
        RECT  0.570 0.695 0.690 0.925 ;
        RECT  0.330 0.695 0.570 0.765 ;
        RECT  0.210 0.695 0.330 0.925 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.660 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.365 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.345 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.725 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.495 4.025 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 3.045 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.320 -0.115 4.900 0.115 ;
        RECT  2.240 -0.115 2.320 0.275 ;
        RECT  1.940 -0.115 2.240 0.115 ;
        RECT  1.860 -0.115 1.940 0.275 ;
        RECT  1.390 -0.115 1.860 0.115 ;
        RECT  1.310 -0.115 1.390 0.275 ;
        RECT  1.030 -0.115 1.310 0.115 ;
        RECT  0.950 -0.115 1.030 0.275 ;
        RECT  0.670 -0.115 0.950 0.115 ;
        RECT  0.590 -0.115 0.670 0.275 ;
        RECT  0.310 -0.115 0.590 0.115 ;
        RECT  0.230 -0.115 0.310 0.275 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.145 4.900 1.375 ;
        RECT  3.140 0.985 3.240 1.375 ;
        RECT  2.860 1.145 3.140 1.375 ;
        RECT  2.780 0.995 2.860 1.375 ;
        RECT  2.490 1.145 2.780 1.375 ;
        RECT  2.410 0.845 2.490 1.375 ;
        RECT  2.120 1.145 2.410 1.375 ;
        RECT  2.040 0.995 2.120 1.375 ;
        RECT  1.760 1.145 2.040 1.375 ;
        RECT  1.660 0.985 1.760 1.375 ;
        RECT  0.000 1.145 1.660 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.345 4.690 0.415 ;
        RECT  4.570 0.695 4.690 0.925 ;
        RECT  4.330 0.695 4.570 0.765 ;
        RECT  4.210 0.695 4.330 0.925 ;
        RECT  3.605 0.695 4.210 0.765 ;
        RECT  2.590 0.345 3.255 0.415 ;
        RECT  0.690 0.695 3.255 0.765 ;
        RECT  0.570 0.695 0.690 0.925 ;
        RECT  0.330 0.695 0.570 0.765 ;
        RECT  0.210 0.695 0.330 0.925 ;
        RECT  4.770 0.205 4.850 0.395 ;
        RECT  4.770 0.735 4.850 1.065 ;
        RECT  2.510 0.205 4.770 0.275 ;
        RECT  4.500 0.995 4.770 1.065 ;
        RECT  4.400 0.845 4.500 1.065 ;
        RECT  4.140 0.995 4.400 1.065 ;
        RECT  4.040 0.845 4.140 1.065 ;
        RECT  3.310 0.995 4.040 1.065 ;
        RECT  3.050 0.845 3.970 0.915 ;
        RECT  2.970 0.845 3.050 1.075 ;
        RECT  2.690 0.845 2.970 0.915 ;
        RECT  2.570 0.845 2.690 1.050 ;
        RECT  2.430 0.205 2.510 0.415 ;
        RECT  2.130 0.345 2.430 0.415 ;
        RECT  2.210 0.845 2.330 1.050 ;
        RECT  1.930 0.845 2.210 0.915 ;
        RECT  2.050 0.185 2.130 0.415 ;
        RECT  1.745 0.345 2.050 0.415 ;
        RECT  1.850 0.845 1.930 1.075 ;
        RECT  0.930 0.845 1.850 0.915 ;
        RECT  1.675 0.185 1.745 0.415 ;
        RECT  1.565 0.340 1.675 0.415 ;
        RECT  0.860 0.995 1.590 1.065 ;
        RECT  1.495 0.185 1.565 0.415 ;
        RECT  1.210 0.345 1.495 0.415 ;
        RECT  1.130 0.185 1.210 0.415 ;
        RECT  0.850 0.345 1.130 0.415 ;
        RECT  0.760 0.845 0.860 1.065 ;
        RECT  0.770 0.185 0.850 0.415 ;
        RECT  0.490 0.345 0.770 0.415 ;
        RECT  0.500 0.995 0.760 1.065 ;
        RECT  0.400 0.845 0.500 1.065 ;
        RECT  0.410 0.185 0.490 0.415 ;
        RECT  0.130 0.345 0.410 0.415 ;
        RECT  0.130 0.995 0.400 1.065 ;
        RECT  0.050 0.255 0.130 0.415 ;
        RECT  0.050 0.735 0.130 1.065 ;
    END
END OAI33XD4BWP

MACRO OD25DCAP16BWP
    CLASS CORE ;
    FOREIGN OD25DCAP16BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.115 2.240 0.115 ;
        RECT  1.740 -0.115 1.840 0.770 ;
        RECT  0.500 -0.115 1.740 0.115 ;
        RECT  0.400 -0.115 0.500 0.770 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.205 1.145 2.240 1.375 ;
        RECT  1.205 0.920 1.680 1.000 ;
        RECT  1.035 0.920 1.205 1.375 ;
        RECT  0.560 0.920 1.035 1.000 ;
        RECT  0.000 1.145 1.035 1.375 ;
        END
    END VDD
END OD25DCAP16BWP

MACRO OD25DCAP32BWP
    CLASS CORE ;
    FOREIGN OD25DCAP32BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.080 -0.115 4.480 0.115 ;
        RECT  3.980 -0.115 4.080 0.770 ;
        RECT  2.290 -0.115 3.980 0.115 ;
        RECT  2.190 -0.115 2.290 0.770 ;
        RECT  0.500 -0.115 2.190 0.115 ;
        RECT  0.400 -0.115 0.500 0.770 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.220 1.145 4.480 1.375 ;
        RECT  3.220 0.920 3.920 1.000 ;
        RECT  3.050 0.920 3.220 1.375 ;
        RECT  2.350 0.920 3.050 1.000 ;
        RECT  1.430 1.145 3.050 1.375 ;
        RECT  1.430 0.920 2.130 1.000 ;
        RECT  1.260 0.920 1.430 1.375 ;
        RECT  0.560 0.920 1.260 1.000 ;
        RECT  0.000 1.145 1.260 1.375 ;
        END
    END VDD
END OD25DCAP32BWP

MACRO OD25DCAP64BWP
    CLASS CORE ;
    FOREIGN OD25DCAP64BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.560 -0.115 8.960 0.115 ;
        RECT  8.460 -0.115 8.560 0.770 ;
        RECT  6.550 -0.115 8.460 0.115 ;
        RECT  6.440 -0.115 6.550 0.770 ;
        RECT  4.530 -0.115 6.440 0.115 ;
        RECT  4.430 -0.115 4.530 0.770 ;
        RECT  2.520 -0.115 4.430 0.115 ;
        RECT  2.410 -0.115 2.520 0.770 ;
        RECT  0.500 -0.115 2.410 0.115 ;
        RECT  0.400 -0.115 0.500 0.770 ;
        RECT  0.000 -0.115 0.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.585 1.145 8.960 1.375 ;
        RECT  7.585 0.910 8.400 0.990 ;
        RECT  7.415 0.910 7.585 1.375 ;
        RECT  6.605 0.910 7.415 0.990 ;
        RECT  5.570 1.145 7.415 1.375 ;
        RECT  5.570 0.910 6.385 0.990 ;
        RECT  5.400 0.910 5.570 1.375 ;
        RECT  4.590 0.910 5.400 0.990 ;
        RECT  3.555 1.145 5.400 1.375 ;
        RECT  3.555 0.910 4.370 0.990 ;
        RECT  3.385 0.910 3.555 1.375 ;
        RECT  2.575 0.910 3.385 0.990 ;
        RECT  1.540 1.145 3.385 1.375 ;
        RECT  1.540 0.910 2.355 0.990 ;
        RECT  1.370 0.910 1.540 1.375 ;
        RECT  0.560 0.910 1.370 0.990 ;
        RECT  0.000 1.145 1.370 1.375 ;
        END
    END VDD
END OD25DCAP64BWP

MACRO OR2D0BWP
    CLASS CORE ;
    FOREIGN OR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.185 0.805 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 -0.115 0.840 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.145 -0.115 0.480 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.000 1.145 0.480 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.565 0.345 0.635 0.915 ;
        RECT  0.340 0.345 0.565 0.415 ;
        RECT  0.130 0.845 0.565 0.915 ;
        RECT  0.260 0.185 0.340 0.415 ;
        RECT  0.050 0.845 0.130 1.050 ;
    END
END OR2D0BWP

MACRO OR2D1BWP
    CLASS CORE ;
    FOREIGN OR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.185 0.805 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 -0.115 0.840 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.145 -0.115 0.480 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.000 1.145 0.480 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.565 0.345 0.635 0.915 ;
        RECT  0.340 0.345 0.565 0.415 ;
        RECT  0.130 0.845 0.565 0.915 ;
        RECT  0.260 0.185 0.340 0.415 ;
        RECT  0.050 0.735 0.130 1.035 ;
    END
END OR2D1BWP

MACRO OR2D2BWP
    CLASS CORE ;
    FOREIGN OR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.745 0.355 0.805 0.905 ;
        RECT  0.735 0.185 0.745 1.035 ;
        RECT  0.675 0.185 0.735 0.465 ;
        RECT  0.675 0.740 0.735 1.035 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.115 0.980 0.115 ;
        RECT  0.835 -0.115 0.945 0.285 ;
        RECT  0.560 -0.115 0.835 0.115 ;
        RECT  0.440 -0.115 0.560 0.275 ;
        RECT  0.165 -0.115 0.440 0.115 ;
        RECT  0.055 -0.115 0.165 0.275 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.960 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.985 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.535 0.345 0.605 0.915 ;
        RECT  0.325 0.345 0.535 0.415 ;
        RECT  0.150 0.845 0.535 0.915 ;
        RECT  0.255 0.185 0.325 0.415 ;
        RECT  0.070 0.735 0.150 1.035 ;
    END
END OR2D2BWP

MACRO OR2D4BWP
    CLASS CORE ;
    FOREIGN OR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.445 0.465 ;
        RECT  1.435 0.695 1.445 1.035 ;
        RECT  1.375 0.185 1.435 1.035 ;
        RECT  1.225 0.355 1.375 0.815 ;
        RECT  1.085 0.355 1.225 0.465 ;
        RECT  1.085 0.695 1.225 0.815 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.695 1.085 1.035 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.520 0.740 0.640 ;
        RECT  0.595 0.520 0.665 0.905 ;
        RECT  0.245 0.835 0.595 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.115 1.680 0.115 ;
        RECT  1.550 -0.115 1.630 0.475 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.280 ;
        RECT  0.900 -0.115 1.170 0.115 ;
        RECT  0.780 -0.115 0.900 0.275 ;
        RECT  0.510 -0.115 0.780 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.390 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.145 1.680 1.375 ;
        RECT  1.550 0.675 1.630 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.885 1.290 1.375 ;
        RECT  0.900 1.145 1.170 1.375 ;
        RECT  0.780 1.115 0.900 1.375 ;
        RECT  0.140 1.145 0.780 1.375 ;
        RECT  0.040 0.975 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.355 1.155 0.465 ;
        RECT  1.085 0.695 1.155 0.815 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.695 1.085 1.035 ;
        RECT  0.935 0.545 1.130 0.615 ;
        RECT  0.865 0.345 0.935 1.045 ;
        RECT  0.665 0.345 0.865 0.415 ;
        RECT  0.390 0.975 0.865 1.045 ;
        RECT  0.595 0.185 0.665 0.415 ;
        RECT  0.305 0.345 0.595 0.415 ;
        RECT  0.235 0.185 0.305 0.415 ;
    END
END OR2D4BWP

MACRO OR2D8BWP
    CLASS CORE ;
    FOREIGN OR2D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.185 2.570 0.470 ;
        RECT  2.490 0.695 2.570 1.035 ;
        RECT  2.190 0.340 2.490 0.470 ;
        RECT  2.190 0.695 2.490 0.815 ;
        RECT  2.135 0.185 2.190 0.470 ;
        RECT  2.135 0.695 2.190 1.045 ;
        RECT  2.110 0.185 2.135 1.045 ;
        RECT  1.925 0.340 2.110 0.815 ;
        RECT  1.810 0.340 1.925 0.465 ;
        RECT  1.810 0.695 1.925 0.815 ;
        RECT  1.730 0.185 1.810 0.465 ;
        RECT  1.730 0.695 1.810 1.035 ;
        RECT  1.430 0.340 1.730 0.465 ;
        RECT  1.430 0.695 1.730 0.815 ;
        RECT  1.350 0.185 1.430 0.465 ;
        RECT  1.350 0.695 1.430 1.035 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.135 0.640 ;
        RECT  1.010 0.495 1.085 0.770 ;
        RECT  0.525 0.700 1.010 0.770 ;
        RECT  0.435 0.495 0.525 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.545 0.875 0.625 ;
        RECT  0.730 0.345 0.805 0.625 ;
        RECT  0.325 0.345 0.730 0.415 ;
        RECT  0.250 0.345 0.325 0.620 ;
        RECT  0.140 0.540 0.250 0.620 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.465 ;
        RECT  2.400 -0.115 2.670 0.115 ;
        RECT  2.280 -0.115 2.400 0.270 ;
        RECT  2.020 -0.115 2.280 0.115 ;
        RECT  1.900 -0.115 2.020 0.270 ;
        RECT  1.640 -0.115 1.900 0.115 ;
        RECT  1.520 -0.115 1.640 0.270 ;
        RECT  1.250 -0.115 1.520 0.115 ;
        RECT  1.170 -0.115 1.250 0.280 ;
        RECT  0.900 -0.115 1.170 0.115 ;
        RECT  0.780 -0.115 0.900 0.135 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.135 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.675 2.750 1.375 ;
        RECT  2.400 1.145 2.670 1.375 ;
        RECT  2.280 0.885 2.400 1.375 ;
        RECT  2.020 1.145 2.280 1.375 ;
        RECT  1.900 0.885 2.020 1.375 ;
        RECT  1.640 1.145 1.900 1.375 ;
        RECT  1.520 0.885 1.640 1.375 ;
        RECT  1.250 1.145 1.520 1.375 ;
        RECT  1.150 0.980 1.250 1.375 ;
        RECT  0.510 1.145 1.150 1.375 ;
        RECT  0.410 0.980 0.510 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.185 2.570 0.470 ;
        RECT  2.490 0.695 2.570 1.035 ;
        RECT  2.205 0.340 2.490 0.470 ;
        RECT  2.205 0.695 2.490 0.815 ;
        RECT  1.810 0.340 1.855 0.465 ;
        RECT  1.810 0.695 1.855 0.815 ;
        RECT  1.730 0.185 1.810 0.465 ;
        RECT  1.730 0.695 1.810 1.035 ;
        RECT  1.430 0.340 1.730 0.465 ;
        RECT  1.430 0.695 1.730 0.815 ;
        RECT  1.350 0.185 1.430 0.465 ;
        RECT  1.090 0.350 1.210 0.420 ;
        RECT  0.870 0.840 1.210 0.910 ;
        RECT  1.010 0.205 1.090 0.420 ;
        RECT  0.210 0.205 1.010 0.275 ;
        RECT  0.790 0.840 0.870 1.075 ;
        RECT  0.125 0.840 0.790 0.910 ;
        RECT  0.055 0.735 0.125 1.035 ;
        RECT  1.350 0.695 1.430 1.035 ;
        RECT  2.275 0.545 2.615 0.615 ;
        RECT  1.280 0.545 1.745 0.615 ;
        RECT  1.210 0.350 1.280 0.910 ;
    END
END OR2D8BWP

MACRO OR2XD1BWP
    CLASS CORE ;
    FOREIGN OR2XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.185 0.805 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.400 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.540 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 -0.115 0.840 0.115 ;
        RECT  0.480 -0.115 0.600 0.275 ;
        RECT  0.145 -0.115 0.480 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.985 0.600 1.375 ;
        RECT  0.000 1.145 0.480 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.565 0.355 0.635 0.915 ;
        RECT  0.350 0.355 0.565 0.425 ;
        RECT  0.130 0.845 0.565 0.915 ;
        RECT  0.240 0.185 0.350 0.425 ;
        RECT  0.050 0.735 0.130 1.035 ;
    END
END OR2XD1BWP

MACRO OR3D0BWP
    CLASS CORE ;
    FOREIGN OR3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.070 ;
        RECT  0.840 0.190 0.875 0.290 ;
        RECT  0.840 0.970 0.875 1.070 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.285 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 0.985 0.740 1.375 ;
        RECT  0.000 1.145 0.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.905 ;
        RECT  0.545 0.355 0.735 0.425 ;
        RECT  0.150 0.835 0.735 0.905 ;
        RECT  0.475 0.215 0.545 0.425 ;
        RECT  0.145 0.215 0.475 0.285 ;
        RECT  0.070 0.835 0.150 1.065 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OR3D0BWP

MACRO OR3D1BWP
    CLASS CORE ;
    FOREIGN OR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.075 ;
        RECT  0.840 0.190 0.875 0.290 ;
        RECT  0.835 0.975 0.875 1.075 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.285 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 0.975 0.740 1.375 ;
        RECT  0.000 1.145 0.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.905 ;
        RECT  0.545 0.355 0.735 0.425 ;
        RECT  0.160 0.835 0.735 0.905 ;
        RECT  0.475 0.215 0.545 0.425 ;
        RECT  0.145 0.215 0.475 0.285 ;
        RECT  0.060 0.835 0.160 1.075 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OR3D1BWP

MACRO OR3D2BWP
    CLASS CORE ;
    FOREIGN OR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.885 0.355 0.945 0.905 ;
        RECT  0.875 0.185 0.885 1.035 ;
        RECT  0.815 0.185 0.875 0.465 ;
        RECT  0.815 0.735 0.875 1.035 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.575 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 -0.115 1.120 0.115 ;
        RECT  0.990 -0.115 1.070 0.300 ;
        RECT  0.720 -0.115 0.990 0.115 ;
        RECT  0.600 -0.115 0.720 0.275 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.120 1.375 ;
        RECT  0.990 0.960 1.070 1.375 ;
        RECT  0.720 1.145 0.990 1.375 ;
        RECT  0.600 0.985 0.720 1.375 ;
        RECT  0.000 1.145 0.600 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.745 0.545 0.795 0.615 ;
        RECT  0.675 0.345 0.745 0.915 ;
        RECT  0.530 0.345 0.675 0.415 ;
        RECT  0.170 0.845 0.675 0.915 ;
        RECT  0.460 0.215 0.530 0.415 ;
        RECT  0.145 0.215 0.460 0.285 ;
        RECT  0.050 0.845 0.170 1.060 ;
        RECT  0.035 0.185 0.145 0.285 ;
    END
END OR3D2BWP

MACRO OR3D4BWP
    CLASS CORE ;
    FOREIGN OR3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.865 0.465 ;
        RECT  1.855 0.695 1.865 1.035 ;
        RECT  1.795 0.185 1.855 1.035 ;
        RECT  1.645 0.355 1.795 0.815 ;
        RECT  1.485 0.355 1.645 0.465 ;
        RECT  1.485 0.695 1.645 0.815 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.695 1.485 1.035 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.355 0.685 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.965 0.775 ;
        RECT  0.385 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.385 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0452 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.495 1.135 0.915 ;
        RECT  0.245 0.845 1.055 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.475 ;
        RECT  1.700 -0.115 1.970 0.115 ;
        RECT  1.580 -0.115 1.700 0.280 ;
        RECT  1.300 -0.115 1.580 0.115 ;
        RECT  1.180 -0.115 1.300 0.145 ;
        RECT  0.900 -0.115 1.180 0.115 ;
        RECT  0.780 -0.115 0.900 0.145 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.145 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.675 2.050 1.375 ;
        RECT  1.700 1.145 1.970 1.375 ;
        RECT  1.580 0.885 1.700 1.375 ;
        RECT  1.300 1.145 1.580 1.375 ;
        RECT  1.180 1.125 1.300 1.375 ;
        RECT  0.145 1.145 1.180 1.375 ;
        RECT  0.035 0.980 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.485 0.355 1.575 0.465 ;
        RECT  1.485 0.695 1.575 0.815 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.695 1.485 1.035 ;
        RECT  1.335 0.545 1.530 0.615 ;
        RECT  1.265 0.215 1.335 1.055 ;
        RECT  0.210 0.215 1.265 0.285 ;
        RECT  0.570 0.985 1.265 1.055 ;
    END
END OR3D4BWP

MACRO OR3D8BWP
    CLASS CORE ;
    FOREIGN OR3D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 0.185 3.130 0.470 ;
        RECT  3.050 0.695 3.130 1.035 ;
        RECT  2.750 0.340 3.050 0.470 ;
        RECT  2.750 0.695 3.050 0.815 ;
        RECT  2.695 0.185 2.750 0.470 ;
        RECT  2.695 0.695 2.750 1.045 ;
        RECT  2.670 0.185 2.695 1.045 ;
        RECT  2.485 0.340 2.670 0.815 ;
        RECT  2.370 0.340 2.485 0.465 ;
        RECT  2.370 0.695 2.485 0.815 ;
        RECT  2.290 0.185 2.370 0.465 ;
        RECT  2.290 0.695 2.370 1.035 ;
        RECT  1.990 0.340 2.290 0.465 ;
        RECT  1.990 0.695 2.290 0.815 ;
        RECT  1.910 0.185 1.990 0.465 ;
        RECT  1.910 0.695 1.990 1.035 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.645 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.085 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0678 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.525 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.465 ;
        RECT  2.960 -0.115 3.230 0.115 ;
        RECT  2.840 -0.115 2.960 0.270 ;
        RECT  2.580 -0.115 2.840 0.115 ;
        RECT  2.460 -0.115 2.580 0.270 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.270 ;
        RECT  1.800 -0.115 2.080 0.115 ;
        RECT  1.680 -0.115 1.800 0.275 ;
        RECT  1.410 -0.115 1.680 0.115 ;
        RECT  1.290 -0.115 1.410 0.275 ;
        RECT  1.050 -0.115 1.290 0.115 ;
        RECT  0.930 -0.115 1.050 0.275 ;
        RECT  0.690 -0.115 0.930 0.115 ;
        RECT  0.570 -0.115 0.690 0.275 ;
        RECT  0.330 -0.115 0.570 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 1.145 3.360 1.375 ;
        RECT  3.230 0.675 3.310 1.375 ;
        RECT  2.960 1.145 3.230 1.375 ;
        RECT  2.840 0.885 2.960 1.375 ;
        RECT  2.580 1.145 2.840 1.375 ;
        RECT  2.460 0.885 2.580 1.375 ;
        RECT  2.200 1.145 2.460 1.375 ;
        RECT  2.080 0.885 2.200 1.375 ;
        RECT  1.780 1.145 2.080 1.375 ;
        RECT  1.700 0.735 1.780 1.375 ;
        RECT  1.400 1.145 1.700 1.375 ;
        RECT  1.300 0.845 1.400 1.375 ;
        RECT  0.000 1.145 1.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.050 0.185 3.130 0.470 ;
        RECT  3.050 0.695 3.130 1.035 ;
        RECT  2.765 0.340 3.050 0.470 ;
        RECT  2.765 0.695 3.050 0.815 ;
        RECT  2.370 0.340 2.415 0.465 ;
        RECT  2.370 0.695 2.415 0.815 ;
        RECT  2.290 0.185 2.370 0.465 ;
        RECT  2.290 0.695 2.370 1.035 ;
        RECT  1.990 0.340 2.290 0.465 ;
        RECT  1.990 0.695 2.290 0.815 ;
        RECT  1.910 0.185 1.990 0.465 ;
        RECT  1.910 0.695 1.990 1.035 ;
        RECT  2.835 0.545 3.175 0.615 ;
        RECT  1.800 0.545 2.310 0.615 ;
        RECT  1.730 0.345 1.800 0.615 ;
        RECT  1.570 0.345 1.730 0.415 ;
        RECT  1.490 0.185 1.570 0.415 ;
        RECT  1.495 0.705 1.565 1.035 ;
        RECT  1.205 0.705 1.495 0.775 ;
        RECT  1.210 0.345 1.490 0.415 ;
        RECT  1.130 0.185 1.210 0.415 ;
        RECT  1.135 0.705 1.205 1.035 ;
        RECT  0.870 0.705 1.135 0.775 ;
        RECT  0.850 0.345 1.130 0.415 ;
        RECT  0.680 0.995 1.050 1.065 ;
        RECT  0.750 0.705 0.870 0.925 ;
        RECT  0.770 0.185 0.850 0.415 ;
        RECT  0.665 0.345 0.770 0.415 ;
        RECT  0.580 0.845 0.680 1.065 ;
        RECT  0.595 0.345 0.665 0.775 ;
        RECT  0.490 0.345 0.595 0.415 ;
        RECT  0.510 0.705 0.595 0.775 ;
        RECT  0.210 0.995 0.580 1.065 ;
        RECT  0.390 0.705 0.510 0.925 ;
        RECT  0.410 0.185 0.490 0.415 ;
        RECT  0.125 0.345 0.410 0.415 ;
        RECT  0.125 0.705 0.390 0.775 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.705 0.125 1.035 ;
    END
END OR3D8BWP

MACRO OR3XD1BWP
    CLASS CORE ;
    FOREIGN OR3XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.075 ;
        RECT  0.840 0.190 0.875 0.290 ;
        RECT  0.835 0.975 0.875 1.075 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.545 0.240 0.615 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 0.980 0.115 ;
        RECT  0.620 -0.115 0.740 0.285 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.220 -0.115 0.340 0.145 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 0.975 0.740 1.375 ;
        RECT  0.000 1.145 0.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.905 ;
        RECT  0.545 0.355 0.735 0.425 ;
        RECT  0.160 0.835 0.735 0.905 ;
        RECT  0.475 0.215 0.545 0.425 ;
        RECT  0.130 0.215 0.475 0.285 ;
        RECT  0.060 0.835 0.160 1.075 ;
        RECT  0.050 0.215 0.130 0.395 ;
    END
END OR3XD1BWP

MACRO OR4D0BWP
    CLASS CORE ;
    FOREIGN OR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0437 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.085 1.060 ;
        RECT  0.995 0.185 1.015 0.305 ;
        RECT  0.995 0.920 1.015 1.060 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.565 0.600 0.635 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.355 0.755 0.905 ;
        RECT  0.595 0.355 0.685 0.485 ;
        RECT  0.595 0.775 0.685 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.140 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.140 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 1.125 0.880 1.375 ;
        RECT  0.000 1.145 0.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.915 0.520 0.945 0.640 ;
        RECT  0.845 0.210 0.915 1.055 ;
        RECT  0.210 0.210 0.845 0.280 ;
        RECT  0.130 0.985 0.845 1.055 ;
        RECT  0.050 0.920 0.130 1.055 ;
    END
END OR4D0BWP

MACRO OR4D1BWP
    CLASS CORE ;
    FOREIGN OR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0874 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.085 1.060 ;
        RECT  0.995 0.185 1.015 0.305 ;
        RECT  0.995 0.920 1.015 1.060 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.600 0.565 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.520 0.755 0.705 ;
        RECT  0.665 0.635 0.685 0.705 ;
        RECT  0.595 0.635 0.665 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.140 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.140 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 1.125 0.880 1.375 ;
        RECT  0.000 1.145 0.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.915 0.520 0.945 0.640 ;
        RECT  0.845 0.210 0.915 1.055 ;
        RECT  0.210 0.210 0.845 0.280 ;
        RECT  0.130 0.985 0.845 1.055 ;
        RECT  0.050 0.845 0.130 1.055 ;
    END
END OR4D1BWP

MACRO OR4D2BWP
    CLASS CORE ;
    FOREIGN OR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.905 ;
        RECT  1.145 0.355 1.155 0.465 ;
        RECT  1.145 0.735 1.155 0.905 ;
        RECT  1.075 0.185 1.145 0.465 ;
        RECT  1.075 0.735 1.145 1.035 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.220 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.905 ;
        RECT  0.555 0.495 0.595 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0226 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.230 -0.115 1.350 0.275 ;
        RECT  0.960 -0.115 1.230 0.115 ;
        RECT  0.840 -0.115 0.960 0.275 ;
        RECT  0.540 -0.115 0.840 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.145 -0.115 0.420 0.115 ;
        RECT  0.035 -0.115 0.145 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.230 0.975 1.350 1.375 ;
        RECT  0.960 1.145 1.230 1.375 ;
        RECT  0.840 1.125 0.960 1.375 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.545 1.030 0.615 ;
        RECT  0.875 0.345 0.955 1.055 ;
        RECT  0.720 0.345 0.875 0.415 ;
        RECT  0.130 0.985 0.875 1.055 ;
        RECT  0.640 0.185 0.720 0.415 ;
        RECT  0.320 0.345 0.640 0.415 ;
        RECT  0.240 0.185 0.320 0.415 ;
        RECT  0.050 0.735 0.130 1.055 ;
    END
END OR4D2BWP

MACRO OR4D4BWP
    CLASS CORE ;
    FOREIGN OR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.195 0.185 2.275 1.035 ;
        RECT  2.065 0.355 2.195 0.815 ;
        RECT  1.905 0.355 2.065 0.465 ;
        RECT  1.905 0.695 2.065 0.815 ;
        RECT  1.835 0.185 1.905 0.465 ;
        RECT  1.835 0.695 1.905 1.035 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.225 0.775 ;
        RECT  0.665 0.705 1.130 0.775 ;
        RECT  0.575 0.495 0.665 0.775 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.545 1.460 0.625 ;
        RECT  1.295 0.345 1.365 0.625 ;
        RECT  0.405 0.345 1.295 0.415 ;
        RECT  0.315 0.345 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.510 1.615 0.915 ;
        RECT  0.245 0.845 1.545 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 -0.115 2.520 0.115 ;
        RECT  2.370 -0.115 2.450 0.475 ;
        RECT  2.110 -0.115 2.370 0.115 ;
        RECT  1.990 -0.115 2.110 0.280 ;
        RECT  1.740 -0.115 1.990 0.115 ;
        RECT  1.620 -0.115 1.740 0.135 ;
        RECT  1.340 -0.115 1.620 0.115 ;
        RECT  1.220 -0.115 1.340 0.135 ;
        RECT  0.940 -0.115 1.220 0.115 ;
        RECT  0.820 -0.115 0.940 0.135 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.145 2.520 1.375 ;
        RECT  2.370 0.675 2.450 1.375 ;
        RECT  2.110 1.145 2.370 1.375 ;
        RECT  1.990 0.885 2.110 1.375 ;
        RECT  1.740 1.145 1.990 1.375 ;
        RECT  1.620 1.125 1.740 1.375 ;
        RECT  0.145 1.145 1.620 1.375 ;
        RECT  0.035 0.985 0.145 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.905 0.355 1.995 0.465 ;
        RECT  1.905 0.695 1.995 0.815 ;
        RECT  1.835 0.185 1.905 0.465 ;
        RECT  1.835 0.695 1.905 1.035 ;
        RECT  1.755 0.545 1.980 0.615 ;
        RECT  1.685 0.205 1.755 1.055 ;
        RECT  1.515 0.205 1.685 0.275 ;
        RECT  0.810 0.985 1.685 1.055 ;
        RECT  1.445 0.205 1.515 0.440 ;
        RECT  0.210 0.205 1.445 0.275 ;
    END
END OR4D4BWP

MACRO OR4D8BWP
    CLASS CORE ;
    FOREIGN OR4D8BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.4032 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.475 0.695 3.545 1.035 ;
        RECT  3.185 0.365 3.475 0.465 ;
        RECT  3.185 0.695 3.475 0.815 ;
        RECT  3.115 0.185 3.185 0.465 ;
        RECT  3.115 0.695 3.185 1.035 ;
        RECT  2.905 0.365 3.115 0.815 ;
        RECT  2.825 0.365 2.905 0.465 ;
        RECT  2.825 0.695 2.905 0.815 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.755 0.695 2.825 1.035 ;
        RECT  2.465 0.365 2.755 0.465 ;
        RECT  2.465 0.695 2.755 0.815 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.395 0.695 2.465 1.035 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 2.100 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.645 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.085 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.525 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.465 ;
        RECT  3.370 -0.115 3.650 0.115 ;
        RECT  3.290 -0.115 3.370 0.285 ;
        RECT  3.010 -0.115 3.290 0.115 ;
        RECT  2.930 -0.115 3.010 0.285 ;
        RECT  2.650 -0.115 2.930 0.115 ;
        RECT  2.570 -0.115 2.650 0.285 ;
        RECT  2.310 -0.115 2.570 0.115 ;
        RECT  2.190 -0.115 2.310 0.275 ;
        RECT  1.950 -0.115 2.190 0.115 ;
        RECT  1.830 -0.115 1.950 0.275 ;
        RECT  1.590 -0.115 1.830 0.115 ;
        RECT  1.470 -0.115 1.590 0.275 ;
        RECT  1.230 -0.115 1.470 0.115 ;
        RECT  1.110 -0.115 1.230 0.275 ;
        RECT  0.870 -0.115 1.110 0.115 ;
        RECT  0.750 -0.115 0.870 0.275 ;
        RECT  0.510 -0.115 0.750 0.115 ;
        RECT  0.390 -0.115 0.510 0.275 ;
        RECT  0.140 -0.115 0.390 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.685 3.730 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 0.885 3.390 1.375 ;
        RECT  3.030 1.145 3.270 1.375 ;
        RECT  2.910 0.885 3.030 1.375 ;
        RECT  2.670 1.145 2.910 1.375 ;
        RECT  2.550 0.885 2.670 1.375 ;
        RECT  2.290 1.145 2.550 1.375 ;
        RECT  2.210 0.735 2.290 1.375 ;
        RECT  1.930 1.145 2.210 1.375 ;
        RECT  1.850 0.860 1.930 1.375 ;
        RECT  0.000 1.145 1.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.475 0.185 3.545 0.465 ;
        RECT  3.475 0.695 3.545 1.035 ;
        RECT  3.185 0.365 3.475 0.465 ;
        RECT  3.185 0.695 3.475 0.815 ;
        RECT  2.825 0.365 2.835 0.465 ;
        RECT  2.825 0.695 2.835 0.815 ;
        RECT  2.755 0.185 2.825 0.465 ;
        RECT  2.755 0.695 2.825 1.035 ;
        RECT  2.465 0.365 2.755 0.465 ;
        RECT  2.465 0.695 2.755 0.815 ;
        RECT  2.395 0.185 2.465 0.465 ;
        RECT  2.395 0.695 2.465 1.035 ;
        RECT  3.280 0.545 3.610 0.615 ;
        RECT  2.290 0.545 2.815 0.615 ;
        RECT  2.210 0.345 2.290 0.615 ;
        RECT  2.105 0.345 2.210 0.415 ;
        RECT  2.030 0.720 2.110 1.035 ;
        RECT  2.035 0.255 2.105 0.415 ;
        RECT  1.745 0.345 2.035 0.415 ;
        RECT  1.745 0.720 2.030 0.790 ;
        RECT  1.675 0.255 1.745 0.415 ;
        RECT  1.675 0.720 1.745 1.065 ;
        RECT  1.385 0.345 1.675 0.415 ;
        RECT  1.410 0.995 1.675 1.065 ;
        RECT  1.210 0.720 1.590 0.790 ;
        RECT  1.290 0.860 1.410 1.065 ;
        RECT  1.315 0.255 1.385 0.415 ;
        RECT  1.025 0.345 1.315 0.415 ;
        RECT  1.130 0.720 1.210 1.035 ;
        RECT  0.750 0.720 1.130 0.790 ;
        RECT  0.930 0.860 1.050 1.065 ;
        RECT  0.955 0.255 1.025 0.415 ;
        RECT  0.665 0.345 0.955 0.415 ;
        RECT  0.690 0.995 0.930 1.065 ;
        RECT  0.570 0.855 0.690 1.065 ;
        RECT  0.595 0.255 0.665 0.785 ;
        RECT  0.305 0.345 0.595 0.415 ;
        RECT  0.125 0.715 0.595 0.785 ;
        RECT  0.330 0.995 0.570 1.065 ;
        RECT  0.210 0.855 0.330 1.065 ;
        RECT  0.235 0.255 0.305 0.415 ;
        RECT  0.055 0.715 0.125 1.035 ;
    END
END OR4D8BWP

MACRO OR4XD1BWP
    CLASS CORE ;
    FOREIGN OR4XD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0874 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.085 1.045 ;
        RECT  0.995 0.185 1.015 0.465 ;
        RECT  0.995 0.735 1.015 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.520 0.755 0.905 ;
        RECT  0.595 0.775 0.685 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.900 -0.115 1.120 0.115 ;
        RECT  0.780 -0.115 0.900 0.145 ;
        RECT  0.520 -0.115 0.780 0.115 ;
        RECT  0.400 -0.115 0.520 0.145 ;
        RECT  0.130 -0.115 0.400 0.115 ;
        RECT  0.050 -0.115 0.130 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.145 1.120 1.375 ;
        RECT  0.760 1.125 0.880 1.375 ;
        RECT  0.000 1.145 0.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.915 0.520 0.945 0.640 ;
        RECT  0.845 0.215 0.915 1.055 ;
        RECT  0.710 0.215 0.845 0.285 ;
        RECT  0.130 0.985 0.845 1.055 ;
        RECT  0.590 0.215 0.710 0.425 ;
        RECT  0.210 0.215 0.590 0.285 ;
        RECT  0.050 0.845 0.130 1.055 ;
    END
END OR4XD1BWP

MACRO SDFCND0BWP
    CLASS CORE ;
    FOREIGN SDFCND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.215 4.585 0.905 ;
        RECT  4.495 0.215 4.515 0.335 ;
        RECT  4.500 0.775 4.515 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 0.715 4.220 0.785 ;
        RECT  4.090 0.215 4.185 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0330 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.355 3.745 0.640 ;
        RECT  3.605 0.520 3.665 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 -0.115 4.620 0.115 ;
        RECT  4.300 -0.115 4.380 0.335 ;
        RECT  3.535 -0.115 4.300 0.115 ;
        RECT  3.465 -0.115 3.535 0.440 ;
        RECT  2.550 -0.115 3.465 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 1.145 4.620 1.375 ;
        RECT  4.260 1.130 4.380 1.375 ;
        RECT  2.660 1.145 4.260 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.650 ;
        RECT  4.355 0.520 4.425 0.925 ;
        RECT  3.360 0.855 4.355 0.925 ;
        RECT  3.945 0.520 4.020 0.640 ;
        RECT  3.875 0.190 3.945 0.785 ;
        RECT  3.500 0.715 3.875 0.785 ;
        RECT  3.740 0.995 3.860 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.785 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.255 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.685 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.760 ;
        RECT  2.260 0.690 2.760 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.030 0.840 2.240 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.490 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFCND0BWP

MACRO SDFCND1BWP
    CLASS CORE ;
    FOREIGN SDFCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0803 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.190 4.585 1.065 ;
        RECT  4.495 0.190 4.515 0.470 ;
        RECT  4.500 0.775 4.515 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0803 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 0.715 4.220 0.785 ;
        RECT  4.090 0.190 4.185 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0330 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.355 3.745 0.640 ;
        RECT  3.605 0.520 3.665 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.375 -0.115 4.620 0.115 ;
        RECT  4.305 -0.115 4.375 0.330 ;
        RECT  3.535 -0.115 4.305 0.115 ;
        RECT  3.465 -0.115 3.535 0.440 ;
        RECT  2.550 -0.115 3.465 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 1.005 4.400 1.375 ;
        RECT  4.020 1.145 4.280 1.375 ;
        RECT  3.900 1.135 4.020 1.375 ;
        RECT  3.620 1.145 3.900 1.375 ;
        RECT  3.500 1.135 3.620 1.375 ;
        RECT  2.660 1.145 3.500 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.430 0.520 4.440 0.640 ;
        RECT  4.360 0.520 4.430 0.925 ;
        RECT  3.360 0.855 4.360 0.925 ;
        RECT  3.945 0.520 4.020 0.640 ;
        RECT  3.875 0.190 3.945 0.785 ;
        RECT  3.500 0.715 3.875 0.785 ;
        RECT  3.740 0.995 3.860 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.785 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.255 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.690 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.760 ;
        RECT  2.260 0.690 2.760 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.015 0.840 2.240 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCND1BWP

MACRO SDFCND2BWP
    CLASS CORE ;
    FOREIGN SDFCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.355 5.005 0.805 ;
        RECT  4.935 0.185 4.945 1.035 ;
        RECT  4.875 0.185 4.935 0.465 ;
        RECT  4.875 0.735 4.935 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.590 0.780 ;
        RECT  4.495 0.185 4.515 0.485 ;
        RECT  4.470 0.710 4.515 0.780 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.580 0.535 3.675 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.300 ;
        RECT  4.755 -0.115 5.050 0.115 ;
        RECT  4.685 -0.115 4.755 0.465 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.275 ;
        RECT  3.555 -0.115 4.280 0.115 ;
        RECT  3.485 -0.115 3.555 0.400 ;
        RECT  2.550 -0.115 3.485 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.055 0.895 5.125 1.375 ;
        RECT  4.780 1.145 5.055 1.375 ;
        RECT  4.660 0.995 4.780 1.375 ;
        RECT  4.410 1.145 4.660 1.375 ;
        RECT  4.290 0.995 4.410 1.375 ;
        RECT  2.660 1.145 4.290 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.805 0.545 4.860 0.615 ;
        RECT  4.735 0.545 4.805 0.925 ;
        RECT  3.360 0.855 4.735 0.925 ;
        RECT  4.375 0.520 4.430 0.640 ;
        RECT  4.305 0.350 4.375 0.780 ;
        RECT  3.840 0.350 4.305 0.420 ;
        RECT  3.500 0.710 4.305 0.780 ;
        RECT  3.740 0.995 3.860 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.780 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.235 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.690 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.760 ;
        RECT  2.260 0.690 2.760 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.030 0.840 2.240 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCND2BWP

MACRO SDFCND4BWP
    CLASS CORE ;
    FOREIGN SDFCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.185 5.925 0.465 ;
        RECT  5.915 0.775 5.925 1.065 ;
        RECT  5.855 0.185 5.915 1.065 ;
        RECT  5.705 0.355 5.855 0.905 ;
        RECT  5.565 0.355 5.705 0.465 ;
        RECT  5.565 0.775 5.705 0.905 ;
        RECT  5.495 0.185 5.565 0.465 ;
        RECT  5.495 0.775 5.565 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.705 5.230 0.795 ;
        RECT  5.135 0.185 5.205 0.485 ;
        RECT  5.075 0.355 5.135 0.485 ;
        RECT  4.865 0.355 5.075 0.795 ;
        RECT  4.845 0.355 4.865 0.485 ;
        RECT  4.750 0.705 4.865 0.795 ;
        RECT  4.775 0.185 4.845 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.535 0.495 3.675 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 -0.115 6.160 0.115 ;
        RECT  6.035 -0.115 6.105 0.465 ;
        RECT  5.770 -0.115 6.035 0.115 ;
        RECT  5.650 -0.115 5.770 0.275 ;
        RECT  5.385 -0.115 5.650 0.115 ;
        RECT  5.315 -0.115 5.385 0.465 ;
        RECT  5.050 -0.115 5.315 0.115 ;
        RECT  4.930 -0.115 5.050 0.275 ;
        RECT  4.665 -0.115 4.930 0.115 ;
        RECT  4.595 -0.115 4.665 0.310 ;
        RECT  4.340 -0.115 4.595 0.115 ;
        RECT  4.220 -0.115 4.340 0.145 ;
        RECT  3.325 -0.115 4.220 0.115 ;
        RECT  3.255 -0.115 3.325 0.250 ;
        RECT  2.570 -0.115 3.255 0.115 ;
        RECT  2.500 -0.115 2.570 0.290 ;
        RECT  1.480 -0.115 2.500 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 1.145 6.160 1.375 ;
        RECT  6.035 0.675 6.105 1.375 ;
        RECT  5.745 1.145 6.035 1.375 ;
        RECT  5.675 0.975 5.745 1.375 ;
        RECT  5.410 1.145 5.675 1.375 ;
        RECT  5.290 1.005 5.410 1.375 ;
        RECT  5.050 1.145 5.290 1.375 ;
        RECT  4.930 1.005 5.050 1.375 ;
        RECT  4.690 1.145 4.930 1.375 ;
        RECT  4.570 1.005 4.690 1.375 ;
        RECT  4.330 1.145 4.570 1.375 ;
        RECT  4.210 1.005 4.330 1.375 ;
        RECT  2.680 1.145 4.210 1.375 ;
        RECT  2.560 1.060 2.680 1.375 ;
        RECT  1.440 1.145 2.560 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.355 5.635 0.465 ;
        RECT  5.565 0.775 5.635 0.905 ;
        RECT  5.495 0.185 5.565 0.465 ;
        RECT  5.495 0.775 5.565 1.065 ;
        RECT  5.145 0.705 5.230 0.795 ;
        RECT  5.145 0.185 5.205 0.485 ;
        RECT  4.775 0.185 4.795 0.485 ;
        RECT  4.750 0.705 4.795 0.795 ;
        RECT  5.400 0.545 5.540 0.615 ;
        RECT  5.330 0.545 5.400 0.935 ;
        RECT  4.680 0.865 5.330 0.935 ;
        RECT  4.610 0.395 4.680 0.935 ;
        RECT  4.485 0.395 4.610 0.465 ;
        RECT  4.485 0.865 4.610 0.935 ;
        RECT  4.415 0.185 4.485 0.465 ;
        RECT  4.415 0.735 4.485 1.035 ;
        RECT  4.150 0.545 4.460 0.615 ;
        RECT  4.150 0.260 4.415 0.330 ;
        RECT  3.270 0.855 4.415 0.925 ;
        RECT  4.080 0.205 4.150 0.330 ;
        RECT  4.080 0.400 4.150 0.780 ;
        RECT  3.595 0.205 4.080 0.275 ;
        RECT  3.820 0.400 4.080 0.470 ;
        RECT  3.455 0.710 4.080 0.780 ;
        RECT  3.720 0.995 3.840 1.075 ;
        RECT  3.180 0.995 3.720 1.065 ;
        RECT  3.525 0.205 3.595 0.400 ;
        RECT  3.325 0.330 3.525 0.400 ;
        RECT  3.385 0.520 3.455 0.780 ;
        RECT  3.255 0.330 3.325 0.450 ;
        RECT  3.185 0.685 3.290 0.755 ;
        RECT  3.115 0.205 3.185 0.755 ;
        RECT  3.110 0.965 3.180 1.065 ;
        RECT  2.710 0.205 3.115 0.275 ;
        RECT  3.045 0.965 3.110 1.035 ;
        RECT  2.975 0.360 3.045 1.035 ;
        RECT  2.850 0.690 2.905 1.040 ;
        RECT  2.835 0.360 2.850 1.040 ;
        RECT  2.780 0.360 2.835 0.760 ;
        RECT  2.280 0.690 2.780 0.760 ;
        RECT  2.640 0.205 2.710 0.440 ;
        RECT  2.570 0.510 2.690 0.615 ;
        RECT  2.360 0.370 2.640 0.440 ;
        RECT  2.025 0.510 2.570 0.580 ;
        RECT  2.320 0.830 2.530 0.900 ;
        RECT  2.290 0.195 2.360 0.440 ;
        RECT  2.260 0.830 2.320 0.910 ;
        RECT  2.040 0.195 2.290 0.265 ;
        RECT  2.160 0.665 2.280 0.760 ;
        RECT  2.050 0.840 2.260 0.910 ;
        RECT  1.965 0.340 2.025 0.580 ;
        RECT  1.955 0.340 1.965 0.930 ;
        RECT  1.895 0.510 1.955 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.655 0.350 1.725 0.795 ;
        RECT  1.540 0.350 1.655 0.420 ;
        RECT  1.510 0.725 1.655 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.940 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCND4BWP

MACRO SDFCNQD0BWP
    CLASS CORE ;
    FOREIGN SDFCNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.045 ;
        RECT  4.075 0.185 4.095 0.305 ;
        RECT  4.075 0.910 4.095 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.655 0.640 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 -0.115 4.200 0.115 ;
        RECT  3.860 -0.115 3.980 0.275 ;
        RECT  3.385 -0.115 3.860 0.115 ;
        RECT  3.315 -0.115 3.385 0.440 ;
        RECT  2.550 -0.115 3.315 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.145 4.200 1.375 ;
        RECT  3.860 1.120 3.980 1.375 ;
        RECT  3.580 1.145 3.860 1.375 ;
        RECT  3.460 1.135 3.580 1.375 ;
        RECT  2.660 1.145 3.460 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.000 0.520 4.020 0.640 ;
        RECT  3.930 0.350 4.000 1.050 ;
        RECT  3.585 0.350 3.930 0.420 ;
        RECT  3.420 0.980 3.930 1.050 ;
        RECT  3.765 0.520 3.835 0.910 ;
        RECT  3.120 0.840 3.765 0.910 ;
        RECT  3.515 0.230 3.585 0.420 ;
        RECT  3.300 0.980 3.420 1.060 ;
        RECT  3.175 0.695 3.290 0.765 ;
        RECT  3.105 0.205 3.175 0.765 ;
        RECT  3.045 0.840 3.120 1.070 ;
        RECT  2.690 0.205 3.105 0.275 ;
        RECT  3.025 0.840 3.045 0.910 ;
        RECT  2.955 0.345 3.025 0.910 ;
        RECT  2.840 0.690 2.885 1.040 ;
        RECT  2.815 0.345 2.840 1.040 ;
        RECT  2.770 0.345 2.815 0.760 ;
        RECT  2.260 0.690 2.770 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.320 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.255 0.830 2.320 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.030 0.840 2.255 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFCNQD0BWP

MACRO SDFCNQD1BWP
    CLASS CORE ;
    FOREIGN SDFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.045 ;
        RECT  4.075 0.185 4.095 0.465 ;
        RECT  4.075 0.735 4.095 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.495 3.655 0.640 ;
        RECT  3.535 0.495 3.625 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 -0.115 4.200 0.115 ;
        RECT  3.860 -0.115 3.980 0.275 ;
        RECT  3.385 -0.115 3.860 0.115 ;
        RECT  3.315 -0.115 3.385 0.440 ;
        RECT  2.550 -0.115 3.315 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.145 4.200 1.375 ;
        RECT  3.860 1.120 3.980 1.375 ;
        RECT  3.580 1.145 3.860 1.375 ;
        RECT  3.460 1.135 3.580 1.375 ;
        RECT  2.660 1.145 3.460 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.000 0.520 4.020 0.640 ;
        RECT  3.930 0.350 4.000 1.050 ;
        RECT  3.585 0.350 3.930 0.420 ;
        RECT  3.420 0.980 3.930 1.050 ;
        RECT  3.765 0.520 3.835 0.910 ;
        RECT  3.025 0.840 3.765 0.910 ;
        RECT  3.515 0.230 3.585 0.420 ;
        RECT  3.300 0.980 3.420 1.060 ;
        RECT  3.175 0.695 3.290 0.765 ;
        RECT  3.105 0.205 3.175 0.765 ;
        RECT  2.690 0.205 3.105 0.275 ;
        RECT  2.955 0.345 3.025 0.910 ;
        RECT  2.840 0.690 2.885 1.040 ;
        RECT  2.815 0.345 2.840 1.040 ;
        RECT  2.770 0.345 2.815 0.760 ;
        RECT  2.260 0.690 2.770 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.320 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.255 0.830 2.320 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.030 0.840 2.255 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCNQD1BWP

MACRO SDFCNQD2BWP
    CLASS CORE ;
    FOREIGN SDFCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 0.355 4.585 0.805 ;
        RECT  4.515 0.185 4.525 1.035 ;
        RECT  4.455 0.185 4.515 0.465 ;
        RECT  4.455 0.735 4.515 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.400 4.175 0.640 ;
        RECT  3.620 0.400 4.095 0.470 ;
        RECT  3.520 0.400 3.620 0.630 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 -0.115 4.760 0.115 ;
        RECT  4.635 -0.115 4.705 0.300 ;
        RECT  4.340 -0.115 4.635 0.115 ;
        RECT  4.220 -0.115 4.340 0.145 ;
        RECT  3.360 -0.115 4.220 0.115 ;
        RECT  3.240 -0.115 3.360 0.200 ;
        RECT  2.550 -0.115 3.240 0.115 ;
        RECT  2.480 -0.115 2.550 0.290 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.705 1.145 4.760 1.375 ;
        RECT  4.635 0.885 4.705 1.375 ;
        RECT  4.315 1.145 4.635 1.375 ;
        RECT  4.245 0.895 4.315 1.375 ;
        RECT  3.950 1.145 4.245 1.375 ;
        RECT  3.830 0.990 3.950 1.375 ;
        RECT  3.560 1.145 3.830 1.375 ;
        RECT  3.440 1.115 3.560 1.375 ;
        RECT  2.660 1.145 3.440 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.355 0.520 4.410 0.640 ;
        RECT  4.285 0.260 4.355 0.805 ;
        RECT  3.470 0.260 4.285 0.330 ;
        RECT  4.105 0.735 4.285 0.805 ;
        RECT  4.035 0.735 4.105 1.035 ;
        RECT  3.640 0.850 4.035 0.920 ;
        RECT  3.890 0.545 3.960 0.615 ;
        RECT  3.820 0.545 3.890 0.780 ;
        RECT  3.490 0.710 3.820 0.780 ;
        RECT  3.420 0.710 3.490 0.960 ;
        RECT  3.400 0.260 3.470 0.340 ;
        RECT  3.025 0.890 3.420 0.960 ;
        RECT  3.395 0.270 3.400 0.340 ;
        RECT  3.325 0.270 3.395 0.640 ;
        RECT  3.165 0.730 3.280 0.800 ;
        RECT  3.095 0.205 3.165 0.800 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  2.955 0.360 3.025 0.960 ;
        RECT  2.840 0.690 2.885 1.040 ;
        RECT  2.815 0.345 2.840 1.040 ;
        RECT  2.770 0.345 2.815 0.760 ;
        RECT  2.260 0.690 2.770 0.760 ;
        RECT  2.620 0.205 2.690 0.440 ;
        RECT  2.550 0.510 2.670 0.615 ;
        RECT  2.340 0.370 2.620 0.440 ;
        RECT  2.005 0.510 2.550 0.580 ;
        RECT  2.320 0.830 2.510 0.900 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.255 0.830 2.320 0.910 ;
        RECT  2.020 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.760 ;
        RECT  2.030 0.840 2.255 0.910 ;
        RECT  1.945 0.340 2.005 0.580 ;
        RECT  1.935 0.340 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCNQD2BWP

MACRO SDFCNQD4BWP
    CLASS CORE ;
    FOREIGN SDFCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.805 0.465 ;
        RECT  4.795 0.775 4.805 1.065 ;
        RECT  4.735 0.185 4.795 1.065 ;
        RECT  4.585 0.355 4.735 0.905 ;
        RECT  4.445 0.355 4.585 0.465 ;
        RECT  4.445 0.775 4.585 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.775 4.445 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.085 0.410 4.165 0.640 ;
        RECT  3.605 0.410 4.085 0.480 ;
        RECT  3.525 0.410 3.605 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.985 0.465 ;
        RECT  4.650 -0.115 4.915 0.115 ;
        RECT  4.530 -0.115 4.650 0.275 ;
        RECT  4.280 -0.115 4.530 0.115 ;
        RECT  4.160 -0.115 4.280 0.145 ;
        RECT  3.485 -0.115 4.160 0.115 ;
        RECT  3.365 -0.115 3.485 0.200 ;
        RECT  2.570 -0.115 3.365 0.115 ;
        RECT  2.500 -0.115 2.570 0.290 ;
        RECT  1.480 -0.115 2.500 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 1.145 5.040 1.375 ;
        RECT  4.915 0.675 4.985 1.375 ;
        RECT  4.625 1.145 4.915 1.375 ;
        RECT  4.555 0.975 4.625 1.375 ;
        RECT  4.255 1.145 4.555 1.375 ;
        RECT  4.185 0.895 4.255 1.375 ;
        RECT  3.910 1.145 4.185 1.375 ;
        RECT  3.790 0.990 3.910 1.375 ;
        RECT  3.550 1.145 3.790 1.375 ;
        RECT  3.430 1.135 3.550 1.375 ;
        RECT  2.680 1.145 3.430 1.375 ;
        RECT  2.560 1.060 2.680 1.375 ;
        RECT  1.440 1.145 2.560 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.355 4.515 0.465 ;
        RECT  4.445 0.775 4.515 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.775 4.445 1.065 ;
        RECT  4.305 0.545 4.410 0.615 ;
        RECT  4.235 0.270 4.305 0.805 ;
        RECT  3.385 0.270 4.235 0.340 ;
        RECT  4.065 0.735 4.235 0.805 ;
        RECT  3.995 0.735 4.065 1.035 ;
        RECT  3.600 0.850 3.995 0.920 ;
        RECT  3.905 0.550 3.970 0.620 ;
        RECT  3.835 0.550 3.905 0.780 ;
        RECT  3.440 0.710 3.835 0.780 ;
        RECT  3.370 0.710 3.440 0.955 ;
        RECT  3.315 0.270 3.385 0.640 ;
        RECT  3.045 0.885 3.370 0.955 ;
        RECT  3.185 0.730 3.300 0.800 ;
        RECT  3.115 0.205 3.185 0.800 ;
        RECT  2.710 0.205 3.115 0.275 ;
        RECT  2.975 0.360 3.045 0.955 ;
        RECT  2.850 0.690 2.905 1.040 ;
        RECT  2.835 0.360 2.850 1.040 ;
        RECT  2.780 0.360 2.835 0.760 ;
        RECT  2.280 0.690 2.780 0.760 ;
        RECT  2.640 0.205 2.710 0.440 ;
        RECT  2.570 0.510 2.690 0.615 ;
        RECT  2.360 0.370 2.640 0.440 ;
        RECT  2.025 0.510 2.570 0.580 ;
        RECT  2.340 0.830 2.530 0.900 ;
        RECT  2.290 0.195 2.360 0.440 ;
        RECT  2.275 0.830 2.340 0.910 ;
        RECT  2.040 0.195 2.290 0.265 ;
        RECT  2.160 0.665 2.280 0.760 ;
        RECT  2.050 0.840 2.275 0.910 ;
        RECT  1.965 0.340 2.025 0.580 ;
        RECT  1.955 0.340 1.965 0.930 ;
        RECT  1.895 0.510 1.955 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.655 0.350 1.725 0.795 ;
        RECT  1.540 0.350 1.655 0.420 ;
        RECT  1.510 0.725 1.655 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.940 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCNQD4BWP

MACRO SDFCSND0BWP
    CLASS CORE ;
    FOREIGN SDFCSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.760 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.195 5.005 1.045 ;
        RECT  4.915 0.195 4.935 0.315 ;
        RECT  4.915 0.910 4.935 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.695 0.775 4.730 1.045 ;
        RECT  4.625 0.350 4.695 1.045 ;
        RECT  4.535 0.350 4.625 0.470 ;
        RECT  4.540 0.920 4.625 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.495 4.165 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.140 ;
        RECT  4.070 -0.115 4.700 0.115 ;
        RECT  3.950 -0.115 4.070 0.275 ;
        RECT  2.560 -0.115 3.950 0.115 ;
        RECT  2.490 -0.115 2.560 0.290 ;
        RECT  1.440 -0.115 2.490 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 1.120 4.820 1.375 ;
        RECT  4.450 1.145 4.700 1.375 ;
        RECT  4.330 1.120 4.450 1.375 ;
        RECT  4.040 1.145 4.330 1.375 ;
        RECT  3.920 1.130 4.040 1.375 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 0.990 3.690 1.375 ;
        RECT  2.900 1.145 3.570 1.375 ;
        RECT  2.780 1.120 2.900 1.375 ;
        RECT  2.380 1.145 2.780 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.835 0.520 4.860 0.640 ;
        RECT  4.765 0.210 4.835 0.640 ;
        RECT  4.220 0.210 4.765 0.280 ;
        RECT  4.460 0.545 4.540 0.615 ;
        RECT  4.390 0.355 4.460 1.050 ;
        RECT  4.320 0.355 4.390 0.425 ;
        RECT  3.820 0.975 4.390 1.050 ;
        RECT  4.245 0.520 4.315 0.905 ;
        RECT  3.305 0.835 4.245 0.905 ;
        RECT  4.150 0.210 4.220 0.425 ;
        RECT  3.450 0.355 4.150 0.425 ;
        RECT  3.450 0.695 3.870 0.765 ;
        RECT  2.700 0.200 3.470 0.270 ;
        RECT  3.380 0.355 3.450 0.765 ;
        RECT  3.250 0.375 3.380 0.445 ;
        RECT  3.235 0.630 3.305 0.905 ;
        RECT  3.145 0.630 3.235 0.700 ;
        RECT  3.095 0.980 3.230 1.050 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  3.025 0.970 3.095 1.050 ;
        RECT  2.965 0.830 3.090 0.900 ;
        RECT  2.700 0.970 3.025 1.040 ;
        RECT  2.895 0.350 2.965 0.900 ;
        RECT  2.685 0.830 2.895 0.900 ;
        RECT  2.620 0.510 2.740 0.615 ;
        RECT  2.630 0.200 2.700 0.440 ;
        RECT  2.630 0.970 2.700 1.065 ;
        RECT  2.615 0.685 2.685 0.900 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.110 0.995 2.630 1.065 ;
        RECT  2.005 0.510 2.620 0.580 ;
        RECT  2.280 0.685 2.615 0.755 ;
        RECT  2.170 0.855 2.530 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.160 0.665 2.280 0.755 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.050 0.835 2.170 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.040 0.995 2.110 1.075 ;
        RECT  1.970 1.005 2.040 1.075 ;
        RECT  1.965 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.965 0.930 ;
        RECT  1.895 0.510 1.935 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFCSND0BWP

MACRO SDFCSND1BWP
    CLASS CORE ;
    FOREIGN SDFCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.760 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.045 ;
        RECT  4.915 0.185 4.935 0.465 ;
        RECT  4.915 0.750 4.935 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.695 0.775 4.730 1.045 ;
        RECT  4.625 0.350 4.695 1.045 ;
        RECT  4.535 0.350 4.625 0.470 ;
        RECT  4.540 0.775 4.625 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.495 4.165 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.140 ;
        RECT  4.070 -0.115 4.700 0.115 ;
        RECT  3.950 -0.115 4.070 0.275 ;
        RECT  2.560 -0.115 3.950 0.115 ;
        RECT  2.490 -0.115 2.560 0.290 ;
        RECT  1.440 -0.115 2.490 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 1.120 4.820 1.375 ;
        RECT  4.450 1.145 4.700 1.375 ;
        RECT  4.330 1.120 4.450 1.375 ;
        RECT  4.040 1.145 4.330 1.375 ;
        RECT  3.920 1.130 4.040 1.375 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 0.990 3.690 1.375 ;
        RECT  2.900 1.145 3.570 1.375 ;
        RECT  2.780 1.120 2.900 1.375 ;
        RECT  2.380 1.145 2.780 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.835 0.520 4.860 0.640 ;
        RECT  4.765 0.210 4.835 0.640 ;
        RECT  4.220 0.210 4.765 0.280 ;
        RECT  4.460 0.545 4.540 0.615 ;
        RECT  4.390 0.355 4.460 1.050 ;
        RECT  4.320 0.355 4.390 0.425 ;
        RECT  3.820 0.975 4.390 1.050 ;
        RECT  4.245 0.520 4.315 0.905 ;
        RECT  3.305 0.835 4.245 0.905 ;
        RECT  4.150 0.210 4.220 0.425 ;
        RECT  3.450 0.355 4.150 0.425 ;
        RECT  3.450 0.695 3.870 0.765 ;
        RECT  2.700 0.200 3.470 0.270 ;
        RECT  3.380 0.355 3.450 0.765 ;
        RECT  3.250 0.375 3.380 0.445 ;
        RECT  3.235 0.630 3.305 0.905 ;
        RECT  3.145 0.630 3.235 0.700 ;
        RECT  3.095 0.980 3.230 1.050 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  3.025 0.970 3.095 1.050 ;
        RECT  2.965 0.830 3.090 0.900 ;
        RECT  2.700 0.970 3.025 1.040 ;
        RECT  2.895 0.350 2.965 0.900 ;
        RECT  2.685 0.830 2.895 0.900 ;
        RECT  2.620 0.510 2.740 0.615 ;
        RECT  2.630 0.200 2.700 0.440 ;
        RECT  2.630 0.970 2.700 1.065 ;
        RECT  2.615 0.685 2.685 0.900 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.110 0.995 2.630 1.065 ;
        RECT  2.005 0.510 2.620 0.580 ;
        RECT  2.280 0.685 2.615 0.755 ;
        RECT  2.170 0.855 2.530 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.160 0.665 2.280 0.755 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.050 0.835 2.170 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.040 0.995 2.110 1.075 ;
        RECT  1.970 1.005 2.040 1.075 ;
        RECT  1.965 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.965 0.930 ;
        RECT  1.895 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.845 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.775 1.580 0.845 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSND1BWP

MACRO SDFCSND2BWP
    CLASS CORE ;
    FOREIGN SDFCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.600 0.540 3.675 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.355 5.145 0.810 ;
        RECT  5.075 0.185 5.085 1.040 ;
        RECT  5.015 0.185 5.075 0.465 ;
        RECT  5.015 0.740 5.075 1.040 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.690 0.350 4.760 1.045 ;
        RECT  4.620 0.350 4.690 0.450 ;
        RECT  4.655 0.735 4.690 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.495 4.165 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.300 ;
        RECT  4.920 -0.115 5.190 0.115 ;
        RECT  4.800 -0.115 4.920 0.140 ;
        RECT  4.540 -0.115 4.800 0.115 ;
        RECT  4.420 -0.115 4.540 0.140 ;
        RECT  4.010 -0.115 4.420 0.115 ;
        RECT  3.890 -0.115 4.010 0.275 ;
        RECT  2.555 -0.115 3.890 0.115 ;
        RECT  2.485 -0.115 2.555 0.290 ;
        RECT  1.440 -0.115 2.485 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 1.145 5.320 1.375 ;
        RECT  5.195 0.905 5.265 1.375 ;
        RECT  4.905 1.145 5.195 1.375 ;
        RECT  4.835 0.745 4.905 1.375 ;
        RECT  4.545 1.145 4.835 1.375 ;
        RECT  4.475 0.980 4.545 1.375 ;
        RECT  4.390 1.145 4.475 1.375 ;
        RECT  4.270 0.980 4.390 1.375 ;
        RECT  4.000 1.145 4.270 1.375 ;
        RECT  3.880 1.130 4.000 1.375 ;
        RECT  3.640 1.145 3.880 1.375 ;
        RECT  3.520 0.990 3.640 1.375 ;
        RECT  2.900 1.145 3.520 1.375 ;
        RECT  2.780 1.135 2.900 1.375 ;
        RECT  2.360 1.145 2.780 1.375 ;
        RECT  2.240 1.135 2.360 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.910 0.545 5.000 0.615 ;
        RECT  4.840 0.210 4.910 0.615 ;
        RECT  4.170 0.210 4.840 0.280 ;
        RECT  4.525 0.520 4.620 0.640 ;
        RECT  4.455 0.350 4.525 0.905 ;
        RECT  4.250 0.350 4.455 0.420 ;
        RECT  4.185 0.835 4.455 0.905 ;
        RECT  4.305 0.520 4.375 0.765 ;
        RECT  4.045 0.695 4.305 0.765 ;
        RECT  4.115 0.835 4.185 1.045 ;
        RECT  4.100 0.210 4.170 0.425 ;
        RECT  3.780 0.975 4.115 1.045 ;
        RECT  3.885 0.355 4.100 0.425 ;
        RECT  3.975 0.695 4.045 0.905 ;
        RECT  3.265 0.835 3.975 0.905 ;
        RECT  3.815 0.355 3.885 0.765 ;
        RECT  3.410 0.695 3.815 0.765 ;
        RECT  3.530 0.305 3.605 0.445 ;
        RECT  3.410 0.375 3.530 0.445 ;
        RECT  2.700 0.205 3.440 0.275 ;
        RECT  3.340 0.375 3.410 0.765 ;
        RECT  3.210 0.375 3.340 0.445 ;
        RECT  3.195 0.630 3.265 0.905 ;
        RECT  3.040 0.985 3.230 1.055 ;
        RECT  3.125 0.630 3.195 0.700 ;
        RECT  3.055 0.350 3.125 0.700 ;
        RECT  2.945 0.825 3.110 0.895 ;
        RECT  2.960 0.985 3.040 1.065 ;
        RECT  2.090 0.995 2.960 1.065 ;
        RECT  2.875 0.350 2.945 0.895 ;
        RECT  2.665 0.825 2.875 0.895 ;
        RECT  2.630 0.205 2.700 0.440 ;
        RECT  2.580 0.510 2.700 0.615 ;
        RECT  2.595 0.685 2.665 0.925 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.260 0.685 2.595 0.755 ;
        RECT  2.005 0.510 2.580 0.580 ;
        RECT  2.150 0.855 2.510 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.755 ;
        RECT  2.030 0.835 2.150 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.020 0.995 2.090 1.075 ;
        RECT  1.950 1.005 2.020 1.075 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.630 0.865 1.790 0.935 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.560 0.865 1.630 1.055 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSND2BWP

MACRO SDFCSND4BWP
    CLASS CORE ;
    FOREIGN SDFCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.745 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.185 6.065 0.465 ;
        RECT  6.055 0.775 6.065 1.055 ;
        RECT  5.995 0.185 6.055 1.055 ;
        RECT  5.845 0.355 5.995 0.905 ;
        RECT  5.705 0.355 5.845 0.465 ;
        RECT  5.705 0.775 5.845 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.775 5.705 1.055 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.350 5.350 0.470 ;
        RECT  5.255 0.775 5.325 1.055 ;
        RECT  5.215 0.775 5.255 0.905 ;
        RECT  5.005 0.350 5.215 0.905 ;
        RECT  4.880 0.350 5.005 0.470 ;
        RECT  4.985 0.775 5.005 0.905 ;
        RECT  4.895 0.775 4.985 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0584 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.585 0.495 4.670 0.640 ;
        RECT  4.515 0.495 4.585 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 -0.115 6.300 0.115 ;
        RECT  6.175 -0.115 6.245 0.465 ;
        RECT  5.885 -0.115 6.175 0.115 ;
        RECT  5.815 -0.115 5.885 0.280 ;
        RECT  5.540 -0.115 5.815 0.115 ;
        RECT  5.420 -0.115 5.540 0.140 ;
        RECT  5.160 -0.115 5.420 0.115 ;
        RECT  5.040 -0.115 5.160 0.140 ;
        RECT  4.780 -0.115 5.040 0.115 ;
        RECT  4.660 -0.115 4.780 0.140 ;
        RECT  4.015 -0.115 4.660 0.115 ;
        RECT  3.945 -0.115 4.015 0.270 ;
        RECT  2.575 -0.115 3.945 0.115 ;
        RECT  2.505 -0.115 2.575 0.290 ;
        RECT  1.480 -0.115 2.505 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 1.145 6.300 1.375 ;
        RECT  6.175 0.675 6.245 1.375 ;
        RECT  5.885 1.145 6.175 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  5.515 1.145 5.815 1.375 ;
        RECT  5.445 0.745 5.515 1.375 ;
        RECT  5.150 1.145 5.445 1.375 ;
        RECT  5.070 0.975 5.150 1.375 ;
        RECT  4.810 1.145 5.070 1.375 ;
        RECT  4.690 1.005 4.810 1.375 ;
        RECT  4.450 1.145 4.690 1.375 ;
        RECT  4.330 1.005 4.450 1.375 ;
        RECT  4.070 1.145 4.330 1.375 ;
        RECT  3.950 1.005 4.070 1.375 ;
        RECT  3.660 1.145 3.950 1.375 ;
        RECT  3.540 1.010 3.660 1.375 ;
        RECT  2.920 1.145 3.540 1.375 ;
        RECT  2.800 1.135 2.920 1.375 ;
        RECT  2.380 1.145 2.800 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.440 1.145 2.260 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.355 5.775 0.465 ;
        RECT  5.705 0.775 5.775 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.775 5.705 1.055 ;
        RECT  5.285 0.350 5.350 0.470 ;
        RECT  5.285 0.775 5.325 1.055 ;
        RECT  4.880 0.350 4.935 0.470 ;
        RECT  4.895 0.775 4.935 1.065 ;
        RECT  5.530 0.545 5.670 0.615 ;
        RECT  5.460 0.210 5.530 0.615 ;
        RECT  4.165 0.210 5.460 0.280 ;
        RECT  4.810 0.545 4.910 0.615 ;
        RECT  4.740 0.350 4.810 0.915 ;
        RECT  4.305 0.350 4.740 0.420 ;
        RECT  4.605 0.845 4.740 0.915 ;
        RECT  4.535 0.845 4.605 1.075 ;
        RECT  4.150 0.845 4.535 0.915 ;
        RECT  4.375 0.520 4.445 0.765 ;
        RECT  4.060 0.695 4.375 0.765 ;
        RECT  4.235 0.350 4.305 0.615 ;
        RECT  3.840 0.545 4.235 0.615 ;
        RECT  4.095 0.210 4.165 0.425 ;
        RECT  3.430 0.355 4.095 0.425 ;
        RECT  3.990 0.695 4.060 0.915 ;
        RECT  3.285 0.845 3.990 0.915 ;
        RECT  3.430 0.705 3.860 0.775 ;
        RECT  2.720 0.205 3.460 0.275 ;
        RECT  3.360 0.355 3.430 0.775 ;
        RECT  3.230 0.375 3.360 0.445 ;
        RECT  3.215 0.630 3.285 0.915 ;
        RECT  3.040 0.985 3.250 1.055 ;
        RECT  3.145 0.630 3.215 0.700 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  2.965 0.825 3.130 0.895 ;
        RECT  2.960 0.985 3.040 1.065 ;
        RECT  2.895 0.350 2.965 0.895 ;
        RECT  2.110 0.995 2.960 1.065 ;
        RECT  2.685 0.825 2.895 0.895 ;
        RECT  2.650 0.205 2.720 0.440 ;
        RECT  2.600 0.510 2.720 0.615 ;
        RECT  2.615 0.685 2.685 0.925 ;
        RECT  2.360 0.370 2.650 0.440 ;
        RECT  2.280 0.685 2.615 0.755 ;
        RECT  2.025 0.510 2.600 0.580 ;
        RECT  2.170 0.855 2.530 0.925 ;
        RECT  2.290 0.195 2.360 0.440 ;
        RECT  2.160 0.195 2.290 0.265 ;
        RECT  2.160 0.665 2.280 0.755 ;
        RECT  2.050 0.835 2.170 0.925 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.040 0.995 2.110 1.075 ;
        RECT  1.970 1.005 2.040 1.075 ;
        RECT  1.965 0.350 2.025 0.580 ;
        RECT  1.955 0.350 1.965 0.930 ;
        RECT  1.895 0.510 1.955 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.665 0.350 1.735 0.795 ;
        RECT  1.540 0.350 1.665 0.420 ;
        RECT  1.510 0.725 1.665 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.940 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSND4BWP

MACRO SDFCSNQD0BWP
    CLASS CORE ;
    FOREIGN SDFCSNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.625 0.505 3.675 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.215 4.725 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.495 4.065 0.640 ;
        RECT  3.955 0.495 4.045 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.115 4.760 0.115 ;
        RECT  4.455 -0.115 4.525 0.305 ;
        RECT  4.010 -0.115 4.455 0.115 ;
        RECT  3.890 -0.115 4.010 0.275 ;
        RECT  2.555 -0.115 3.890 0.115 ;
        RECT  2.485 -0.115 2.555 0.290 ;
        RECT  1.440 -0.115 2.485 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.145 4.760 1.375 ;
        RECT  4.455 0.920 4.525 1.375 ;
        RECT  4.380 1.145 4.455 1.375 ;
        RECT  4.260 1.120 4.380 1.375 ;
        RECT  4.000 1.145 4.260 1.375 ;
        RECT  3.880 1.110 4.000 1.375 ;
        RECT  3.640 1.145 3.880 1.375 ;
        RECT  3.520 0.990 3.640 1.375 ;
        RECT  2.900 1.145 3.520 1.375 ;
        RECT  2.780 1.135 2.900 1.375 ;
        RECT  2.360 1.145 2.780 1.375 ;
        RECT  2.240 1.135 2.360 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.385 0.545 4.560 0.615 ;
        RECT  4.345 0.350 4.385 1.045 ;
        RECT  4.315 0.185 4.345 1.045 ;
        RECT  4.275 0.185 4.315 0.420 ;
        RECT  4.070 0.975 4.315 1.045 ;
        RECT  3.885 0.350 4.275 0.420 ;
        RECT  4.175 0.520 4.245 0.905 ;
        RECT  3.990 0.835 4.175 0.905 ;
        RECT  3.920 0.835 3.990 0.920 ;
        RECT  3.265 0.850 3.920 0.920 ;
        RECT  3.815 0.350 3.885 0.630 ;
        RECT  3.410 0.710 3.840 0.780 ;
        RECT  3.530 0.280 3.605 0.425 ;
        RECT  3.410 0.355 3.530 0.425 ;
        RECT  2.700 0.205 3.440 0.275 ;
        RECT  3.340 0.355 3.410 0.780 ;
        RECT  3.210 0.375 3.340 0.445 ;
        RECT  3.195 0.630 3.265 0.920 ;
        RECT  3.035 0.990 3.230 1.060 ;
        RECT  3.125 0.630 3.195 0.700 ;
        RECT  3.055 0.350 3.125 0.700 ;
        RECT  2.945 0.825 3.110 0.895 ;
        RECT  2.940 0.990 3.035 1.065 ;
        RECT  2.875 0.350 2.945 0.895 ;
        RECT  2.090 0.995 2.940 1.065 ;
        RECT  2.665 0.825 2.875 0.895 ;
        RECT  2.630 0.205 2.700 0.440 ;
        RECT  2.580 0.510 2.700 0.615 ;
        RECT  2.595 0.685 2.665 0.925 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.260 0.685 2.595 0.755 ;
        RECT  2.005 0.510 2.580 0.580 ;
        RECT  2.150 0.855 2.510 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.755 ;
        RECT  2.030 0.835 2.150 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.020 0.995 2.090 1.075 ;
        RECT  1.950 1.005 2.020 1.075 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.660 0.575 1.730 0.645 ;
        RECT  1.590 0.350 1.660 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.725 1.590 0.795 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.480 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFCSNQD0BWP

MACRO SDFCSNQD1BWP
    CLASS CORE ;
    FOREIGN SDFCSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.630 ;
        RECT  3.600 0.550 3.675 0.630 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0803 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.195 4.725 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.495 4.065 0.640 ;
        RECT  3.955 0.495 4.045 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.115 4.760 0.115 ;
        RECT  4.455 -0.115 4.525 0.465 ;
        RECT  4.010 -0.115 4.455 0.115 ;
        RECT  3.890 -0.115 4.010 0.275 ;
        RECT  2.555 -0.115 3.890 0.115 ;
        RECT  2.485 -0.115 2.555 0.290 ;
        RECT  1.440 -0.115 2.485 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.145 4.760 1.375 ;
        RECT  4.455 0.760 4.525 1.375 ;
        RECT  4.000 1.145 4.455 1.375 ;
        RECT  3.880 1.110 4.000 1.375 ;
        RECT  3.640 1.145 3.880 1.375 ;
        RECT  3.520 0.990 3.640 1.375 ;
        RECT  2.900 1.145 3.520 1.375 ;
        RECT  2.780 1.135 2.900 1.375 ;
        RECT  2.360 1.145 2.780 1.375 ;
        RECT  2.240 1.135 2.360 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.385 0.545 4.560 0.615 ;
        RECT  4.345 0.350 4.385 1.065 ;
        RECT  4.315 0.185 4.345 1.065 ;
        RECT  4.275 0.185 4.315 0.420 ;
        RECT  4.070 0.995 4.315 1.065 ;
        RECT  3.885 0.350 4.275 0.420 ;
        RECT  4.175 0.520 4.245 0.920 ;
        RECT  3.265 0.850 4.175 0.920 ;
        RECT  3.815 0.350 3.885 0.630 ;
        RECT  3.410 0.710 3.840 0.780 ;
        RECT  3.530 0.280 3.605 0.445 ;
        RECT  3.410 0.375 3.530 0.445 ;
        RECT  2.700 0.205 3.440 0.275 ;
        RECT  3.340 0.375 3.410 0.780 ;
        RECT  3.210 0.375 3.340 0.445 ;
        RECT  3.195 0.630 3.265 0.920 ;
        RECT  3.035 0.990 3.230 1.060 ;
        RECT  3.125 0.630 3.195 0.700 ;
        RECT  3.055 0.350 3.125 0.700 ;
        RECT  2.945 0.825 3.110 0.895 ;
        RECT  2.940 0.990 3.035 1.065 ;
        RECT  2.875 0.350 2.945 0.895 ;
        RECT  2.090 0.995 2.940 1.065 ;
        RECT  2.665 0.825 2.875 0.895 ;
        RECT  2.630 0.205 2.700 0.440 ;
        RECT  2.580 0.510 2.700 0.615 ;
        RECT  2.595 0.685 2.665 0.925 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.260 0.685 2.595 0.755 ;
        RECT  2.005 0.510 2.580 0.580 ;
        RECT  2.150 0.855 2.510 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.755 ;
        RECT  2.030 0.835 2.150 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.020 0.995 2.090 1.075 ;
        RECT  1.950 1.005 2.020 1.075 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.650 0.875 1.790 0.945 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  1.580 0.350 1.650 0.805 ;
        RECT  1.580 0.875 1.650 1.055 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.735 1.580 0.805 ;
        RECT  0.685 0.985 1.580 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSNQD1BWP

MACRO SDFCSNQD2BWP
    CLASS CORE ;
    FOREIGN SDFCSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.630 ;
        RECT  3.600 0.530 3.675 0.630 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.355 5.005 0.905 ;
        RECT  4.935 0.185 4.945 1.065 ;
        RECT  4.875 0.185 4.935 0.465 ;
        RECT  4.875 0.765 4.935 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.585 0.520 4.635 0.640 ;
        RECT  4.515 0.410 4.585 0.640 ;
        RECT  4.165 0.410 4.515 0.480 ;
        RECT  4.095 0.410 4.165 0.765 ;
        RECT  3.990 0.540 4.095 0.620 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.300 ;
        RECT  4.780 -0.115 5.050 0.115 ;
        RECT  4.660 -0.115 4.780 0.145 ;
        RECT  3.980 -0.115 4.660 0.115 ;
        RECT  3.860 -0.115 3.980 0.200 ;
        RECT  2.555 -0.115 3.860 0.115 ;
        RECT  2.485 -0.115 2.555 0.290 ;
        RECT  1.440 -0.115 2.485 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.145 5.180 1.375 ;
        RECT  5.050 0.960 5.130 1.375 ;
        RECT  4.755 1.145 5.050 1.375 ;
        RECT  4.685 0.905 4.755 1.375 ;
        RECT  4.400 1.145 4.685 1.375 ;
        RECT  4.280 1.125 4.400 1.375 ;
        RECT  4.020 1.145 4.280 1.375 ;
        RECT  3.900 1.110 4.020 1.375 ;
        RECT  3.640 1.145 3.900 1.375 ;
        RECT  3.520 0.990 3.640 1.375 ;
        RECT  2.900 1.145 3.520 1.375 ;
        RECT  2.780 1.135 2.900 1.375 ;
        RECT  2.360 1.145 2.780 1.375 ;
        RECT  2.240 1.135 2.360 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.775 0.545 4.860 0.615 ;
        RECT  4.705 0.270 4.775 0.805 ;
        RECT  3.885 0.270 4.705 0.340 ;
        RECT  4.565 0.735 4.705 0.805 ;
        RECT  4.495 0.735 4.565 1.055 ;
        RECT  4.090 0.985 4.495 1.055 ;
        RECT  4.330 0.550 4.400 0.620 ;
        RECT  4.260 0.550 4.330 0.915 ;
        RECT  3.990 0.845 4.260 0.915 ;
        RECT  3.920 0.845 3.990 0.920 ;
        RECT  3.265 0.850 3.920 0.920 ;
        RECT  3.815 0.270 3.885 0.630 ;
        RECT  3.410 0.710 3.840 0.780 ;
        RECT  3.510 0.310 3.585 0.450 ;
        RECT  3.410 0.375 3.510 0.450 ;
        RECT  2.700 0.205 3.440 0.275 ;
        RECT  3.340 0.375 3.410 0.780 ;
        RECT  3.210 0.375 3.340 0.445 ;
        RECT  3.195 0.630 3.265 0.920 ;
        RECT  3.110 0.990 3.230 1.065 ;
        RECT  3.125 0.630 3.195 0.700 ;
        RECT  3.055 0.350 3.125 0.700 ;
        RECT  2.945 0.825 3.110 0.895 ;
        RECT  2.090 0.995 3.110 1.065 ;
        RECT  2.875 0.350 2.945 0.895 ;
        RECT  2.665 0.825 2.875 0.895 ;
        RECT  2.630 0.205 2.700 0.440 ;
        RECT  2.580 0.510 2.700 0.615 ;
        RECT  2.595 0.685 2.665 0.925 ;
        RECT  2.340 0.370 2.630 0.440 ;
        RECT  2.260 0.685 2.595 0.755 ;
        RECT  2.005 0.510 2.580 0.580 ;
        RECT  2.150 0.855 2.510 0.925 ;
        RECT  2.270 0.195 2.340 0.440 ;
        RECT  2.140 0.195 2.270 0.265 ;
        RECT  2.140 0.665 2.260 0.755 ;
        RECT  2.030 0.835 2.150 0.925 ;
        RECT  2.020 0.185 2.140 0.265 ;
        RECT  2.020 0.995 2.090 1.075 ;
        RECT  1.950 1.005 2.020 1.075 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.930 ;
        RECT  1.875 0.510 1.935 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.650 0.875 1.790 0.945 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  1.580 0.350 1.650 0.805 ;
        RECT  1.580 0.875 1.650 1.055 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.735 1.580 0.805 ;
        RECT  0.685 0.985 1.580 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSNQD2BWP

MACRO SDFCSNQD4BWP
    CLASS CORE ;
    FOREIGN SDFCSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.630 ;
        RECT  3.620 0.540 3.675 0.630 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.355 0.185 5.365 0.465 ;
        RECT  5.355 0.775 5.365 1.065 ;
        RECT  5.295 0.185 5.355 1.065 ;
        RECT  5.145 0.355 5.295 0.905 ;
        RECT  5.005 0.355 5.145 0.465 ;
        RECT  5.005 0.775 5.145 0.905 ;
        RECT  4.935 0.185 5.005 0.465 ;
        RECT  4.935 0.775 5.005 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.605 0.520 4.655 0.640 ;
        RECT  4.535 0.410 4.605 0.640 ;
        RECT  4.165 0.410 4.535 0.480 ;
        RECT  4.095 0.410 4.165 0.765 ;
        RECT  4.000 0.545 4.095 0.615 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 -0.115 5.600 0.115 ;
        RECT  5.475 -0.115 5.545 0.465 ;
        RECT  5.210 -0.115 5.475 0.115 ;
        RECT  5.090 -0.115 5.210 0.280 ;
        RECT  4.820 -0.115 5.090 0.115 ;
        RECT  4.700 -0.115 4.820 0.145 ;
        RECT  4.000 -0.115 4.700 0.115 ;
        RECT  3.880 -0.115 4.000 0.200 ;
        RECT  2.575 -0.115 3.880 0.115 ;
        RECT  2.505 -0.115 2.575 0.290 ;
        RECT  1.480 -0.115 2.505 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 1.145 5.600 1.375 ;
        RECT  5.475 0.685 5.545 1.375 ;
        RECT  5.190 1.145 5.475 1.375 ;
        RECT  5.110 0.975 5.190 1.375 ;
        RECT  4.795 1.145 5.110 1.375 ;
        RECT  4.725 0.905 4.795 1.375 ;
        RECT  4.420 1.145 4.725 1.375 ;
        RECT  4.300 1.125 4.420 1.375 ;
        RECT  4.040 1.145 4.300 1.375 ;
        RECT  3.920 1.110 4.040 1.375 ;
        RECT  3.660 1.145 3.920 1.375 ;
        RECT  3.540 0.990 3.660 1.375 ;
        RECT  2.920 1.145 3.540 1.375 ;
        RECT  2.800 1.135 2.920 1.375 ;
        RECT  2.380 1.145 2.800 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.440 1.145 2.260 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.005 0.355 5.075 0.465 ;
        RECT  5.005 0.775 5.075 0.905 ;
        RECT  4.935 0.185 5.005 0.465 ;
        RECT  4.935 0.775 5.005 1.065 ;
        RECT  4.800 0.545 4.940 0.615 ;
        RECT  4.730 0.270 4.800 0.805 ;
        RECT  3.895 0.270 4.730 0.340 ;
        RECT  4.585 0.735 4.730 0.805 ;
        RECT  4.515 0.735 4.585 1.055 ;
        RECT  4.110 0.985 4.515 1.055 ;
        RECT  4.350 0.550 4.420 0.620 ;
        RECT  4.280 0.550 4.350 0.915 ;
        RECT  3.285 0.845 4.280 0.915 ;
        RECT  3.825 0.270 3.895 0.630 ;
        RECT  3.430 0.705 3.860 0.775 ;
        RECT  3.530 0.310 3.605 0.450 ;
        RECT  3.430 0.375 3.530 0.450 ;
        RECT  2.720 0.205 3.460 0.275 ;
        RECT  3.360 0.375 3.430 0.775 ;
        RECT  3.230 0.375 3.360 0.445 ;
        RECT  3.215 0.630 3.285 0.915 ;
        RECT  3.130 0.990 3.250 1.065 ;
        RECT  3.145 0.630 3.215 0.700 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  2.965 0.825 3.130 0.895 ;
        RECT  2.110 0.995 3.130 1.065 ;
        RECT  2.895 0.350 2.965 0.895 ;
        RECT  2.685 0.825 2.895 0.895 ;
        RECT  2.650 0.205 2.720 0.440 ;
        RECT  2.600 0.510 2.720 0.615 ;
        RECT  2.615 0.685 2.685 0.925 ;
        RECT  2.360 0.370 2.650 0.440 ;
        RECT  2.280 0.685 2.615 0.755 ;
        RECT  2.025 0.510 2.600 0.580 ;
        RECT  2.170 0.855 2.530 0.925 ;
        RECT  2.290 0.195 2.360 0.440 ;
        RECT  2.160 0.195 2.290 0.265 ;
        RECT  2.160 0.665 2.280 0.755 ;
        RECT  2.050 0.835 2.170 0.925 ;
        RECT  2.040 0.185 2.160 0.265 ;
        RECT  2.040 0.995 2.110 1.075 ;
        RECT  1.970 1.005 2.040 1.075 ;
        RECT  1.965 0.350 2.025 0.580 ;
        RECT  1.955 0.350 1.965 0.930 ;
        RECT  1.895 0.510 1.955 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.665 0.350 1.735 0.795 ;
        RECT  1.540 0.350 1.665 0.420 ;
        RECT  1.510 0.725 1.665 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.940 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFCSNQD4BWP

MACRO SDFD0BWP
    CLASS CORE ;
    FOREIGN SDFD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.350 4.025 0.905 ;
        RECT  3.935 0.350 3.955 0.470 ;
        RECT  3.935 0.710 3.955 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.350 3.410 0.420 ;
        RECT  3.325 0.790 3.385 0.910 ;
        RECT  3.255 0.350 3.325 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.700 -0.115 3.820 0.140 ;
        RECT  3.200 -0.115 3.700 0.115 ;
        RECT  3.080 -0.115 3.200 0.130 ;
        RECT  2.360 -0.115 3.080 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 1.145 4.060 1.375 ;
        RECT  3.700 1.130 3.820 1.375 ;
        RECT  3.240 1.145 3.700 1.375 ;
        RECT  3.120 1.130 3.240 1.375 ;
        RECT  2.380 1.145 3.120 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.885 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.075 0.210 3.790 0.280 ;
        RECT  3.650 0.520 3.720 1.060 ;
        RECT  3.630 0.520 3.650 0.640 ;
        RECT  2.765 0.990 3.650 1.060 ;
        RECT  3.560 0.350 3.610 0.420 ;
        RECT  3.560 0.790 3.580 0.910 ;
        RECT  3.490 0.350 3.560 0.910 ;
        RECT  3.395 0.520 3.490 0.640 ;
        RECT  3.005 0.210 3.075 0.920 ;
        RECT  2.940 0.315 3.005 0.415 ;
        RECT  2.910 0.850 3.005 0.920 ;
        RECT  2.870 0.500 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.570 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.480 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFD0BWP

MACRO SDFD1BWP
    CLASS CORE ;
    FOREIGN SDFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.350 3.410 0.420 ;
        RECT  3.325 0.790 3.385 0.910 ;
        RECT  3.255 0.350 3.325 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.700 -0.115 3.820 0.140 ;
        RECT  3.200 -0.115 3.700 0.115 ;
        RECT  3.080 -0.115 3.200 0.130 ;
        RECT  2.360 -0.115 3.080 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 1.145 4.060 1.375 ;
        RECT  3.700 1.130 3.820 1.375 ;
        RECT  3.220 1.145 3.700 1.375 ;
        RECT  3.100 1.130 3.220 1.375 ;
        RECT  2.380 1.145 3.100 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.885 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.075 0.210 3.790 0.280 ;
        RECT  3.650 0.520 3.720 1.060 ;
        RECT  3.630 0.520 3.650 0.640 ;
        RECT  2.765 0.990 3.650 1.060 ;
        RECT  3.560 0.350 3.610 0.420 ;
        RECT  3.560 0.790 3.580 0.910 ;
        RECT  3.490 0.350 3.560 0.910 ;
        RECT  3.395 0.520 3.490 0.640 ;
        RECT  3.005 0.210 3.075 0.920 ;
        RECT  2.940 0.325 3.005 0.425 ;
        RECT  2.910 0.850 3.005 0.920 ;
        RECT  2.870 0.500 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.570 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFD1BWP

MACRO SDFD2BWP
    CLASS CORE ;
    FOREIGN SDFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.805 ;
        RECT  4.235 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.235 0.465 ;
        RECT  4.175 0.735 4.235 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.350 3.885 0.910 ;
        RECT  3.795 0.350 3.815 0.470 ;
        RECT  3.795 0.770 3.815 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.300 ;
        RECT  4.080 -0.115 4.350 0.115 ;
        RECT  3.960 -0.115 4.080 0.140 ;
        RECT  3.650 -0.115 3.960 0.115 ;
        RECT  3.530 -0.115 3.650 0.140 ;
        RECT  3.260 -0.115 3.530 0.115 ;
        RECT  3.140 -0.115 3.260 0.140 ;
        RECT  2.360 -0.115 3.140 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.905 4.430 1.375 ;
        RECT  4.080 1.145 4.350 1.375 ;
        RECT  3.960 1.120 4.080 1.375 ;
        RECT  3.650 1.145 3.960 1.375 ;
        RECT  3.530 1.120 3.650 1.375 ;
        RECT  3.280 1.145 3.530 1.375 ;
        RECT  3.160 1.120 3.280 1.375 ;
        RECT  2.380 1.145 3.160 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.545 4.160 0.615 ;
        RECT  4.000 0.210 4.070 1.050 ;
        RECT  3.020 0.210 4.000 0.280 ;
        RECT  3.070 0.980 4.000 1.050 ;
        RECT  3.680 0.520 3.745 0.640 ;
        RECT  3.610 0.365 3.680 0.830 ;
        RECT  3.160 0.365 3.610 0.435 ;
        RECT  3.445 0.760 3.610 0.830 ;
        RECT  3.375 0.760 3.445 0.900 ;
        RECT  3.300 0.545 3.400 0.615 ;
        RECT  3.230 0.545 3.300 0.910 ;
        RECT  2.765 0.840 3.230 0.910 ;
        RECT  3.090 0.365 3.160 0.615 ;
        RECT  3.040 0.545 3.090 0.615 ;
        RECT  2.930 0.980 3.070 1.065 ;
        RECT  2.950 0.185 3.020 0.465 ;
        RECT  2.870 0.580 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.650 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFD2BWP

MACRO SDFD4BWP
    CLASS CORE ;
    FOREIGN SDFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.775 4.945 1.065 ;
        RECT  4.795 0.355 4.875 0.465 ;
        RECT  4.795 0.775 4.875 0.905 ;
        RECT  4.585 0.355 4.795 0.905 ;
        RECT  4.565 0.355 4.585 0.465 ;
        RECT  4.495 0.775 4.585 1.075 ;
        RECT  4.495 0.185 4.565 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.710 4.230 0.800 ;
        RECT  4.095 0.355 4.210 0.445 ;
        RECT  3.885 0.355 4.095 0.800 ;
        RECT  3.710 0.355 3.885 0.445 ;
        RECT  3.750 0.710 3.885 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.055 -0.115 5.125 0.465 ;
        RECT  4.755 -0.115 5.055 0.115 ;
        RECT  4.685 -0.115 4.755 0.285 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.145 ;
        RECT  4.020 -0.115 4.280 0.115 ;
        RECT  3.900 -0.115 4.020 0.145 ;
        RECT  3.640 -0.115 3.900 0.115 ;
        RECT  3.520 -0.115 3.640 0.145 ;
        RECT  3.260 -0.115 3.520 0.115 ;
        RECT  3.140 -0.115 3.260 0.145 ;
        RECT  2.380 -0.115 3.140 0.115 ;
        RECT  2.260 -0.115 2.380 0.125 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.055 0.685 5.125 1.375 ;
        RECT  4.755 1.145 5.055 1.375 ;
        RECT  4.685 0.975 4.755 1.375 ;
        RECT  4.410 1.145 4.685 1.375 ;
        RECT  4.290 1.010 4.410 1.375 ;
        RECT  4.050 1.145 4.290 1.375 ;
        RECT  3.930 1.010 4.050 1.375 ;
        RECT  3.680 1.145 3.930 1.375 ;
        RECT  3.560 1.010 3.680 1.375 ;
        RECT  3.300 1.145 3.560 1.375 ;
        RECT  3.180 1.130 3.300 1.375 ;
        RECT  2.400 1.145 3.180 1.375 ;
        RECT  2.280 0.870 2.400 1.375 ;
        RECT  1.440 1.145 2.280 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.775 4.945 1.065 ;
        RECT  4.865 0.355 4.875 0.465 ;
        RECT  4.865 0.775 4.875 0.905 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.775 4.515 1.075 ;
        RECT  4.165 0.710 4.230 0.800 ;
        RECT  4.165 0.355 4.210 0.445 ;
        RECT  3.710 0.355 3.815 0.445 ;
        RECT  3.750 0.710 3.815 0.800 ;
        RECT  4.370 0.545 4.490 0.615 ;
        RECT  4.300 0.215 4.370 0.940 ;
        RECT  3.030 0.215 4.300 0.285 ;
        RECT  3.475 0.870 4.300 0.940 ;
        RECT  3.600 0.545 3.780 0.615 ;
        RECT  3.530 0.365 3.600 0.800 ;
        RECT  3.170 0.365 3.530 0.435 ;
        RECT  3.380 0.700 3.530 0.800 ;
        RECT  3.405 0.870 3.475 1.060 ;
        RECT  3.310 0.545 3.450 0.615 ;
        RECT  2.920 0.990 3.405 1.060 ;
        RECT  3.240 0.545 3.310 0.920 ;
        RECT  2.795 0.850 3.240 0.920 ;
        RECT  3.100 0.365 3.170 0.630 ;
        RECT  3.070 0.530 3.100 0.630 ;
        RECT  2.960 0.215 3.030 0.425 ;
        RECT  2.890 0.710 3.000 0.780 ;
        RECT  2.820 0.195 2.890 0.780 ;
        RECT  2.700 0.195 2.820 0.265 ;
        RECT  2.750 0.850 2.795 1.070 ;
        RECT  2.725 0.350 2.750 1.070 ;
        RECT  2.680 0.350 2.725 0.920 ;
        RECT  2.580 0.185 2.700 0.265 ;
        RECT  2.540 0.355 2.610 1.040 ;
        RECT  2.040 0.195 2.580 0.265 ;
        RECT  2.470 0.355 2.540 0.425 ;
        RECT  2.535 0.730 2.540 1.040 ;
        RECT  2.275 0.730 2.535 0.800 ;
        RECT  2.400 0.510 2.470 0.640 ;
        RECT  2.025 0.510 2.400 0.580 ;
        RECT  2.205 0.650 2.275 0.800 ;
        RECT  1.965 0.350 2.025 0.580 ;
        RECT  1.955 0.350 1.965 0.950 ;
        RECT  1.895 0.510 1.955 0.950 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.655 0.350 1.725 0.795 ;
        RECT  1.540 0.350 1.655 0.420 ;
        RECT  1.510 0.725 1.655 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.940 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFD4BWP

MACRO SDFKCND0BWP
    CLASS CORE ;
    FOREIGN SDFKCND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0232 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.335 4.445 0.905 ;
        RECT  4.355 0.335 4.375 0.455 ;
        RECT  4.360 0.765 4.375 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.355 4.045 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.625 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 -0.115 4.480 0.115 ;
        RECT  4.140 -0.115 4.260 0.420 ;
        RECT  3.685 -0.115 4.140 0.115 ;
        RECT  3.615 -0.115 3.685 0.280 ;
        RECT  2.915 -0.115 3.615 0.115 ;
        RECT  2.845 -0.115 2.915 0.420 ;
        RECT  2.000 -0.115 2.845 0.115 ;
        RECT  1.880 -0.115 2.000 0.135 ;
        RECT  1.440 -0.115 1.880 0.115 ;
        RECT  1.320 -0.115 1.440 0.265 ;
        RECT  1.040 -0.115 1.320 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.235 1.145 4.480 1.375 ;
        RECT  4.165 1.010 4.235 1.375 ;
        RECT  3.700 1.145 4.165 1.375 ;
        RECT  3.580 1.120 3.700 1.375 ;
        RECT  2.940 1.145 3.580 1.375 ;
        RECT  2.820 0.870 2.940 1.375 ;
        RECT  2.000 1.145 2.820 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.440 1.145 1.880 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.010 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.280 0.520 4.305 0.650 ;
        RECT  4.210 0.520 4.280 0.940 ;
        RECT  3.880 0.870 4.210 0.940 ;
        RECT  3.865 0.460 3.880 0.940 ;
        RECT  3.810 0.185 3.865 0.940 ;
        RECT  3.795 0.185 3.810 0.530 ;
        RECT  3.760 0.870 3.810 0.940 ;
        RECT  3.500 0.460 3.795 0.530 ;
        RECT  3.580 0.635 3.735 0.755 ;
        RECT  3.510 0.635 3.580 1.050 ;
        RECT  3.400 0.635 3.510 0.705 ;
        RECT  3.180 0.980 3.510 1.050 ;
        RECT  3.260 0.825 3.430 0.895 ;
        RECT  3.330 0.195 3.400 0.705 ;
        RECT  3.210 0.195 3.330 0.265 ;
        RECT  3.190 0.410 3.260 0.895 ;
        RECT  3.105 0.220 3.120 0.800 ;
        RECT  3.050 0.220 3.105 1.050 ;
        RECT  3.035 0.730 3.050 1.050 ;
        RECT  2.795 0.730 3.035 0.800 ;
        RECT  2.910 0.510 2.980 0.640 ;
        RECT  2.535 0.510 2.910 0.580 ;
        RECT  2.725 0.680 2.795 0.800 ;
        RECT  2.530 0.300 2.535 0.580 ;
        RECT  2.460 0.300 2.530 0.960 ;
        RECT  2.320 0.205 2.390 0.935 ;
        RECT  1.605 0.205 2.320 0.275 ;
        RECT  2.250 0.865 2.320 1.040 ;
        RECT  1.690 0.970 2.250 1.040 ;
        RECT  2.165 0.355 2.235 0.765 ;
        RECT  2.070 0.355 2.165 0.425 ;
        RECT  2.095 0.695 2.165 0.850 ;
        RECT  1.980 0.545 2.080 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.690 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.535 0.205 1.605 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.250 0.665 0.990 ;
        RECT  0.485 0.215 0.525 0.920 ;
        RECT  0.455 0.215 0.485 1.020 ;
        RECT  0.390 0.215 0.455 0.285 ;
        RECT  0.415 0.850 0.455 1.020 ;
        RECT  0.125 0.850 0.415 0.920 ;
        RECT  0.055 0.850 0.125 1.020 ;
    END
END SDFKCND0BWP

MACRO SDFKCND1BWP
    CLASS CORE ;
    FOREIGN SDFKCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.185 4.445 1.045 ;
        RECT  4.355 0.185 4.375 0.465 ;
        RECT  4.355 0.735 4.375 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.215 4.045 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.240 -0.115 4.480 0.115 ;
        RECT  4.160 -0.115 4.240 0.440 ;
        RECT  3.685 -0.115 4.160 0.115 ;
        RECT  3.615 -0.115 3.685 0.280 ;
        RECT  2.915 -0.115 3.615 0.115 ;
        RECT  2.845 -0.115 2.915 0.420 ;
        RECT  2.000 -0.115 2.845 0.115 ;
        RECT  1.880 -0.115 2.000 0.135 ;
        RECT  1.440 -0.115 1.880 0.115 ;
        RECT  1.320 -0.115 1.440 0.265 ;
        RECT  1.040 -0.115 1.320 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.145 4.480 1.375 ;
        RECT  4.140 1.025 4.260 1.375 ;
        RECT  3.700 1.145 4.140 1.375 ;
        RECT  3.580 1.120 3.700 1.375 ;
        RECT  2.940 1.145 3.580 1.375 ;
        RECT  2.820 0.870 2.940 1.375 ;
        RECT  2.000 1.145 2.820 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.440 1.145 1.880 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.280 0.520 4.305 0.640 ;
        RECT  4.210 0.520 4.280 0.940 ;
        RECT  3.880 0.870 4.210 0.940 ;
        RECT  3.865 0.460 3.880 0.940 ;
        RECT  3.810 0.185 3.865 0.940 ;
        RECT  3.795 0.185 3.810 0.530 ;
        RECT  3.760 0.870 3.810 0.940 ;
        RECT  3.500 0.460 3.795 0.530 ;
        RECT  3.580 0.635 3.735 0.755 ;
        RECT  3.510 0.635 3.580 1.050 ;
        RECT  3.400 0.635 3.510 0.705 ;
        RECT  3.180 0.980 3.510 1.050 ;
        RECT  3.260 0.825 3.430 0.895 ;
        RECT  3.330 0.195 3.400 0.705 ;
        RECT  3.210 0.195 3.330 0.265 ;
        RECT  3.190 0.410 3.260 0.895 ;
        RECT  3.105 0.220 3.120 0.800 ;
        RECT  3.050 0.220 3.105 1.050 ;
        RECT  3.035 0.730 3.050 1.050 ;
        RECT  2.795 0.730 3.035 0.800 ;
        RECT  2.910 0.510 2.980 0.640 ;
        RECT  2.535 0.510 2.910 0.580 ;
        RECT  2.725 0.680 2.795 0.800 ;
        RECT  2.530 0.300 2.535 0.580 ;
        RECT  2.460 0.300 2.530 0.960 ;
        RECT  2.320 0.205 2.390 0.935 ;
        RECT  1.605 0.205 2.320 0.275 ;
        RECT  2.250 0.865 2.320 1.040 ;
        RECT  1.690 0.970 2.250 1.040 ;
        RECT  2.165 0.355 2.235 0.765 ;
        RECT  2.070 0.355 2.165 0.425 ;
        RECT  2.095 0.695 2.165 0.850 ;
        RECT  1.980 0.545 2.080 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.690 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.535 0.205 1.605 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCND1BWP

MACRO SDFKCND2BWP
    CLASS CORE ;
    FOREIGN SDFKCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 0.355 4.585 0.805 ;
        RECT  4.515 0.185 4.525 1.035 ;
        RECT  4.455 0.185 4.515 0.465 ;
        RECT  4.455 0.735 4.515 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.195 4.165 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.300 ;
        RECT  4.345 -0.115 4.630 0.115 ;
        RECT  4.275 -0.115 4.345 0.465 ;
        RECT  3.985 -0.115 4.275 0.115 ;
        RECT  3.915 -0.115 3.985 0.475 ;
        RECT  3.625 -0.115 3.915 0.115 ;
        RECT  3.555 -0.115 3.625 0.260 ;
        RECT  2.885 -0.115 3.555 0.115 ;
        RECT  2.815 -0.115 2.885 0.420 ;
        RECT  1.980 -0.115 2.815 0.115 ;
        RECT  1.860 -0.115 1.980 0.135 ;
        RECT  1.440 -0.115 1.860 0.115 ;
        RECT  1.320 -0.115 1.440 0.265 ;
        RECT  1.040 -0.115 1.320 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.905 4.710 1.375 ;
        RECT  4.370 1.145 4.630 1.375 ;
        RECT  4.250 1.010 4.370 1.375 ;
        RECT  4.010 1.145 4.250 1.375 ;
        RECT  3.890 1.010 4.010 1.375 ;
        RECT  3.640 1.145 3.890 1.375 ;
        RECT  3.520 1.120 3.640 1.375 ;
        RECT  2.900 1.145 3.520 1.375 ;
        RECT  2.780 0.870 2.900 1.375 ;
        RECT  1.980 1.145 2.780 1.375 ;
        RECT  1.860 1.110 1.980 1.375 ;
        RECT  1.440 1.145 1.860 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.370 0.545 4.440 0.615 ;
        RECT  4.300 0.545 4.370 0.940 ;
        RECT  3.840 0.870 4.300 0.940 ;
        RECT  3.805 0.460 3.840 0.940 ;
        RECT  3.770 0.185 3.805 0.940 ;
        RECT  3.735 0.185 3.770 0.530 ;
        RECT  3.700 0.870 3.770 0.940 ;
        RECT  3.460 0.460 3.735 0.530 ;
        RECT  3.520 0.635 3.695 0.755 ;
        RECT  3.450 0.635 3.520 1.050 ;
        RECT  3.370 0.635 3.450 0.705 ;
        RECT  3.140 0.980 3.450 1.050 ;
        RECT  3.230 0.815 3.380 0.885 ;
        RECT  3.300 0.185 3.370 0.705 ;
        RECT  3.170 0.185 3.300 0.255 ;
        RECT  3.160 0.440 3.230 0.885 ;
        RECT  3.065 0.220 3.090 0.800 ;
        RECT  3.020 0.220 3.065 1.050 ;
        RECT  3.005 0.220 3.020 0.340 ;
        RECT  2.995 0.730 3.020 1.050 ;
        RECT  2.755 0.730 2.995 0.800 ;
        RECT  2.880 0.510 2.950 0.640 ;
        RECT  2.515 0.510 2.880 0.580 ;
        RECT  2.685 0.680 2.755 0.800 ;
        RECT  2.510 0.300 2.515 0.580 ;
        RECT  2.440 0.300 2.510 0.960 ;
        RECT  2.300 0.205 2.370 0.935 ;
        RECT  1.605 0.205 2.300 0.275 ;
        RECT  2.230 0.865 2.300 1.040 ;
        RECT  1.690 0.970 2.230 1.040 ;
        RECT  2.145 0.355 2.215 0.765 ;
        RECT  2.050 0.355 2.145 0.425 ;
        RECT  2.075 0.695 2.145 0.850 ;
        RECT  1.980 0.545 2.065 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.690 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.535 0.205 1.605 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCND2BWP

MACRO SDFKCND4BWP
    CLASS CORE ;
    FOREIGN SDFKCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.185 5.785 0.465 ;
        RECT  5.775 0.765 5.785 1.065 ;
        RECT  5.715 0.185 5.775 1.065 ;
        RECT  5.565 0.355 5.715 0.905 ;
        RECT  5.425 0.355 5.565 0.465 ;
        RECT  5.425 0.765 5.565 0.905 ;
        RECT  5.355 0.185 5.425 0.465 ;
        RECT  5.355 0.765 5.425 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.700 5.090 0.800 ;
        RECT  4.995 0.185 5.065 0.485 ;
        RECT  4.935 0.355 4.995 0.485 ;
        RECT  4.725 0.355 4.935 0.800 ;
        RECT  4.705 0.355 4.725 0.485 ;
        RECT  4.610 0.700 4.725 0.800 ;
        RECT  4.635 0.185 4.705 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 -0.115 6.020 0.115 ;
        RECT  5.890 -0.115 5.970 0.465 ;
        RECT  5.630 -0.115 5.890 0.115 ;
        RECT  5.510 -0.115 5.630 0.275 ;
        RECT  5.245 -0.115 5.510 0.115 ;
        RECT  5.175 -0.115 5.245 0.465 ;
        RECT  4.910 -0.115 5.175 0.115 ;
        RECT  4.790 -0.115 4.910 0.275 ;
        RECT  4.525 -0.115 4.790 0.115 ;
        RECT  4.455 -0.115 4.525 0.305 ;
        RECT  4.165 -0.115 4.455 0.115 ;
        RECT  4.095 -0.115 4.165 0.320 ;
        RECT  3.245 -0.115 4.095 0.115 ;
        RECT  3.175 -0.115 3.245 0.460 ;
        RECT  2.885 -0.115 3.175 0.115 ;
        RECT  2.815 -0.115 2.885 0.400 ;
        RECT  1.980 -0.115 2.815 0.115 ;
        RECT  1.860 -0.115 1.980 0.135 ;
        RECT  1.430 -0.115 1.860 0.115 ;
        RECT  1.310 -0.115 1.430 0.265 ;
        RECT  1.040 -0.115 1.310 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 1.145 6.020 1.375 ;
        RECT  5.890 0.675 5.970 1.375 ;
        RECT  5.605 1.145 5.890 1.375 ;
        RECT  5.535 0.975 5.605 1.375 ;
        RECT  5.270 1.145 5.535 1.375 ;
        RECT  5.150 1.010 5.270 1.375 ;
        RECT  4.910 1.145 5.150 1.375 ;
        RECT  4.790 1.010 4.910 1.375 ;
        RECT  4.550 1.145 4.790 1.375 ;
        RECT  4.430 1.010 4.550 1.375 ;
        RECT  4.170 1.145 4.430 1.375 ;
        RECT  4.100 0.950 4.170 1.375 ;
        RECT  3.245 1.145 4.100 1.375 ;
        RECT  3.175 0.850 3.245 1.375 ;
        RECT  2.885 1.145 3.175 1.375 ;
        RECT  2.815 0.860 2.885 1.375 ;
        RECT  2.000 1.145 2.815 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.440 1.145 1.880 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.355 5.495 0.465 ;
        RECT  5.425 0.765 5.495 0.905 ;
        RECT  5.355 0.185 5.425 0.465 ;
        RECT  5.355 0.765 5.425 1.065 ;
        RECT  5.005 0.700 5.090 0.800 ;
        RECT  5.005 0.185 5.065 0.485 ;
        RECT  4.635 0.185 4.655 0.485 ;
        RECT  4.610 0.700 4.655 0.800 ;
        RECT  5.250 0.545 5.390 0.615 ;
        RECT  5.180 0.545 5.250 0.940 ;
        RECT  4.500 0.870 5.180 0.940 ;
        RECT  4.430 0.435 4.500 0.940 ;
        RECT  4.345 0.435 4.430 0.505 ;
        RECT  4.345 0.870 4.430 0.940 ;
        RECT  4.275 0.200 4.345 0.505 ;
        RECT  4.275 0.870 4.345 1.010 ;
        RECT  4.030 0.585 4.310 0.655 ;
        RECT  4.000 0.435 4.275 0.505 ;
        RECT  3.960 0.585 4.030 1.055 ;
        RECT  3.920 0.585 3.960 0.655 ;
        RECT  3.425 0.985 3.960 1.055 ;
        RECT  3.850 0.270 3.920 0.655 ;
        RECT  3.800 0.780 3.890 0.910 ;
        RECT  3.805 0.270 3.850 0.340 ;
        RECT  3.735 0.195 3.805 0.340 ;
        RECT  3.750 0.780 3.800 0.850 ;
        RECT  3.680 0.485 3.750 0.850 ;
        RECT  3.420 0.195 3.735 0.265 ;
        RECT  3.630 0.485 3.680 0.555 ;
        RECT  3.560 0.335 3.630 0.405 ;
        RECT  3.560 0.710 3.605 0.890 ;
        RECT  3.535 0.335 3.560 0.890 ;
        RECT  3.490 0.335 3.535 0.780 ;
        RECT  3.105 0.710 3.490 0.780 ;
        RECT  3.355 0.850 3.425 1.055 ;
        RECT  3.350 0.195 3.420 0.350 ;
        RECT  3.065 0.335 3.105 0.780 ;
        RECT  3.035 0.335 3.065 0.980 ;
        RECT  2.970 0.335 3.035 0.405 ;
        RECT  2.995 0.710 3.035 0.980 ;
        RECT  2.775 0.710 2.995 0.780 ;
        RECT  2.885 0.510 2.955 0.640 ;
        RECT  2.525 0.510 2.885 0.580 ;
        RECT  2.705 0.660 2.775 0.780 ;
        RECT  2.515 0.510 2.525 0.980 ;
        RECT  2.445 0.280 2.515 0.980 ;
        RECT  2.320 0.205 2.375 0.935 ;
        RECT  2.305 0.205 2.320 1.040 ;
        RECT  1.585 0.205 2.305 0.275 ;
        RECT  2.250 0.865 2.305 1.040 ;
        RECT  1.690 0.970 2.250 1.040 ;
        RECT  2.165 0.355 2.235 0.765 ;
        RECT  2.050 0.355 2.165 0.425 ;
        RECT  2.095 0.695 2.165 0.850 ;
        RECT  1.980 0.545 2.080 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.670 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.515 0.205 1.585 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCND4BWP

MACRO SDFKCNQD0BWP
    CLASS CORE ;
    FOREIGN SDFKCNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.665 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.630 0.825 0.905 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0096 ;
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.195 4.025 1.045 ;
        RECT  3.935 0.195 3.955 0.415 ;
        RECT  3.935 0.905 3.955 1.045 ;
        RECT  3.705 0.345 3.935 0.415 ;
        RECT  3.635 0.345 3.705 0.610 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.770 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.015 0.640 ;
        RECT  1.850 0.495 1.925 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.770 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 -0.115 4.060 0.115 ;
        RECT  3.720 -0.115 3.840 0.255 ;
        RECT  3.045 -0.115 3.720 0.115 ;
        RECT  2.975 -0.115 3.045 0.420 ;
        RECT  2.120 -0.115 2.975 0.115 ;
        RECT  2.000 -0.115 2.120 0.125 ;
        RECT  1.620 -0.115 2.000 0.115 ;
        RECT  1.500 -0.115 1.620 0.125 ;
        RECT  0.860 -0.115 1.500 0.115 ;
        RECT  0.760 -0.115 0.860 0.400 ;
        RECT  0.510 -0.115 0.760 0.115 ;
        RECT  0.390 -0.115 0.510 0.270 ;
        RECT  0.000 -0.115 0.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.145 4.060 1.375 ;
        RECT  3.760 0.915 3.830 1.375 ;
        RECT  3.060 1.145 3.760 1.375 ;
        RECT  2.940 0.870 3.060 1.375 ;
        RECT  2.120 1.145 2.940 1.375 ;
        RECT  2.000 1.130 2.120 1.375 ;
        RECT  1.620 1.145 2.000 1.375 ;
        RECT  1.500 1.135 1.620 1.375 ;
        RECT  0.840 1.145 1.500 1.375 ;
        RECT  0.720 1.135 0.840 1.375 ;
        RECT  0.540 1.145 0.720 1.375 ;
        RECT  0.420 1.135 0.540 1.375 ;
        RECT  0.125 1.145 0.420 1.375 ;
        RECT  0.055 0.890 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.815 0.510 3.885 0.750 ;
        RECT  3.690 0.680 3.815 0.750 ;
        RECT  3.620 0.680 3.690 1.060 ;
        RECT  3.530 0.680 3.620 0.750 ;
        RECT  3.300 0.990 3.620 1.060 ;
        RECT  3.390 0.830 3.540 0.900 ;
        RECT  3.460 0.195 3.530 0.750 ;
        RECT  3.330 0.195 3.460 0.265 ;
        RECT  3.320 0.430 3.390 0.900 ;
        RECT  3.225 0.220 3.250 0.800 ;
        RECT  3.180 0.220 3.225 1.050 ;
        RECT  3.165 0.220 3.180 0.340 ;
        RECT  3.155 0.730 3.180 1.050 ;
        RECT  2.935 0.730 3.155 0.800 ;
        RECT  3.040 0.510 3.110 0.640 ;
        RECT  2.675 0.510 3.040 0.580 ;
        RECT  2.865 0.675 2.935 0.800 ;
        RECT  2.665 0.300 2.675 0.580 ;
        RECT  2.595 0.300 2.665 0.960 ;
        RECT  1.220 0.195 2.520 0.265 ;
        RECT  2.415 0.840 2.485 1.060 ;
        RECT  1.100 0.990 2.415 1.060 ;
        RECT  2.310 0.340 2.375 0.765 ;
        RECT  2.305 0.340 2.310 0.850 ;
        RECT  2.235 0.340 2.305 0.460 ;
        RECT  2.235 0.695 2.305 0.850 ;
        RECT  2.155 0.520 2.190 0.640 ;
        RECT  2.085 0.355 2.155 0.915 ;
        RECT  1.850 0.355 2.085 0.425 ;
        RECT  1.850 0.845 2.085 0.915 ;
        RECT  1.465 0.335 1.770 0.405 ;
        RECT  1.465 0.845 1.770 0.915 ;
        RECT  1.395 0.335 1.465 0.915 ;
        RECT  1.215 0.475 1.285 0.760 ;
        RECT  1.120 0.195 1.220 0.400 ;
        RECT  0.665 0.475 1.215 0.545 ;
        RECT  1.000 0.665 1.130 0.735 ;
        RECT  0.930 0.665 1.000 1.065 ;
        RECT  0.525 0.995 0.930 1.065 ;
        RECT  0.595 0.190 0.665 0.910 ;
        RECT  0.455 0.350 0.525 1.065 ;
        RECT  0.130 0.350 0.455 0.420 ;
        RECT  0.210 0.920 0.455 0.990 ;
        RECT  0.055 0.190 0.130 0.420 ;
    END
END SDFKCNQD0BWP

MACRO SDFKCNQD1BWP
    CLASS CORE ;
    FOREIGN SDFKCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.195 4.165 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.965 -0.115 4.200 0.115 ;
        RECT  3.895 -0.115 3.965 0.305 ;
        RECT  3.605 -0.115 3.895 0.115 ;
        RECT  3.535 -0.115 3.605 0.285 ;
        RECT  2.865 -0.115 3.535 0.115 ;
        RECT  2.795 -0.115 2.865 0.420 ;
        RECT  1.960 -0.115 2.795 0.115 ;
        RECT  1.840 -0.115 1.960 0.135 ;
        RECT  1.430 -0.115 1.840 0.115 ;
        RECT  1.310 -0.115 1.430 0.265 ;
        RECT  1.040 -0.115 1.310 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.965 1.145 4.200 1.375 ;
        RECT  3.895 0.905 3.965 1.375 ;
        RECT  3.610 1.145 3.895 1.375 ;
        RECT  3.540 0.955 3.610 1.375 ;
        RECT  2.890 1.145 3.540 1.375 ;
        RECT  2.770 0.870 2.890 1.375 ;
        RECT  1.980 1.145 2.770 1.375 ;
        RECT  1.860 1.110 1.980 1.375 ;
        RECT  1.440 1.145 1.860 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.925 0.395 3.995 0.820 ;
        RECT  3.785 0.395 3.925 0.465 ;
        RECT  3.785 0.750 3.925 0.820 ;
        RECT  3.470 0.545 3.830 0.615 ;
        RECT  3.715 0.185 3.785 0.465 ;
        RECT  3.715 0.750 3.785 1.075 ;
        RECT  3.440 0.395 3.715 0.465 ;
        RECT  3.400 0.545 3.470 1.060 ;
        RECT  3.350 0.545 3.400 0.615 ;
        RECT  3.130 0.990 3.400 1.060 ;
        RECT  3.280 0.195 3.350 0.615 ;
        RECT  3.210 0.800 3.330 0.920 ;
        RECT  3.150 0.195 3.280 0.265 ;
        RECT  3.140 0.440 3.210 0.920 ;
        RECT  3.045 0.220 3.070 0.800 ;
        RECT  3.000 0.220 3.045 1.050 ;
        RECT  2.985 0.220 3.000 0.340 ;
        RECT  2.975 0.730 3.000 1.050 ;
        RECT  2.755 0.730 2.975 0.800 ;
        RECT  2.860 0.510 2.930 0.640 ;
        RECT  2.510 0.510 2.860 0.580 ;
        RECT  2.685 0.680 2.755 0.800 ;
        RECT  2.495 0.510 2.510 0.960 ;
        RECT  2.425 0.300 2.495 0.960 ;
        RECT  2.300 0.205 2.355 0.935 ;
        RECT  2.285 0.205 2.300 1.040 ;
        RECT  1.585 0.205 2.285 0.275 ;
        RECT  2.230 0.865 2.285 1.040 ;
        RECT  1.690 0.970 2.230 1.040 ;
        RECT  2.145 0.355 2.215 0.765 ;
        RECT  2.030 0.355 2.145 0.425 ;
        RECT  2.075 0.695 2.145 0.850 ;
        RECT  1.950 0.545 2.065 0.615 ;
        RECT  1.880 0.355 1.950 0.855 ;
        RECT  1.670 0.355 1.880 0.425 ;
        RECT  1.715 0.735 1.880 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.515 0.205 1.585 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCNQD1BWP

MACRO SDFKCNQD2BWP
    CLASS CORE ;
    FOREIGN SDFKCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.805 ;
        RECT  4.235 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.235 0.465 ;
        RECT  4.175 0.735 4.235 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.300 ;
        RECT  4.065 -0.115 4.350 0.115 ;
        RECT  3.995 -0.115 4.065 0.305 ;
        RECT  3.685 -0.115 3.995 0.115 ;
        RECT  3.615 -0.115 3.685 0.290 ;
        RECT  2.925 -0.115 3.615 0.115 ;
        RECT  2.855 -0.115 2.925 0.420 ;
        RECT  2.000 -0.115 2.855 0.115 ;
        RECT  1.880 -0.115 2.000 0.135 ;
        RECT  1.440 -0.115 1.880 0.115 ;
        RECT  1.320 -0.115 1.440 0.265 ;
        RECT  1.040 -0.115 1.320 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.905 4.430 1.375 ;
        RECT  4.065 1.145 4.350 1.375 ;
        RECT  3.995 0.905 4.065 1.375 ;
        RECT  3.700 1.145 3.995 1.375 ;
        RECT  3.580 1.120 3.700 1.375 ;
        RECT  2.940 1.145 3.580 1.375 ;
        RECT  2.820 0.870 2.940 1.375 ;
        RECT  2.000 1.145 2.820 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.440 1.145 1.880 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.025 0.395 4.095 0.835 ;
        RECT  3.865 0.395 4.025 0.465 ;
        RECT  3.865 0.765 4.025 0.835 ;
        RECT  3.580 0.545 3.900 0.615 ;
        RECT  3.795 0.190 3.865 0.465 ;
        RECT  3.795 0.765 3.865 1.070 ;
        RECT  3.520 0.395 3.795 0.465 ;
        RECT  3.510 0.545 3.580 1.050 ;
        RECT  3.410 0.545 3.510 0.615 ;
        RECT  3.180 0.980 3.510 1.050 ;
        RECT  3.270 0.815 3.420 0.885 ;
        RECT  3.340 0.185 3.410 0.615 ;
        RECT  3.210 0.185 3.340 0.255 ;
        RECT  3.200 0.440 3.270 0.885 ;
        RECT  3.105 0.220 3.130 0.800 ;
        RECT  3.060 0.220 3.105 1.050 ;
        RECT  3.045 0.220 3.060 0.340 ;
        RECT  3.035 0.730 3.060 1.050 ;
        RECT  2.795 0.730 3.035 0.800 ;
        RECT  2.920 0.510 2.990 0.640 ;
        RECT  2.535 0.510 2.920 0.580 ;
        RECT  2.725 0.680 2.795 0.800 ;
        RECT  2.530 0.300 2.535 0.580 ;
        RECT  2.460 0.300 2.530 0.960 ;
        RECT  2.320 0.205 2.390 0.935 ;
        RECT  1.605 0.205 2.320 0.275 ;
        RECT  2.250 0.865 2.320 1.040 ;
        RECT  1.690 0.970 2.250 1.040 ;
        RECT  2.165 0.355 2.235 0.765 ;
        RECT  2.070 0.355 2.165 0.425 ;
        RECT  2.095 0.695 2.165 0.850 ;
        RECT  1.980 0.545 2.080 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.690 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.535 0.205 1.605 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCNQD2BWP

MACRO SDFKCNQD4BWP
    CLASS CORE ;
    FOREIGN SDFKCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.925 0.500 0.995 0.650 ;
        RECT  0.805 0.500 0.925 0.570 ;
        RECT  0.735 0.215 0.805 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0320 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.650 ;
        RECT  1.260 0.520 1.295 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.185 5.085 0.465 ;
        RECT  5.075 0.765 5.085 1.065 ;
        RECT  5.015 0.185 5.075 1.065 ;
        RECT  4.865 0.355 5.015 0.905 ;
        RECT  4.730 0.355 4.865 0.465 ;
        RECT  4.730 0.765 4.865 0.905 ;
        RECT  4.660 0.185 4.730 0.465 ;
        RECT  4.660 0.765 4.730 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.540 1.750 0.620 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.355 0.385 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.930 -0.115 5.190 0.115 ;
        RECT  4.810 -0.115 4.930 0.275 ;
        RECT  4.545 -0.115 4.810 0.115 ;
        RECT  4.475 -0.115 4.545 0.305 ;
        RECT  4.165 -0.115 4.475 0.115 ;
        RECT  4.095 -0.115 4.165 0.320 ;
        RECT  3.245 -0.115 4.095 0.115 ;
        RECT  3.175 -0.115 3.245 0.460 ;
        RECT  2.885 -0.115 3.175 0.115 ;
        RECT  2.815 -0.115 2.885 0.400 ;
        RECT  1.980 -0.115 2.815 0.115 ;
        RECT  1.860 -0.115 1.980 0.135 ;
        RECT  1.430 -0.115 1.860 0.115 ;
        RECT  1.310 -0.115 1.430 0.265 ;
        RECT  1.040 -0.115 1.310 0.115 ;
        RECT  0.970 -0.115 1.040 0.430 ;
        RECT  0.125 -0.115 0.970 0.115 ;
        RECT  0.055 -0.115 0.125 0.345 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.675 5.270 1.375 ;
        RECT  4.905 1.145 5.190 1.375 ;
        RECT  4.835 0.975 4.905 1.375 ;
        RECT  4.545 1.145 4.835 1.375 ;
        RECT  4.475 0.905 4.545 1.375 ;
        RECT  4.170 1.145 4.475 1.375 ;
        RECT  4.100 0.940 4.170 1.375 ;
        RECT  3.270 1.145 4.100 1.375 ;
        RECT  3.150 0.880 3.270 1.375 ;
        RECT  2.885 1.145 3.150 1.375 ;
        RECT  2.815 0.860 2.885 1.375 ;
        RECT  2.000 1.145 2.815 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.440 1.145 1.880 1.375 ;
        RECT  1.320 1.110 1.440 1.375 ;
        RECT  1.100 1.145 1.320 1.375 ;
        RECT  0.980 1.040 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.355 4.795 0.465 ;
        RECT  4.730 0.765 4.795 0.905 ;
        RECT  4.660 0.185 4.730 0.465 ;
        RECT  4.660 0.765 4.730 1.065 ;
        RECT  4.520 0.395 4.590 0.835 ;
        RECT  4.345 0.395 4.520 0.465 ;
        RECT  4.345 0.765 4.520 0.835 ;
        RECT  4.030 0.545 4.450 0.615 ;
        RECT  4.275 0.200 4.345 0.465 ;
        RECT  4.275 0.765 4.345 1.070 ;
        RECT  4.000 0.395 4.275 0.465 ;
        RECT  3.960 0.545 4.030 1.055 ;
        RECT  3.920 0.545 3.960 0.615 ;
        RECT  3.425 0.985 3.960 1.055 ;
        RECT  3.850 0.270 3.920 0.615 ;
        RECT  3.800 0.780 3.890 0.910 ;
        RECT  3.805 0.270 3.850 0.340 ;
        RECT  3.735 0.195 3.805 0.340 ;
        RECT  3.750 0.780 3.800 0.850 ;
        RECT  3.680 0.485 3.750 0.850 ;
        RECT  3.420 0.195 3.735 0.265 ;
        RECT  3.630 0.485 3.680 0.555 ;
        RECT  3.560 0.335 3.630 0.405 ;
        RECT  3.560 0.710 3.605 0.890 ;
        RECT  3.535 0.335 3.560 0.890 ;
        RECT  3.490 0.335 3.535 0.780 ;
        RECT  3.105 0.710 3.490 0.780 ;
        RECT  3.355 0.850 3.425 1.055 ;
        RECT  3.350 0.195 3.420 0.350 ;
        RECT  3.065 0.335 3.105 0.780 ;
        RECT  3.035 0.335 3.065 0.980 ;
        RECT  2.970 0.335 3.035 0.405 ;
        RECT  2.995 0.710 3.035 0.980 ;
        RECT  2.775 0.710 2.995 0.780 ;
        RECT  2.885 0.510 2.955 0.640 ;
        RECT  2.525 0.510 2.885 0.580 ;
        RECT  2.705 0.660 2.775 0.780 ;
        RECT  2.515 0.510 2.525 0.980 ;
        RECT  2.445 0.280 2.515 0.980 ;
        RECT  2.320 0.205 2.375 0.935 ;
        RECT  2.305 0.205 2.320 1.040 ;
        RECT  1.585 0.205 2.305 0.275 ;
        RECT  2.250 0.865 2.305 1.040 ;
        RECT  1.690 0.970 2.250 1.040 ;
        RECT  2.165 0.355 2.235 0.765 ;
        RECT  2.050 0.355 2.165 0.425 ;
        RECT  2.095 0.695 2.165 0.850 ;
        RECT  1.980 0.545 2.080 0.615 ;
        RECT  1.910 0.355 1.980 0.855 ;
        RECT  1.670 0.355 1.910 0.425 ;
        RECT  1.715 0.735 1.910 0.855 ;
        RECT  1.620 0.970 1.690 1.060 ;
        RECT  1.510 0.990 1.620 1.060 ;
        RECT  1.515 0.205 1.585 0.410 ;
        RECT  1.435 0.510 1.505 0.910 ;
        RECT  1.405 0.840 1.435 0.910 ;
        RECT  1.345 0.840 1.405 0.930 ;
        RECT  0.665 0.860 1.345 0.930 ;
        RECT  1.190 0.720 1.280 0.790 ;
        RECT  1.190 0.190 1.225 0.310 ;
        RECT  1.120 0.190 1.190 0.790 ;
        RECT  0.815 0.720 1.120 0.790 ;
        RECT  0.745 0.640 0.815 0.790 ;
        RECT  0.595 0.200 0.665 1.075 ;
        RECT  0.485 0.205 0.525 0.915 ;
        RECT  0.455 0.205 0.485 1.075 ;
        RECT  0.370 0.205 0.455 0.275 ;
        RECT  0.415 0.845 0.455 1.075 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCNQD4BWP

MACRO SDFKCSND0BWP
    CLASS CORE ;
    FOREIGN SDFKCSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0246 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.335 5.005 0.905 ;
        RECT  4.915 0.335 4.935 0.455 ;
        RECT  4.920 0.765 4.935 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.355 4.605 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0126 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.760 0.795 0.875 0.865 ;
        RECT  0.345 0.380 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.420 ;
        RECT  4.245 -0.115 4.700 0.115 ;
        RECT  4.175 -0.115 4.245 0.280 ;
        RECT  3.475 -0.115 4.175 0.115 ;
        RECT  3.405 -0.115 3.475 0.420 ;
        RECT  2.560 -0.115 3.405 0.115 ;
        RECT  2.440 -0.115 2.560 0.135 ;
        RECT  2.000 -0.115 2.440 0.115 ;
        RECT  1.880 -0.115 2.000 0.265 ;
        RECT  1.600 -0.115 1.880 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.795 1.145 5.040 1.375 ;
        RECT  4.725 1.010 4.795 1.375 ;
        RECT  4.260 1.145 4.725 1.375 ;
        RECT  4.140 1.120 4.260 1.375 ;
        RECT  3.500 1.145 4.140 1.375 ;
        RECT  3.380 0.870 3.500 1.375 ;
        RECT  2.560 1.145 3.380 1.375 ;
        RECT  2.440 1.110 2.560 1.375 ;
        RECT  2.000 1.145 2.440 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.010 1.660 1.375 ;
        RECT  0.900 1.145 1.540 1.375 ;
        RECT  0.780 1.110 0.900 1.375 ;
        RECT  0.330 1.145 0.780 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.840 0.520 4.865 0.650 ;
        RECT  4.770 0.520 4.840 0.940 ;
        RECT  4.440 0.870 4.770 0.940 ;
        RECT  4.425 0.460 4.440 0.940 ;
        RECT  4.370 0.185 4.425 0.940 ;
        RECT  4.355 0.185 4.370 0.530 ;
        RECT  4.320 0.870 4.370 0.940 ;
        RECT  4.060 0.460 4.355 0.530 ;
        RECT  4.140 0.635 4.295 0.755 ;
        RECT  4.070 0.635 4.140 1.050 ;
        RECT  3.960 0.635 4.070 0.705 ;
        RECT  3.740 0.980 4.070 1.050 ;
        RECT  3.820 0.825 3.990 0.895 ;
        RECT  3.890 0.195 3.960 0.705 ;
        RECT  3.770 0.195 3.890 0.265 ;
        RECT  3.750 0.410 3.820 0.895 ;
        RECT  3.665 0.220 3.680 0.800 ;
        RECT  3.610 0.220 3.665 1.050 ;
        RECT  3.595 0.730 3.610 1.050 ;
        RECT  3.355 0.730 3.595 0.800 ;
        RECT  3.470 0.510 3.540 0.640 ;
        RECT  3.095 0.510 3.470 0.580 ;
        RECT  3.285 0.680 3.355 0.800 ;
        RECT  3.090 0.300 3.095 0.580 ;
        RECT  3.020 0.300 3.090 0.960 ;
        RECT  2.880 0.205 2.950 0.935 ;
        RECT  2.165 0.205 2.880 0.275 ;
        RECT  2.810 0.865 2.880 1.040 ;
        RECT  2.250 0.970 2.810 1.040 ;
        RECT  2.725 0.355 2.795 0.765 ;
        RECT  2.630 0.355 2.725 0.425 ;
        RECT  2.655 0.695 2.725 0.850 ;
        RECT  2.540 0.545 2.640 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.250 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.095 0.205 2.165 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.225 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.155 0.250 1.225 0.990 ;
        RECT  1.045 0.335 1.085 1.005 ;
        RECT  1.015 0.235 1.045 1.005 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.670 0.935 1.015 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSND0BWP

MACRO SDFKCSND1BWP
    CLASS CORE ;
    FOREIGN SDFKCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.045 ;
        RECT  4.915 0.185 4.935 0.465 ;
        RECT  4.915 0.735 4.935 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.215 4.605 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.800 -0.115 5.040 0.115 ;
        RECT  4.720 -0.115 4.800 0.440 ;
        RECT  4.245 -0.115 4.720 0.115 ;
        RECT  4.175 -0.115 4.245 0.280 ;
        RECT  3.475 -0.115 4.175 0.115 ;
        RECT  3.405 -0.115 3.475 0.420 ;
        RECT  2.560 -0.115 3.405 0.115 ;
        RECT  2.440 -0.115 2.560 0.135 ;
        RECT  2.000 -0.115 2.440 0.115 ;
        RECT  1.880 -0.115 2.000 0.265 ;
        RECT  1.600 -0.115 1.880 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 1.025 4.820 1.375 ;
        RECT  4.260 1.145 4.700 1.375 ;
        RECT  4.140 1.120 4.260 1.375 ;
        RECT  3.500 1.145 4.140 1.375 ;
        RECT  3.380 0.870 3.500 1.375 ;
        RECT  2.560 1.145 3.380 1.375 ;
        RECT  2.440 1.110 2.560 1.375 ;
        RECT  2.000 1.145 2.440 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.840 0.520 4.865 0.640 ;
        RECT  4.770 0.520 4.840 0.940 ;
        RECT  4.440 0.870 4.770 0.940 ;
        RECT  4.425 0.460 4.440 0.940 ;
        RECT  4.370 0.185 4.425 0.940 ;
        RECT  4.355 0.185 4.370 0.530 ;
        RECT  4.320 0.870 4.370 0.940 ;
        RECT  4.060 0.460 4.355 0.530 ;
        RECT  4.140 0.635 4.295 0.755 ;
        RECT  4.070 0.635 4.140 1.050 ;
        RECT  3.960 0.635 4.070 0.705 ;
        RECT  3.740 0.980 4.070 1.050 ;
        RECT  3.820 0.825 3.990 0.895 ;
        RECT  3.890 0.195 3.960 0.705 ;
        RECT  3.770 0.195 3.890 0.265 ;
        RECT  3.750 0.410 3.820 0.895 ;
        RECT  3.665 0.220 3.680 0.800 ;
        RECT  3.610 0.220 3.665 1.050 ;
        RECT  3.595 0.730 3.610 1.050 ;
        RECT  3.355 0.730 3.595 0.800 ;
        RECT  3.470 0.510 3.540 0.640 ;
        RECT  3.095 0.510 3.470 0.580 ;
        RECT  3.285 0.680 3.355 0.800 ;
        RECT  3.090 0.300 3.095 0.580 ;
        RECT  3.020 0.300 3.090 0.960 ;
        RECT  2.880 0.205 2.950 0.935 ;
        RECT  2.165 0.205 2.880 0.275 ;
        RECT  2.810 0.865 2.880 1.040 ;
        RECT  2.250 0.970 2.810 1.040 ;
        RECT  2.725 0.355 2.795 0.765 ;
        RECT  2.630 0.355 2.725 0.425 ;
        RECT  2.655 0.695 2.725 0.850 ;
        RECT  2.540 0.545 2.640 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.250 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.095 0.205 2.165 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSND1BWP

MACRO SDFKCSND2BWP
    CLASS CORE ;
    FOREIGN SDFKCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.355 5.145 0.805 ;
        RECT  5.075 0.185 5.085 1.035 ;
        RECT  5.015 0.185 5.075 0.465 ;
        RECT  5.015 0.735 5.075 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.195 4.725 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.300 ;
        RECT  4.905 -0.115 5.190 0.115 ;
        RECT  4.835 -0.115 4.905 0.465 ;
        RECT  4.545 -0.115 4.835 0.115 ;
        RECT  4.475 -0.115 4.545 0.475 ;
        RECT  4.185 -0.115 4.475 0.115 ;
        RECT  4.115 -0.115 4.185 0.260 ;
        RECT  3.445 -0.115 4.115 0.115 ;
        RECT  3.375 -0.115 3.445 0.420 ;
        RECT  2.540 -0.115 3.375 0.115 ;
        RECT  2.420 -0.115 2.540 0.135 ;
        RECT  2.000 -0.115 2.420 0.115 ;
        RECT  1.880 -0.115 2.000 0.265 ;
        RECT  1.600 -0.115 1.880 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.905 5.270 1.375 ;
        RECT  4.930 1.145 5.190 1.375 ;
        RECT  4.810 1.010 4.930 1.375 ;
        RECT  4.570 1.145 4.810 1.375 ;
        RECT  4.450 1.010 4.570 1.375 ;
        RECT  4.200 1.145 4.450 1.375 ;
        RECT  4.080 1.120 4.200 1.375 ;
        RECT  3.460 1.145 4.080 1.375 ;
        RECT  3.340 0.870 3.460 1.375 ;
        RECT  2.540 1.145 3.340 1.375 ;
        RECT  2.420 1.110 2.540 1.375 ;
        RECT  2.000 1.145 2.420 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.930 0.545 5.000 0.615 ;
        RECT  4.860 0.545 4.930 0.940 ;
        RECT  4.400 0.870 4.860 0.940 ;
        RECT  4.365 0.460 4.400 0.940 ;
        RECT  4.330 0.185 4.365 0.940 ;
        RECT  4.295 0.185 4.330 0.530 ;
        RECT  4.260 0.870 4.330 0.940 ;
        RECT  4.020 0.460 4.295 0.530 ;
        RECT  4.080 0.635 4.255 0.755 ;
        RECT  4.010 0.635 4.080 1.050 ;
        RECT  3.930 0.635 4.010 0.705 ;
        RECT  3.700 0.980 4.010 1.050 ;
        RECT  3.790 0.815 3.940 0.885 ;
        RECT  3.860 0.185 3.930 0.705 ;
        RECT  3.730 0.185 3.860 0.255 ;
        RECT  3.720 0.440 3.790 0.885 ;
        RECT  3.625 0.220 3.650 0.800 ;
        RECT  3.580 0.220 3.625 1.050 ;
        RECT  3.565 0.220 3.580 0.340 ;
        RECT  3.555 0.730 3.580 1.050 ;
        RECT  3.315 0.730 3.555 0.800 ;
        RECT  3.440 0.510 3.510 0.640 ;
        RECT  3.075 0.510 3.440 0.580 ;
        RECT  3.245 0.680 3.315 0.800 ;
        RECT  3.070 0.300 3.075 0.580 ;
        RECT  3.000 0.300 3.070 0.960 ;
        RECT  2.860 0.205 2.930 0.935 ;
        RECT  2.165 0.205 2.860 0.275 ;
        RECT  2.790 0.865 2.860 1.040 ;
        RECT  2.250 0.970 2.790 1.040 ;
        RECT  2.705 0.355 2.775 0.765 ;
        RECT  2.610 0.355 2.705 0.425 ;
        RECT  2.635 0.695 2.705 0.850 ;
        RECT  2.540 0.545 2.625 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.250 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.095 0.205 2.165 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSND2BWP

MACRO SDFKCSND4BWP
    CLASS CORE ;
    FOREIGN SDFKCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.335 0.185 6.345 0.465 ;
        RECT  6.335 0.765 6.345 1.065 ;
        RECT  6.275 0.185 6.335 1.065 ;
        RECT  6.125 0.355 6.275 0.905 ;
        RECT  5.985 0.355 6.125 0.465 ;
        RECT  5.985 0.765 6.125 0.905 ;
        RECT  5.915 0.185 5.985 0.465 ;
        RECT  5.915 0.765 5.985 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.700 5.650 0.800 ;
        RECT  5.555 0.185 5.625 0.485 ;
        RECT  5.495 0.355 5.555 0.485 ;
        RECT  5.285 0.355 5.495 0.800 ;
        RECT  5.265 0.355 5.285 0.485 ;
        RECT  5.170 0.700 5.285 0.800 ;
        RECT  5.195 0.185 5.265 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 -0.115 6.580 0.115 ;
        RECT  6.450 -0.115 6.530 0.465 ;
        RECT  6.190 -0.115 6.450 0.115 ;
        RECT  6.070 -0.115 6.190 0.275 ;
        RECT  5.805 -0.115 6.070 0.115 ;
        RECT  5.735 -0.115 5.805 0.465 ;
        RECT  5.470 -0.115 5.735 0.115 ;
        RECT  5.350 -0.115 5.470 0.275 ;
        RECT  5.085 -0.115 5.350 0.115 ;
        RECT  5.015 -0.115 5.085 0.305 ;
        RECT  4.725 -0.115 5.015 0.115 ;
        RECT  4.655 -0.115 4.725 0.320 ;
        RECT  3.805 -0.115 4.655 0.115 ;
        RECT  3.735 -0.115 3.805 0.460 ;
        RECT  3.445 -0.115 3.735 0.115 ;
        RECT  3.375 -0.115 3.445 0.400 ;
        RECT  2.540 -0.115 3.375 0.115 ;
        RECT  2.420 -0.115 2.540 0.135 ;
        RECT  1.990 -0.115 2.420 0.115 ;
        RECT  1.870 -0.115 1.990 0.265 ;
        RECT  1.600 -0.115 1.870 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.580 1.375 ;
        RECT  6.450 0.675 6.530 1.375 ;
        RECT  6.165 1.145 6.450 1.375 ;
        RECT  6.095 0.975 6.165 1.375 ;
        RECT  5.830 1.145 6.095 1.375 ;
        RECT  5.710 1.010 5.830 1.375 ;
        RECT  5.470 1.145 5.710 1.375 ;
        RECT  5.350 1.010 5.470 1.375 ;
        RECT  5.110 1.145 5.350 1.375 ;
        RECT  4.990 1.010 5.110 1.375 ;
        RECT  4.730 1.145 4.990 1.375 ;
        RECT  4.660 0.950 4.730 1.375 ;
        RECT  3.820 1.145 4.660 1.375 ;
        RECT  3.720 0.860 3.820 1.375 ;
        RECT  3.445 1.145 3.720 1.375 ;
        RECT  3.375 0.860 3.445 1.375 ;
        RECT  2.560 1.145 3.375 1.375 ;
        RECT  2.440 1.110 2.560 1.375 ;
        RECT  2.000 1.145 2.440 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.985 0.355 6.055 0.465 ;
        RECT  5.985 0.765 6.055 0.905 ;
        RECT  5.915 0.185 5.985 0.465 ;
        RECT  5.915 0.765 5.985 1.065 ;
        RECT  5.565 0.700 5.650 0.800 ;
        RECT  5.565 0.185 5.625 0.485 ;
        RECT  5.195 0.185 5.215 0.485 ;
        RECT  5.170 0.700 5.215 0.800 ;
        RECT  5.810 0.545 5.950 0.615 ;
        RECT  5.740 0.545 5.810 0.940 ;
        RECT  5.060 0.870 5.740 0.940 ;
        RECT  4.990 0.435 5.060 0.940 ;
        RECT  4.905 0.435 4.990 0.505 ;
        RECT  4.905 0.870 4.990 0.940 ;
        RECT  4.835 0.200 4.905 0.505 ;
        RECT  4.835 0.870 4.905 1.010 ;
        RECT  4.590 0.585 4.870 0.655 ;
        RECT  4.560 0.435 4.835 0.505 ;
        RECT  4.520 0.585 4.590 1.055 ;
        RECT  4.480 0.585 4.520 0.655 ;
        RECT  3.985 0.985 4.520 1.055 ;
        RECT  4.410 0.270 4.480 0.655 ;
        RECT  4.360 0.780 4.450 0.910 ;
        RECT  4.365 0.270 4.410 0.340 ;
        RECT  4.295 0.195 4.365 0.340 ;
        RECT  4.310 0.780 4.360 0.850 ;
        RECT  4.240 0.485 4.310 0.850 ;
        RECT  3.980 0.195 4.295 0.265 ;
        RECT  4.190 0.485 4.240 0.555 ;
        RECT  4.120 0.335 4.190 0.405 ;
        RECT  4.120 0.710 4.165 0.890 ;
        RECT  4.095 0.335 4.120 0.890 ;
        RECT  4.050 0.335 4.095 0.780 ;
        RECT  3.665 0.710 4.050 0.780 ;
        RECT  3.915 0.850 3.985 1.055 ;
        RECT  3.910 0.195 3.980 0.350 ;
        RECT  3.625 0.335 3.665 0.780 ;
        RECT  3.595 0.335 3.625 0.980 ;
        RECT  3.530 0.335 3.595 0.405 ;
        RECT  3.555 0.710 3.595 0.980 ;
        RECT  3.335 0.710 3.555 0.780 ;
        RECT  3.445 0.510 3.515 0.640 ;
        RECT  3.085 0.510 3.445 0.580 ;
        RECT  3.265 0.660 3.335 0.780 ;
        RECT  3.075 0.510 3.085 0.980 ;
        RECT  3.005 0.280 3.075 0.980 ;
        RECT  2.880 0.205 2.935 0.935 ;
        RECT  2.865 0.205 2.880 1.040 ;
        RECT  2.145 0.205 2.865 0.275 ;
        RECT  2.810 0.865 2.865 1.040 ;
        RECT  2.250 0.970 2.810 1.040 ;
        RECT  2.725 0.355 2.795 0.765 ;
        RECT  2.610 0.355 2.725 0.425 ;
        RECT  2.655 0.695 2.725 0.850 ;
        RECT  2.540 0.545 2.640 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.230 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.075 0.205 2.145 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSND4BWP

MACRO SDFKCSNQD0BWP
    CLASS CORE ;
    FOREIGN SDFKCSNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.635 0.945 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.225 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.630 1.385 0.905 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0096 ;
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.195 4.585 1.045 ;
        RECT  4.495 0.195 4.515 0.415 ;
        RECT  4.495 0.905 4.515 1.045 ;
        RECT  4.265 0.345 4.495 0.415 ;
        RECT  4.195 0.345 4.265 0.610 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0152 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.415 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.495 2.575 0.640 ;
        RECT  2.410 0.495 2.485 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.525 0.240 0.605 ;
        RECT  0.105 0.495 0.125 0.605 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.255 ;
        RECT  3.605 -0.115 4.280 0.115 ;
        RECT  3.535 -0.115 3.605 0.420 ;
        RECT  2.680 -0.115 3.535 0.115 ;
        RECT  2.560 -0.115 2.680 0.125 ;
        RECT  2.180 -0.115 2.560 0.115 ;
        RECT  2.060 -0.115 2.180 0.125 ;
        RECT  1.405 -0.115 2.060 0.115 ;
        RECT  1.335 -0.115 1.405 0.400 ;
        RECT  1.040 -0.115 1.335 0.115 ;
        RECT  0.920 -0.115 1.040 0.125 ;
        RECT  0.125 -0.115 0.920 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.390 1.145 4.620 1.375 ;
        RECT  4.320 0.915 4.390 1.375 ;
        RECT  3.620 1.145 4.320 1.375 ;
        RECT  3.500 0.870 3.620 1.375 ;
        RECT  2.680 1.145 3.500 1.375 ;
        RECT  2.560 1.130 2.680 1.375 ;
        RECT  2.180 1.145 2.560 1.375 ;
        RECT  2.060 1.135 2.180 1.375 ;
        RECT  1.400 1.145 2.060 1.375 ;
        RECT  1.280 1.135 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.135 1.100 1.375 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.620 1.135 0.740 1.375 ;
        RECT  0.125 1.145 0.620 1.375 ;
        RECT  0.055 0.970 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.375 0.510 4.445 0.750 ;
        RECT  4.250 0.680 4.375 0.750 ;
        RECT  4.180 0.680 4.250 1.060 ;
        RECT  4.090 0.680 4.180 0.750 ;
        RECT  3.860 0.990 4.180 1.060 ;
        RECT  3.950 0.830 4.100 0.900 ;
        RECT  4.020 0.195 4.090 0.750 ;
        RECT  3.890 0.195 4.020 0.265 ;
        RECT  3.880 0.430 3.950 0.900 ;
        RECT  3.785 0.220 3.810 0.800 ;
        RECT  3.740 0.220 3.785 1.050 ;
        RECT  3.725 0.220 3.740 0.340 ;
        RECT  3.715 0.730 3.740 1.050 ;
        RECT  3.495 0.730 3.715 0.800 ;
        RECT  3.600 0.510 3.670 0.640 ;
        RECT  3.235 0.510 3.600 0.580 ;
        RECT  3.425 0.675 3.495 0.800 ;
        RECT  3.225 0.300 3.235 0.580 ;
        RECT  3.155 0.300 3.225 0.960 ;
        RECT  1.765 0.195 3.080 0.265 ;
        RECT  2.975 0.840 3.045 1.060 ;
        RECT  1.660 0.990 2.975 1.060 ;
        RECT  2.870 0.340 2.935 0.765 ;
        RECT  2.865 0.340 2.870 0.850 ;
        RECT  2.795 0.340 2.865 0.460 ;
        RECT  2.795 0.695 2.865 0.850 ;
        RECT  2.715 0.520 2.750 0.640 ;
        RECT  2.645 0.355 2.715 0.915 ;
        RECT  2.410 0.355 2.645 0.425 ;
        RECT  2.410 0.845 2.645 0.915 ;
        RECT  2.025 0.335 2.330 0.405 ;
        RECT  2.025 0.845 2.330 0.915 ;
        RECT  1.955 0.335 2.025 0.915 ;
        RECT  1.775 0.475 1.845 0.760 ;
        RECT  1.225 0.475 1.775 0.545 ;
        RECT  1.695 0.195 1.765 0.400 ;
        RECT  1.560 0.665 1.690 0.735 ;
        RECT  1.490 0.665 1.560 1.065 ;
        RECT  1.085 0.995 1.490 1.065 ;
        RECT  1.155 0.210 1.225 0.910 ;
        RECT  1.015 0.195 1.085 1.065 ;
        RECT  0.400 0.195 1.015 0.265 ;
        RECT  0.400 0.995 1.015 1.065 ;
        RECT  0.605 0.840 0.900 0.910 ;
        RECT  0.795 0.350 0.865 0.555 ;
        RECT  0.605 0.485 0.795 0.555 ;
        RECT  0.210 0.335 0.710 0.405 ;
        RECT  0.535 0.485 0.605 0.910 ;
        RECT  0.245 0.840 0.535 0.910 ;
        RECT  0.175 0.725 0.245 0.910 ;
    END
END SDFKCSNQD0BWP

MACRO SDFKCSNQD1BWP
    CLASS CORE ;
    FOREIGN SDFKCSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.195 4.725 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 -0.115 4.760 0.115 ;
        RECT  4.455 -0.115 4.525 0.305 ;
        RECT  4.165 -0.115 4.455 0.115 ;
        RECT  4.095 -0.115 4.165 0.285 ;
        RECT  3.425 -0.115 4.095 0.115 ;
        RECT  3.355 -0.115 3.425 0.420 ;
        RECT  2.520 -0.115 3.355 0.115 ;
        RECT  2.400 -0.115 2.520 0.135 ;
        RECT  1.990 -0.115 2.400 0.115 ;
        RECT  1.870 -0.115 1.990 0.265 ;
        RECT  1.600 -0.115 1.870 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.145 4.760 1.375 ;
        RECT  4.455 0.905 4.525 1.375 ;
        RECT  4.170 1.145 4.455 1.375 ;
        RECT  4.100 0.955 4.170 1.375 ;
        RECT  3.450 1.145 4.100 1.375 ;
        RECT  3.330 0.870 3.450 1.375 ;
        RECT  2.540 1.145 3.330 1.375 ;
        RECT  2.420 1.110 2.540 1.375 ;
        RECT  2.000 1.145 2.420 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.485 0.395 4.555 0.820 ;
        RECT  4.345 0.395 4.485 0.465 ;
        RECT  4.345 0.750 4.485 0.820 ;
        RECT  4.030 0.545 4.390 0.615 ;
        RECT  4.275 0.185 4.345 0.465 ;
        RECT  4.275 0.750 4.345 1.075 ;
        RECT  4.000 0.395 4.275 0.465 ;
        RECT  3.960 0.545 4.030 1.060 ;
        RECT  3.910 0.545 3.960 0.615 ;
        RECT  3.690 0.990 3.960 1.060 ;
        RECT  3.840 0.195 3.910 0.615 ;
        RECT  3.770 0.800 3.890 0.920 ;
        RECT  3.710 0.195 3.840 0.265 ;
        RECT  3.700 0.440 3.770 0.920 ;
        RECT  3.605 0.220 3.630 0.800 ;
        RECT  3.560 0.220 3.605 1.050 ;
        RECT  3.545 0.220 3.560 0.340 ;
        RECT  3.535 0.730 3.560 1.050 ;
        RECT  3.315 0.730 3.535 0.800 ;
        RECT  3.420 0.510 3.490 0.640 ;
        RECT  3.070 0.510 3.420 0.580 ;
        RECT  3.245 0.680 3.315 0.800 ;
        RECT  3.055 0.510 3.070 0.960 ;
        RECT  2.985 0.300 3.055 0.960 ;
        RECT  2.860 0.205 2.915 0.935 ;
        RECT  2.845 0.205 2.860 1.040 ;
        RECT  2.145 0.205 2.845 0.275 ;
        RECT  2.790 0.865 2.845 1.040 ;
        RECT  2.250 0.970 2.790 1.040 ;
        RECT  2.705 0.355 2.775 0.765 ;
        RECT  2.590 0.355 2.705 0.425 ;
        RECT  2.635 0.695 2.705 0.850 ;
        RECT  2.510 0.545 2.625 0.615 ;
        RECT  2.440 0.355 2.510 0.855 ;
        RECT  2.230 0.355 2.440 0.425 ;
        RECT  2.275 0.735 2.440 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.075 0.205 2.145 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSNQD1BWP

MACRO SDFKCSNQD2BWP
    CLASS CORE ;
    FOREIGN SDFKCSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.805 0.355 4.865 0.805 ;
        RECT  4.795 0.185 4.805 1.035 ;
        RECT  4.735 0.185 4.795 0.465 ;
        RECT  4.735 0.735 4.795 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.300 ;
        RECT  4.625 -0.115 4.910 0.115 ;
        RECT  4.555 -0.115 4.625 0.305 ;
        RECT  4.245 -0.115 4.555 0.115 ;
        RECT  4.175 -0.115 4.245 0.290 ;
        RECT  3.485 -0.115 4.175 0.115 ;
        RECT  3.415 -0.115 3.485 0.420 ;
        RECT  2.560 -0.115 3.415 0.115 ;
        RECT  2.440 -0.115 2.560 0.135 ;
        RECT  2.000 -0.115 2.440 0.115 ;
        RECT  1.880 -0.115 2.000 0.265 ;
        RECT  1.600 -0.115 1.880 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.905 4.990 1.375 ;
        RECT  4.625 1.145 4.910 1.375 ;
        RECT  4.555 0.905 4.625 1.375 ;
        RECT  4.260 1.145 4.555 1.375 ;
        RECT  4.140 1.120 4.260 1.375 ;
        RECT  3.500 1.145 4.140 1.375 ;
        RECT  3.380 0.870 3.500 1.375 ;
        RECT  2.560 1.145 3.380 1.375 ;
        RECT  2.440 1.110 2.560 1.375 ;
        RECT  2.000 1.145 2.440 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.395 4.655 0.835 ;
        RECT  4.425 0.395 4.585 0.465 ;
        RECT  4.425 0.765 4.585 0.835 ;
        RECT  4.140 0.545 4.460 0.615 ;
        RECT  4.355 0.190 4.425 0.465 ;
        RECT  4.355 0.765 4.425 1.070 ;
        RECT  4.080 0.395 4.355 0.465 ;
        RECT  4.070 0.545 4.140 1.050 ;
        RECT  3.970 0.545 4.070 0.615 ;
        RECT  3.740 0.980 4.070 1.050 ;
        RECT  3.830 0.815 3.980 0.885 ;
        RECT  3.900 0.185 3.970 0.615 ;
        RECT  3.770 0.185 3.900 0.255 ;
        RECT  3.760 0.440 3.830 0.885 ;
        RECT  3.665 0.220 3.690 0.800 ;
        RECT  3.620 0.220 3.665 1.050 ;
        RECT  3.605 0.220 3.620 0.340 ;
        RECT  3.595 0.730 3.620 1.050 ;
        RECT  3.355 0.730 3.595 0.800 ;
        RECT  3.480 0.510 3.550 0.640 ;
        RECT  3.095 0.510 3.480 0.580 ;
        RECT  3.285 0.680 3.355 0.800 ;
        RECT  3.090 0.300 3.095 0.580 ;
        RECT  3.020 0.300 3.090 0.960 ;
        RECT  2.880 0.205 2.950 0.935 ;
        RECT  2.165 0.205 2.880 0.275 ;
        RECT  2.810 0.865 2.880 1.040 ;
        RECT  2.250 0.970 2.810 1.040 ;
        RECT  2.725 0.355 2.795 0.765 ;
        RECT  2.630 0.355 2.725 0.425 ;
        RECT  2.655 0.695 2.725 0.850 ;
        RECT  2.540 0.545 2.640 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.250 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.095 0.205 2.165 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSNQD2BWP

MACRO SDFKCSNQD4BWP
    CLASS CORE ;
    FOREIGN SDFKCSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.755 0.220 0.825 ;
        RECT  0.035 0.495 0.125 0.825 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.500 1.555 0.650 ;
        RECT  1.365 0.500 1.485 0.570 ;
        RECT  1.295 0.215 1.365 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 1.925 0.650 ;
        RECT  1.820 0.520 1.855 0.650 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.185 5.645 0.465 ;
        RECT  5.635 0.765 5.645 1.065 ;
        RECT  5.575 0.185 5.635 1.065 ;
        RECT  5.425 0.355 5.575 0.905 ;
        RECT  5.290 0.355 5.425 0.465 ;
        RECT  5.290 0.765 5.425 0.905 ;
        RECT  5.220 0.185 5.290 0.465 ;
        RECT  5.220 0.765 5.290 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0184 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.755 0.580 0.825 ;
        RECT  0.455 0.755 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.540 2.310 0.620 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0160 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.865 ;
        RECT  0.415 0.475 0.875 0.545 ;
        RECT  0.690 0.795 0.875 0.865 ;
        RECT  0.345 0.410 0.415 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.825 -0.115 5.880 0.115 ;
        RECT  5.755 -0.115 5.825 0.465 ;
        RECT  5.490 -0.115 5.755 0.115 ;
        RECT  5.370 -0.115 5.490 0.275 ;
        RECT  5.105 -0.115 5.370 0.115 ;
        RECT  5.035 -0.115 5.105 0.305 ;
        RECT  4.725 -0.115 5.035 0.115 ;
        RECT  4.655 -0.115 4.725 0.320 ;
        RECT  3.805 -0.115 4.655 0.115 ;
        RECT  3.735 -0.115 3.805 0.460 ;
        RECT  3.445 -0.115 3.735 0.115 ;
        RECT  3.375 -0.115 3.445 0.400 ;
        RECT  2.540 -0.115 3.375 0.115 ;
        RECT  2.420 -0.115 2.540 0.135 ;
        RECT  1.990 -0.115 2.420 0.115 ;
        RECT  1.870 -0.115 1.990 0.265 ;
        RECT  1.600 -0.115 1.870 0.115 ;
        RECT  1.530 -0.115 1.600 0.430 ;
        RECT  0.305 -0.115 1.530 0.115 ;
        RECT  0.235 -0.115 0.305 0.285 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.825 1.145 5.880 1.375 ;
        RECT  5.755 0.675 5.825 1.375 ;
        RECT  5.465 1.145 5.755 1.375 ;
        RECT  5.395 0.975 5.465 1.375 ;
        RECT  5.105 1.145 5.395 1.375 ;
        RECT  5.035 0.905 5.105 1.375 ;
        RECT  4.730 1.145 5.035 1.375 ;
        RECT  4.660 0.940 4.730 1.375 ;
        RECT  3.820 1.145 4.660 1.375 ;
        RECT  3.720 0.860 3.820 1.375 ;
        RECT  3.445 1.145 3.720 1.375 ;
        RECT  3.375 0.860 3.445 1.375 ;
        RECT  2.560 1.145 3.375 1.375 ;
        RECT  2.440 1.110 2.560 1.375 ;
        RECT  2.000 1.145 2.440 1.375 ;
        RECT  1.880 1.110 2.000 1.375 ;
        RECT  1.660 1.145 1.880 1.375 ;
        RECT  1.540 1.040 1.660 1.375 ;
        RECT  0.910 1.145 1.540 1.375 ;
        RECT  0.790 1.110 0.910 1.375 ;
        RECT  0.330 1.145 0.790 1.375 ;
        RECT  0.210 1.035 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.290 0.355 5.355 0.465 ;
        RECT  5.290 0.765 5.355 0.905 ;
        RECT  5.220 0.185 5.290 0.465 ;
        RECT  5.220 0.765 5.290 1.065 ;
        RECT  5.080 0.395 5.150 0.835 ;
        RECT  4.905 0.395 5.080 0.465 ;
        RECT  4.905 0.765 5.080 0.835 ;
        RECT  4.590 0.545 5.010 0.615 ;
        RECT  4.835 0.200 4.905 0.465 ;
        RECT  4.835 0.765 4.905 1.070 ;
        RECT  4.560 0.395 4.835 0.465 ;
        RECT  4.520 0.545 4.590 1.055 ;
        RECT  4.480 0.545 4.520 0.615 ;
        RECT  3.985 0.985 4.520 1.055 ;
        RECT  4.410 0.270 4.480 0.615 ;
        RECT  4.360 0.780 4.450 0.910 ;
        RECT  4.365 0.270 4.410 0.340 ;
        RECT  4.295 0.195 4.365 0.340 ;
        RECT  4.310 0.780 4.360 0.850 ;
        RECT  4.240 0.485 4.310 0.850 ;
        RECT  3.980 0.195 4.295 0.265 ;
        RECT  4.190 0.485 4.240 0.555 ;
        RECT  4.120 0.335 4.190 0.405 ;
        RECT  4.120 0.710 4.165 0.890 ;
        RECT  4.095 0.335 4.120 0.890 ;
        RECT  4.050 0.335 4.095 0.780 ;
        RECT  3.665 0.710 4.050 0.780 ;
        RECT  3.915 0.850 3.985 1.055 ;
        RECT  3.910 0.195 3.980 0.350 ;
        RECT  3.625 0.335 3.665 0.780 ;
        RECT  3.595 0.335 3.625 0.980 ;
        RECT  3.530 0.335 3.595 0.405 ;
        RECT  3.555 0.710 3.595 0.980 ;
        RECT  3.335 0.710 3.555 0.780 ;
        RECT  3.445 0.510 3.515 0.640 ;
        RECT  3.085 0.510 3.445 0.580 ;
        RECT  3.265 0.660 3.335 0.780 ;
        RECT  3.075 0.510 3.085 0.980 ;
        RECT  3.005 0.280 3.075 0.980 ;
        RECT  2.880 0.205 2.935 0.935 ;
        RECT  2.865 0.205 2.880 1.040 ;
        RECT  2.145 0.205 2.865 0.275 ;
        RECT  2.810 0.865 2.865 1.040 ;
        RECT  2.250 0.970 2.810 1.040 ;
        RECT  2.725 0.355 2.795 0.765 ;
        RECT  2.610 0.355 2.725 0.425 ;
        RECT  2.655 0.695 2.725 0.850 ;
        RECT  2.540 0.545 2.640 0.615 ;
        RECT  2.470 0.355 2.540 0.855 ;
        RECT  2.230 0.355 2.470 0.425 ;
        RECT  2.275 0.735 2.470 0.855 ;
        RECT  2.180 0.970 2.250 1.060 ;
        RECT  2.070 0.990 2.180 1.060 ;
        RECT  2.075 0.205 2.145 0.410 ;
        RECT  1.995 0.510 2.065 0.910 ;
        RECT  1.965 0.840 1.995 0.910 ;
        RECT  1.905 0.840 1.965 0.930 ;
        RECT  1.260 0.860 1.905 0.930 ;
        RECT  1.750 0.720 1.840 0.790 ;
        RECT  1.750 0.190 1.785 0.310 ;
        RECT  1.680 0.190 1.750 0.790 ;
        RECT  1.375 0.720 1.680 0.790 ;
        RECT  1.305 0.640 1.375 0.790 ;
        RECT  1.225 0.860 1.260 0.960 ;
        RECT  1.155 0.195 1.225 0.960 ;
        RECT  1.045 0.335 1.085 1.060 ;
        RECT  1.015 0.235 1.045 1.060 ;
        RECT  0.975 0.235 1.015 0.405 ;
        RECT  0.995 0.935 1.015 1.060 ;
        RECT  0.670 0.935 0.995 1.005 ;
        RECT  0.580 0.335 0.975 0.405 ;
        RECT  0.390 0.195 0.890 0.265 ;
        RECT  0.375 0.615 0.790 0.685 ;
        RECT  0.600 0.935 0.670 1.060 ;
        RECT  0.305 0.615 0.375 0.965 ;
        RECT  0.265 0.615 0.305 0.685 ;
        RECT  0.125 0.895 0.305 0.965 ;
        RECT  0.195 0.355 0.265 0.685 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.895 0.125 1.070 ;
    END
END SDFKCSNQD4BWP

MACRO SDFKSND0BWP
    CLASS CORE ;
    FOREIGN SDFKSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.335 4.725 0.905 ;
        RECT  4.635 0.335 4.655 0.455 ;
        RECT  4.640 0.765 4.655 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.215 4.445 0.485 ;
        RECT  4.330 0.360 4.375 0.485 ;
        RECT  4.260 0.360 4.330 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.635 0.735 0.780 ;
        RECT  0.595 0.635 0.665 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.145 ;
        RECT  3.965 -0.115 4.420 0.115 ;
        RECT  3.895 -0.115 3.965 0.285 ;
        RECT  3.225 -0.115 3.895 0.115 ;
        RECT  3.155 -0.115 3.225 0.420 ;
        RECT  2.320 -0.115 3.155 0.115 ;
        RECT  2.200 -0.115 2.320 0.135 ;
        RECT  1.790 -0.115 2.200 0.115 ;
        RECT  1.670 -0.115 1.790 0.275 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 1.145 4.760 1.375 ;
        RECT  4.445 1.010 4.515 1.375 ;
        RECT  3.970 1.145 4.445 1.375 ;
        RECT  3.900 0.955 3.970 1.375 ;
        RECT  3.250 1.145 3.900 1.375 ;
        RECT  3.130 0.870 3.250 1.375 ;
        RECT  2.340 1.145 3.130 1.375 ;
        RECT  2.220 1.115 2.340 1.375 ;
        RECT  1.800 1.145 2.220 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.975 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.560 0.520 4.580 0.675 ;
        RECT  4.510 0.520 4.560 0.940 ;
        RECT  4.490 0.605 4.510 0.940 ;
        RECT  4.180 0.870 4.490 0.940 ;
        RECT  4.145 0.395 4.180 0.940 ;
        RECT  4.110 0.185 4.145 1.075 ;
        RECT  4.075 0.185 4.110 0.465 ;
        RECT  4.075 0.870 4.110 1.075 ;
        RECT  3.800 0.395 4.075 0.465 ;
        RECT  3.830 0.600 4.035 0.720 ;
        RECT  3.760 0.600 3.830 1.060 ;
        RECT  3.710 0.600 3.760 0.720 ;
        RECT  3.490 0.990 3.760 1.060 ;
        RECT  3.640 0.195 3.710 0.720 ;
        RECT  3.570 0.800 3.690 0.920 ;
        RECT  3.510 0.195 3.640 0.265 ;
        RECT  3.500 0.440 3.570 0.920 ;
        RECT  3.405 0.220 3.430 0.800 ;
        RECT  3.360 0.220 3.405 1.050 ;
        RECT  3.345 0.220 3.360 0.340 ;
        RECT  3.335 0.730 3.360 1.050 ;
        RECT  3.115 0.730 3.335 0.800 ;
        RECT  3.220 0.510 3.290 0.640 ;
        RECT  2.870 0.510 3.220 0.580 ;
        RECT  3.045 0.680 3.115 0.800 ;
        RECT  2.855 0.510 2.870 0.960 ;
        RECT  2.785 0.300 2.855 0.960 ;
        RECT  2.660 0.205 2.715 0.935 ;
        RECT  2.645 0.205 2.660 1.045 ;
        RECT  1.945 0.205 2.645 0.275 ;
        RECT  2.590 0.865 2.645 1.045 ;
        RECT  2.080 0.975 2.590 1.045 ;
        RECT  2.505 0.345 2.575 0.765 ;
        RECT  2.415 0.345 2.505 0.465 ;
        RECT  2.435 0.695 2.505 0.850 ;
        RECT  2.345 0.545 2.420 0.615 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.250 1.025 1.050 ;
        RECT  0.810 0.280 0.880 1.040 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.900 0.810 1.040 ;
        RECT  0.485 0.995 0.700 1.065 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.065 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.905 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.835 0.260 0.905 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.835 0.125 1.025 ;
    END
END SDFKSND0BWP

MACRO SDFKSND1BWP
    CLASS CORE ;
    FOREIGN SDFKSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.045 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.735 4.655 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.330 0.215 4.445 0.485 ;
        RECT  4.260 0.215 4.330 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.145 ;
        RECT  3.965 -0.115 4.420 0.115 ;
        RECT  3.895 -0.115 3.965 0.270 ;
        RECT  3.225 -0.115 3.895 0.115 ;
        RECT  3.155 -0.115 3.225 0.420 ;
        RECT  2.320 -0.115 3.155 0.115 ;
        RECT  2.200 -0.115 2.320 0.135 ;
        RECT  1.790 -0.115 2.200 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.760 1.375 ;
        RECT  4.420 1.025 4.540 1.375 ;
        RECT  3.970 1.145 4.420 1.375 ;
        RECT  3.900 0.955 3.970 1.375 ;
        RECT  3.250 1.145 3.900 1.375 ;
        RECT  3.130 0.870 3.250 1.375 ;
        RECT  2.340 1.145 3.130 1.375 ;
        RECT  2.220 1.115 2.340 1.375 ;
        RECT  1.800 1.145 2.220 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.560 0.515 4.580 0.665 ;
        RECT  4.510 0.515 4.560 0.940 ;
        RECT  4.490 0.595 4.510 0.940 ;
        RECT  4.180 0.870 4.490 0.940 ;
        RECT  4.145 0.395 4.180 0.940 ;
        RECT  4.110 0.185 4.145 1.075 ;
        RECT  4.075 0.185 4.110 0.465 ;
        RECT  4.075 0.870 4.110 1.075 ;
        RECT  3.800 0.395 4.075 0.465 ;
        RECT  3.830 0.600 4.035 0.720 ;
        RECT  3.760 0.600 3.830 1.060 ;
        RECT  3.710 0.600 3.760 0.720 ;
        RECT  3.490 0.990 3.760 1.060 ;
        RECT  3.640 0.195 3.710 0.720 ;
        RECT  3.570 0.800 3.690 0.920 ;
        RECT  3.510 0.195 3.640 0.265 ;
        RECT  3.500 0.440 3.570 0.920 ;
        RECT  3.405 0.220 3.430 0.800 ;
        RECT  3.360 0.220 3.405 1.050 ;
        RECT  3.345 0.220 3.360 0.340 ;
        RECT  3.335 0.730 3.360 1.050 ;
        RECT  3.115 0.730 3.335 0.800 ;
        RECT  3.220 0.510 3.290 0.640 ;
        RECT  2.870 0.510 3.220 0.580 ;
        RECT  3.045 0.680 3.115 0.800 ;
        RECT  2.855 0.510 2.870 0.960 ;
        RECT  2.785 0.300 2.855 0.960 ;
        RECT  2.660 0.205 2.715 0.935 ;
        RECT  2.645 0.205 2.660 1.045 ;
        RECT  1.945 0.205 2.645 0.275 ;
        RECT  2.590 0.865 2.645 1.045 ;
        RECT  2.080 0.975 2.590 1.045 ;
        RECT  2.505 0.345 2.575 0.765 ;
        RECT  2.415 0.345 2.505 0.465 ;
        RECT  2.435 0.695 2.505 0.890 ;
        RECT  2.345 0.545 2.420 0.615 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSND1BWP

MACRO SDFKSND2BWP
    CLASS CORE ;
    FOREIGN SDFKSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.355 5.005 0.805 ;
        RECT  4.935 0.185 4.945 1.035 ;
        RECT  4.875 0.185 4.935 0.465 ;
        RECT  4.875 0.735 4.935 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.195 4.585 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.300 ;
        RECT  4.765 -0.115 5.050 0.115 ;
        RECT  4.695 -0.115 4.765 0.465 ;
        RECT  4.405 -0.115 4.695 0.115 ;
        RECT  4.335 -0.115 4.405 0.315 ;
        RECT  4.015 -0.115 4.335 0.115 ;
        RECT  3.945 -0.115 4.015 0.270 ;
        RECT  3.265 -0.115 3.945 0.115 ;
        RECT  3.195 -0.115 3.265 0.420 ;
        RECT  2.340 -0.115 3.195 0.115 ;
        RECT  2.220 -0.115 2.340 0.135 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.145 5.180 1.375 ;
        RECT  5.050 0.905 5.130 1.375 ;
        RECT  4.790 1.145 5.050 1.375 ;
        RECT  4.670 1.010 4.790 1.375 ;
        RECT  4.430 1.145 4.670 1.375 ;
        RECT  4.310 1.010 4.430 1.375 ;
        RECT  4.020 1.145 4.310 1.375 ;
        RECT  3.950 0.955 4.020 1.375 ;
        RECT  3.290 1.145 3.950 1.375 ;
        RECT  3.170 0.870 3.290 1.375 ;
        RECT  2.360 1.145 3.170 1.375 ;
        RECT  2.240 1.115 2.360 1.375 ;
        RECT  1.800 1.145 2.240 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.790 0.545 4.860 0.615 ;
        RECT  4.720 0.545 4.790 0.940 ;
        RECT  4.410 0.870 4.720 0.940 ;
        RECT  4.340 0.395 4.410 0.940 ;
        RECT  4.205 0.395 4.340 0.465 ;
        RECT  4.205 0.870 4.340 0.940 ;
        RECT  3.870 0.545 4.240 0.615 ;
        RECT  4.135 0.185 4.205 0.465 ;
        RECT  4.135 0.870 4.205 1.045 ;
        RECT  3.840 0.395 4.135 0.465 ;
        RECT  3.800 0.545 3.870 1.060 ;
        RECT  3.750 0.545 3.800 0.615 ;
        RECT  3.530 0.990 3.800 1.060 ;
        RECT  3.680 0.195 3.750 0.615 ;
        RECT  3.610 0.800 3.730 0.920 ;
        RECT  3.550 0.195 3.680 0.265 ;
        RECT  3.540 0.440 3.610 0.920 ;
        RECT  3.445 0.220 3.470 0.800 ;
        RECT  3.400 0.220 3.445 1.050 ;
        RECT  3.385 0.220 3.400 0.340 ;
        RECT  3.375 0.730 3.400 1.050 ;
        RECT  3.155 0.730 3.375 0.800 ;
        RECT  3.260 0.510 3.330 0.640 ;
        RECT  2.890 0.510 3.260 0.580 ;
        RECT  3.085 0.680 3.155 0.800 ;
        RECT  2.875 0.510 2.890 0.960 ;
        RECT  2.805 0.300 2.875 0.960 ;
        RECT  2.680 0.205 2.735 0.935 ;
        RECT  2.665 0.205 2.680 1.045 ;
        RECT  1.945 0.205 2.665 0.275 ;
        RECT  2.610 0.865 2.665 1.045 ;
        RECT  2.080 0.975 2.610 1.045 ;
        RECT  2.525 0.345 2.595 0.765 ;
        RECT  2.435 0.345 2.525 0.465 ;
        RECT  2.455 0.695 2.525 0.890 ;
        RECT  2.345 0.545 2.440 0.620 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSND2BWP

MACRO SDFKSND4BWP
    CLASS CORE ;
    FOREIGN SDFKSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.195 0.185 6.205 0.465 ;
        RECT  6.195 0.765 6.205 1.065 ;
        RECT  6.135 0.185 6.195 1.065 ;
        RECT  5.985 0.355 6.135 0.905 ;
        RECT  5.845 0.355 5.985 0.465 ;
        RECT  5.845 0.765 5.985 0.905 ;
        RECT  5.775 0.185 5.845 0.465 ;
        RECT  5.775 0.765 5.845 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.355 0.700 5.510 0.800 ;
        RECT  5.415 0.185 5.485 0.485 ;
        RECT  5.355 0.355 5.415 0.485 ;
        RECT  5.145 0.355 5.355 0.800 ;
        RECT  5.125 0.355 5.145 0.485 ;
        RECT  5.030 0.700 5.145 0.800 ;
        RECT  5.055 0.185 5.125 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.390 -0.115 6.440 0.115 ;
        RECT  6.310 -0.115 6.390 0.465 ;
        RECT  6.050 -0.115 6.310 0.115 ;
        RECT  5.930 -0.115 6.050 0.275 ;
        RECT  5.665 -0.115 5.930 0.115 ;
        RECT  5.595 -0.115 5.665 0.465 ;
        RECT  5.330 -0.115 5.595 0.115 ;
        RECT  5.210 -0.115 5.330 0.275 ;
        RECT  4.945 -0.115 5.210 0.115 ;
        RECT  4.875 -0.115 4.945 0.305 ;
        RECT  4.565 -0.115 4.875 0.115 ;
        RECT  4.495 -0.115 4.565 0.320 ;
        RECT  3.625 -0.115 4.495 0.115 ;
        RECT  3.555 -0.115 3.625 0.460 ;
        RECT  3.265 -0.115 3.555 0.115 ;
        RECT  3.195 -0.115 3.265 0.400 ;
        RECT  2.340 -0.115 3.195 0.115 ;
        RECT  2.220 -0.115 2.340 0.135 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.390 1.145 6.440 1.375 ;
        RECT  6.310 0.675 6.390 1.375 ;
        RECT  6.025 1.145 6.310 1.375 ;
        RECT  5.955 0.975 6.025 1.375 ;
        RECT  5.690 1.145 5.955 1.375 ;
        RECT  5.570 1.010 5.690 1.375 ;
        RECT  5.330 1.145 5.570 1.375 ;
        RECT  5.210 1.010 5.330 1.375 ;
        RECT  4.970 1.145 5.210 1.375 ;
        RECT  4.850 1.010 4.970 1.375 ;
        RECT  4.570 1.145 4.850 1.375 ;
        RECT  4.500 0.950 4.570 1.375 ;
        RECT  3.640 1.145 4.500 1.375 ;
        RECT  3.540 0.860 3.640 1.375 ;
        RECT  3.265 1.145 3.540 1.375 ;
        RECT  3.195 0.860 3.265 1.375 ;
        RECT  2.360 1.145 3.195 1.375 ;
        RECT  2.240 1.115 2.360 1.375 ;
        RECT  1.800 1.145 2.240 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.845 0.355 5.915 0.465 ;
        RECT  5.845 0.765 5.915 0.905 ;
        RECT  5.775 0.185 5.845 0.465 ;
        RECT  5.775 0.765 5.845 1.065 ;
        RECT  5.425 0.700 5.510 0.800 ;
        RECT  5.425 0.185 5.485 0.485 ;
        RECT  5.055 0.185 5.075 0.485 ;
        RECT  5.030 0.700 5.075 0.800 ;
        RECT  5.670 0.545 5.810 0.615 ;
        RECT  5.600 0.545 5.670 0.940 ;
        RECT  4.920 0.870 5.600 0.940 ;
        RECT  4.850 0.435 4.920 0.940 ;
        RECT  4.745 0.435 4.850 0.505 ;
        RECT  4.745 0.870 4.850 0.940 ;
        RECT  4.675 0.200 4.745 0.505 ;
        RECT  4.675 0.870 4.745 1.010 ;
        RECT  4.410 0.585 4.710 0.655 ;
        RECT  4.380 0.435 4.675 0.505 ;
        RECT  4.340 0.585 4.410 1.055 ;
        RECT  4.300 0.585 4.340 0.655 ;
        RECT  3.805 0.985 4.340 1.055 ;
        RECT  4.230 0.270 4.300 0.655 ;
        RECT  4.180 0.780 4.270 0.910 ;
        RECT  4.185 0.270 4.230 0.340 ;
        RECT  4.115 0.195 4.185 0.340 ;
        RECT  4.130 0.780 4.180 0.850 ;
        RECT  4.060 0.485 4.130 0.850 ;
        RECT  3.800 0.195 4.115 0.265 ;
        RECT  4.010 0.485 4.060 0.555 ;
        RECT  3.940 0.335 4.010 0.405 ;
        RECT  3.940 0.710 3.985 0.890 ;
        RECT  3.915 0.335 3.940 0.890 ;
        RECT  3.870 0.335 3.915 0.780 ;
        RECT  3.485 0.710 3.870 0.780 ;
        RECT  3.735 0.850 3.805 1.055 ;
        RECT  3.730 0.195 3.800 0.350 ;
        RECT  3.445 0.335 3.485 0.780 ;
        RECT  3.415 0.335 3.445 0.980 ;
        RECT  3.350 0.335 3.415 0.405 ;
        RECT  3.375 0.710 3.415 0.980 ;
        RECT  3.155 0.710 3.375 0.780 ;
        RECT  3.265 0.510 3.335 0.640 ;
        RECT  2.885 0.510 3.265 0.580 ;
        RECT  3.085 0.660 3.155 0.780 ;
        RECT  2.875 0.510 2.885 0.980 ;
        RECT  2.805 0.280 2.875 0.980 ;
        RECT  2.680 0.205 2.735 0.935 ;
        RECT  2.665 0.205 2.680 1.045 ;
        RECT  1.945 0.205 2.665 0.275 ;
        RECT  2.610 0.865 2.665 1.045 ;
        RECT  2.080 0.975 2.610 1.045 ;
        RECT  2.525 0.345 2.595 0.765 ;
        RECT  2.435 0.345 2.525 0.465 ;
        RECT  2.455 0.695 2.525 0.850 ;
        RECT  2.345 0.545 2.440 0.620 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSND4BWP

MACRO SDFKSNQD0BWP
    CLASS CORE ;
    FOREIGN SDFKSNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.495 1.925 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.630 1.085 0.905 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0096 ;
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.195 4.305 1.045 ;
        RECT  4.215 0.195 4.235 0.415 ;
        RECT  4.215 0.905 4.235 1.045 ;
        RECT  3.985 0.345 4.215 0.415 ;
        RECT  3.915 0.345 3.985 0.610 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.635 0.550 0.755 ;
        RECT  0.445 0.635 0.525 0.905 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.495 2.235 0.640 ;
        RECT  2.135 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.120 -0.115 4.340 0.115 ;
        RECT  4.000 -0.115 4.120 0.255 ;
        RECT  3.315 -0.115 4.000 0.115 ;
        RECT  3.245 -0.115 3.315 0.420 ;
        RECT  2.360 -0.115 3.245 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.840 -0.115 2.240 0.115 ;
        RECT  1.720 -0.115 1.840 0.125 ;
        RECT  1.025 -0.115 1.720 0.115 ;
        RECT  0.955 -0.115 1.025 0.400 ;
        RECT  0.690 -0.115 0.955 0.115 ;
        RECT  0.570 -0.115 0.690 0.285 ;
        RECT  0.330 -0.115 0.570 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.110 1.145 4.340 1.375 ;
        RECT  4.040 0.915 4.110 1.375 ;
        RECT  3.320 1.145 4.040 1.375 ;
        RECT  3.200 0.870 3.320 1.375 ;
        RECT  2.360 1.145 3.200 1.375 ;
        RECT  2.240 1.130 2.360 1.375 ;
        RECT  1.840 1.145 2.240 1.375 ;
        RECT  1.720 1.135 1.840 1.375 ;
        RECT  1.020 1.145 1.720 1.375 ;
        RECT  0.900 1.135 1.020 1.375 ;
        RECT  0.330 1.145 0.900 1.375 ;
        RECT  0.210 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.510 4.165 0.750 ;
        RECT  3.970 0.680 4.095 0.750 ;
        RECT  3.900 0.680 3.970 1.060 ;
        RECT  3.810 0.680 3.900 0.750 ;
        RECT  3.580 0.990 3.900 1.060 ;
        RECT  3.670 0.830 3.820 0.900 ;
        RECT  3.740 0.195 3.810 0.750 ;
        RECT  3.610 0.195 3.740 0.265 ;
        RECT  3.600 0.430 3.670 0.900 ;
        RECT  3.495 0.220 3.530 0.800 ;
        RECT  3.460 0.220 3.495 1.070 ;
        RECT  3.445 0.220 3.460 0.340 ;
        RECT  3.425 0.730 3.460 1.070 ;
        RECT  3.195 0.730 3.425 0.800 ;
        RECT  3.315 0.510 3.385 0.640 ;
        RECT  2.915 0.510 3.315 0.580 ;
        RECT  3.125 0.675 3.195 0.800 ;
        RECT  2.905 0.300 2.915 0.580 ;
        RECT  2.835 0.300 2.905 0.960 ;
        RECT  1.405 0.195 2.760 0.265 ;
        RECT  2.655 0.840 2.725 1.060 ;
        RECT  1.300 0.990 2.655 1.060 ;
        RECT  2.550 0.355 2.615 0.765 ;
        RECT  2.545 0.355 2.550 0.850 ;
        RECT  2.450 0.355 2.545 0.425 ;
        RECT  2.475 0.695 2.545 0.850 ;
        RECT  2.375 0.520 2.430 0.640 ;
        RECT  2.305 0.355 2.375 0.915 ;
        RECT  2.070 0.355 2.305 0.425 ;
        RECT  2.070 0.845 2.305 0.915 ;
        RECT  1.675 0.335 1.990 0.405 ;
        RECT  1.675 0.845 1.990 0.915 ;
        RECT  1.605 0.335 1.675 0.915 ;
        RECT  1.415 0.475 1.485 0.760 ;
        RECT  0.845 0.475 1.415 0.545 ;
        RECT  1.335 0.195 1.405 0.400 ;
        RECT  1.225 0.665 1.330 0.735 ;
        RECT  1.155 0.665 1.225 1.065 ;
        RECT  0.690 0.995 1.155 1.065 ;
        RECT  0.775 0.210 0.845 0.920 ;
        RECT  0.620 0.355 0.690 1.065 ;
        RECT  0.485 0.355 0.620 0.425 ;
        RECT  0.595 0.920 0.620 1.065 ;
        RECT  0.415 0.215 0.485 0.425 ;
        RECT  0.345 0.520 0.375 0.640 ;
        RECT  0.275 0.355 0.345 0.915 ;
        RECT  0.125 0.355 0.275 0.425 ;
        RECT  0.125 0.845 0.275 0.915 ;
        RECT  0.055 0.210 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFKSNQD0BWP

MACRO SDFKSNQD1BWP
    CLASS CORE ;
    FOREIGN SDFKSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.195 4.585 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.385 -0.115 4.620 0.115 ;
        RECT  4.315 -0.115 4.385 0.305 ;
        RECT  4.025 -0.115 4.315 0.115 ;
        RECT  3.955 -0.115 4.025 0.285 ;
        RECT  3.265 -0.115 3.955 0.115 ;
        RECT  3.195 -0.115 3.265 0.420 ;
        RECT  2.340 -0.115 3.195 0.115 ;
        RECT  2.220 -0.115 2.340 0.135 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.385 1.145 4.620 1.375 ;
        RECT  4.315 0.905 4.385 1.375 ;
        RECT  4.030 1.145 4.315 1.375 ;
        RECT  3.960 0.955 4.030 1.375 ;
        RECT  3.290 1.145 3.960 1.375 ;
        RECT  3.170 0.870 3.290 1.375 ;
        RECT  2.360 1.145 3.170 1.375 ;
        RECT  2.240 1.115 2.360 1.375 ;
        RECT  1.800 1.145 2.240 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.345 0.395 4.415 0.820 ;
        RECT  4.205 0.395 4.345 0.465 ;
        RECT  4.205 0.750 4.345 0.820 ;
        RECT  3.890 0.545 4.250 0.615 ;
        RECT  4.135 0.185 4.205 0.465 ;
        RECT  4.135 0.750 4.205 1.075 ;
        RECT  3.860 0.395 4.135 0.465 ;
        RECT  3.820 0.545 3.890 1.060 ;
        RECT  3.770 0.545 3.820 0.615 ;
        RECT  3.530 0.990 3.820 1.060 ;
        RECT  3.700 0.195 3.770 0.615 ;
        RECT  3.610 0.800 3.750 0.920 ;
        RECT  3.550 0.195 3.700 0.265 ;
        RECT  3.540 0.440 3.610 0.920 ;
        RECT  3.445 0.220 3.470 0.800 ;
        RECT  3.400 0.220 3.445 1.050 ;
        RECT  3.385 0.220 3.400 0.340 ;
        RECT  3.375 0.730 3.400 1.050 ;
        RECT  3.155 0.730 3.375 0.800 ;
        RECT  3.260 0.510 3.330 0.640 ;
        RECT  2.890 0.510 3.260 0.580 ;
        RECT  3.085 0.680 3.155 0.800 ;
        RECT  2.875 0.510 2.890 0.960 ;
        RECT  2.805 0.300 2.875 0.960 ;
        RECT  2.680 0.205 2.735 0.935 ;
        RECT  2.665 0.205 2.680 1.045 ;
        RECT  1.945 0.205 2.665 0.275 ;
        RECT  2.610 0.865 2.665 1.045 ;
        RECT  2.080 0.975 2.610 1.045 ;
        RECT  2.525 0.345 2.595 0.765 ;
        RECT  2.435 0.345 2.525 0.465 ;
        RECT  2.455 0.695 2.525 0.890 ;
        RECT  2.345 0.545 2.440 0.620 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSNQD1BWP

MACRO SDFKSNQD2BWP
    CLASS CORE ;
    FOREIGN SDFKSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 0.355 4.585 0.805 ;
        RECT  4.515 0.185 4.525 1.035 ;
        RECT  4.455 0.185 4.515 0.465 ;
        RECT  4.455 0.735 4.515 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.300 ;
        RECT  4.345 -0.115 4.630 0.115 ;
        RECT  4.275 -0.115 4.345 0.305 ;
        RECT  3.965 -0.115 4.275 0.115 ;
        RECT  3.895 -0.115 3.965 0.290 ;
        RECT  3.225 -0.115 3.895 0.115 ;
        RECT  3.155 -0.115 3.225 0.420 ;
        RECT  2.320 -0.115 3.155 0.115 ;
        RECT  2.200 -0.115 2.320 0.135 ;
        RECT  1.790 -0.115 2.200 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.905 4.710 1.375 ;
        RECT  4.345 1.145 4.630 1.375 ;
        RECT  4.275 0.905 4.345 1.375 ;
        RECT  3.980 1.145 4.275 1.375 ;
        RECT  3.860 1.120 3.980 1.375 ;
        RECT  3.250 1.145 3.860 1.375 ;
        RECT  3.130 0.870 3.250 1.375 ;
        RECT  2.340 1.145 3.130 1.375 ;
        RECT  2.220 1.115 2.340 1.375 ;
        RECT  1.800 1.145 2.220 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.395 4.375 0.835 ;
        RECT  4.145 0.395 4.305 0.465 ;
        RECT  4.145 0.765 4.305 0.835 ;
        RECT  3.860 0.545 4.180 0.615 ;
        RECT  4.075 0.190 4.145 0.465 ;
        RECT  4.075 0.765 4.145 1.070 ;
        RECT  3.800 0.395 4.075 0.465 ;
        RECT  3.790 0.545 3.860 1.050 ;
        RECT  3.710 0.545 3.790 0.615 ;
        RECT  3.480 0.980 3.790 1.050 ;
        RECT  3.570 0.815 3.720 0.885 ;
        RECT  3.640 0.185 3.710 0.615 ;
        RECT  3.510 0.185 3.640 0.255 ;
        RECT  3.500 0.440 3.570 0.885 ;
        RECT  3.405 0.220 3.430 0.800 ;
        RECT  3.360 0.220 3.405 1.050 ;
        RECT  3.345 0.220 3.360 0.340 ;
        RECT  3.335 0.730 3.360 1.050 ;
        RECT  3.115 0.730 3.335 0.800 ;
        RECT  3.220 0.510 3.290 0.640 ;
        RECT  2.865 0.510 3.220 0.580 ;
        RECT  3.045 0.680 3.115 0.800 ;
        RECT  2.855 0.510 2.865 0.960 ;
        RECT  2.785 0.300 2.855 0.960 ;
        RECT  2.660 0.205 2.715 0.935 ;
        RECT  2.645 0.205 2.660 1.045 ;
        RECT  1.945 0.205 2.645 0.275 ;
        RECT  2.590 0.865 2.645 1.045 ;
        RECT  2.080 0.975 2.590 1.045 ;
        RECT  2.505 0.345 2.575 0.765 ;
        RECT  2.415 0.345 2.505 0.465 ;
        RECT  2.435 0.695 2.505 0.890 ;
        RECT  2.345 0.545 2.420 0.615 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSNQD2BWP

MACRO SDFKSNQD4BWP
    CLASS CORE ;
    FOREIGN SDFKSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.365 0.650 ;
        RECT  1.225 0.495 1.275 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0312 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.620 0.520 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.185 5.505 0.465 ;
        RECT  5.495 0.765 5.505 1.065 ;
        RECT  5.435 0.185 5.495 1.065 ;
        RECT  5.285 0.355 5.435 0.905 ;
        RECT  5.150 0.355 5.285 0.465 ;
        RECT  5.150 0.765 5.285 0.905 ;
        RECT  5.080 0.185 5.150 0.465 ;
        RECT  5.080 0.765 5.150 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.735 0.640 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.465 ;
        RECT  5.350 -0.115 5.610 0.115 ;
        RECT  5.230 -0.115 5.350 0.275 ;
        RECT  4.965 -0.115 5.230 0.115 ;
        RECT  4.895 -0.115 4.965 0.305 ;
        RECT  4.585 -0.115 4.895 0.115 ;
        RECT  4.515 -0.115 4.585 0.320 ;
        RECT  3.645 -0.115 4.515 0.115 ;
        RECT  3.575 -0.115 3.645 0.460 ;
        RECT  3.275 -0.115 3.575 0.115 ;
        RECT  3.205 -0.115 3.275 0.400 ;
        RECT  2.340 -0.115 3.205 0.115 ;
        RECT  2.220 -0.115 2.340 0.135 ;
        RECT  1.790 -0.115 2.220 0.115 ;
        RECT  1.670 -0.115 1.790 0.265 ;
        RECT  1.405 -0.115 1.670 0.115 ;
        RECT  1.315 -0.115 1.405 0.425 ;
        RECT  0.690 -0.115 1.315 0.115 ;
        RECT  0.550 -0.115 0.690 0.150 ;
        RECT  0.330 -0.115 0.550 0.115 ;
        RECT  0.210 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.675 5.690 1.375 ;
        RECT  5.325 1.145 5.610 1.375 ;
        RECT  5.255 0.975 5.325 1.375 ;
        RECT  4.965 1.145 5.255 1.375 ;
        RECT  4.895 0.905 4.965 1.375 ;
        RECT  4.575 1.145 4.895 1.375 ;
        RECT  4.505 0.940 4.575 1.375 ;
        RECT  3.660 1.145 4.505 1.375 ;
        RECT  3.560 0.860 3.660 1.375 ;
        RECT  3.275 1.145 3.560 1.375 ;
        RECT  3.205 0.860 3.275 1.375 ;
        RECT  2.360 1.145 3.205 1.375 ;
        RECT  2.240 1.115 2.360 1.375 ;
        RECT  1.800 1.145 2.240 1.375 ;
        RECT  1.680 1.110 1.800 1.375 ;
        RECT  1.460 1.145 1.680 1.375 ;
        RECT  1.340 1.010 1.460 1.375 ;
        RECT  0.330 1.145 1.340 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.150 0.355 5.215 0.465 ;
        RECT  5.150 0.765 5.215 0.905 ;
        RECT  5.080 0.185 5.150 0.465 ;
        RECT  5.080 0.765 5.150 1.065 ;
        RECT  4.940 0.395 5.010 0.835 ;
        RECT  4.765 0.395 4.940 0.465 ;
        RECT  4.765 0.765 4.940 0.835 ;
        RECT  4.430 0.545 4.870 0.615 ;
        RECT  4.695 0.200 4.765 0.465 ;
        RECT  4.695 0.765 4.765 1.070 ;
        RECT  4.400 0.395 4.695 0.465 ;
        RECT  4.360 0.545 4.430 1.055 ;
        RECT  4.320 0.545 4.360 0.615 ;
        RECT  3.825 0.985 4.360 1.055 ;
        RECT  4.250 0.270 4.320 0.615 ;
        RECT  4.200 0.780 4.290 0.910 ;
        RECT  4.205 0.270 4.250 0.340 ;
        RECT  4.135 0.195 4.205 0.340 ;
        RECT  4.150 0.780 4.200 0.850 ;
        RECT  4.080 0.485 4.150 0.850 ;
        RECT  3.820 0.195 4.135 0.265 ;
        RECT  4.030 0.485 4.080 0.555 ;
        RECT  3.960 0.335 4.030 0.405 ;
        RECT  3.960 0.710 4.005 0.890 ;
        RECT  3.935 0.335 3.960 0.890 ;
        RECT  3.890 0.335 3.935 0.780 ;
        RECT  3.505 0.710 3.890 0.780 ;
        RECT  3.755 0.850 3.825 1.055 ;
        RECT  3.750 0.195 3.820 0.350 ;
        RECT  3.465 0.335 3.505 0.780 ;
        RECT  3.435 0.335 3.465 0.980 ;
        RECT  3.370 0.335 3.435 0.405 ;
        RECT  3.395 0.710 3.435 0.980 ;
        RECT  3.155 0.710 3.395 0.780 ;
        RECT  3.285 0.510 3.355 0.640 ;
        RECT  2.885 0.510 3.285 0.580 ;
        RECT  3.085 0.660 3.155 0.780 ;
        RECT  2.875 0.510 2.885 0.980 ;
        RECT  2.805 0.280 2.875 0.980 ;
        RECT  2.680 0.205 2.735 0.935 ;
        RECT  2.665 0.205 2.680 1.045 ;
        RECT  1.945 0.205 2.665 0.275 ;
        RECT  2.610 0.865 2.665 1.045 ;
        RECT  2.080 0.975 2.610 1.045 ;
        RECT  2.525 0.345 2.595 0.765 ;
        RECT  2.435 0.345 2.525 0.465 ;
        RECT  2.455 0.695 2.525 0.850 ;
        RECT  2.345 0.545 2.440 0.620 ;
        RECT  2.275 0.355 2.345 0.905 ;
        RECT  2.030 0.355 2.275 0.425 ;
        RECT  2.050 0.835 2.275 0.905 ;
        RECT  2.010 0.975 2.080 1.060 ;
        RECT  1.870 0.990 2.010 1.060 ;
        RECT  1.875 0.205 1.945 0.410 ;
        RECT  1.855 0.510 1.930 0.915 ;
        RECT  1.765 0.845 1.855 0.915 ;
        RECT  1.705 0.845 1.765 0.930 ;
        RECT  1.025 0.860 1.705 0.930 ;
        RECT  1.545 0.720 1.630 0.790 ;
        RECT  1.545 0.190 1.585 0.310 ;
        RECT  1.475 0.190 1.545 0.790 ;
        RECT  1.175 0.720 1.475 0.790 ;
        RECT  1.105 0.640 1.175 0.790 ;
        RECT  0.955 0.210 1.025 1.060 ;
        RECT  0.845 0.280 0.880 0.840 ;
        RECT  0.810 0.280 0.845 1.060 ;
        RECT  0.485 0.280 0.810 0.350 ;
        RECT  0.775 0.770 0.810 1.060 ;
        RECT  0.485 0.935 0.700 1.005 ;
        RECT  0.415 0.230 0.485 0.350 ;
        RECT  0.415 0.935 0.485 1.070 ;
        RECT  0.330 0.545 0.400 0.615 ;
        RECT  0.260 0.345 0.330 0.915 ;
        RECT  0.125 0.345 0.260 0.415 ;
        RECT  0.125 0.845 0.260 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END SDFKSNQD4BWP

MACRO SDFNCND0BWP
    CLASS CORE ;
    FOREIGN SDFNCND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.215 4.585 0.905 ;
        RECT  4.495 0.215 4.515 0.335 ;
        RECT  4.500 0.775 4.515 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 0.715 4.220 0.785 ;
        RECT  4.090 0.215 4.185 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0330 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.355 3.745 0.640 ;
        RECT  3.605 0.520 3.665 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 -0.115 4.620 0.115 ;
        RECT  4.300 -0.115 4.380 0.335 ;
        RECT  3.555 -0.115 4.300 0.115 ;
        RECT  3.485 -0.115 3.555 0.440 ;
        RECT  2.550 -0.115 3.485 0.115 ;
        RECT  2.480 -0.115 2.550 0.320 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 1.145 4.620 1.375 ;
        RECT  4.260 1.130 4.380 1.375 ;
        RECT  3.620 1.145 4.260 1.375 ;
        RECT  3.500 1.135 3.620 1.375 ;
        RECT  2.660 1.145 3.500 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.650 ;
        RECT  4.355 0.520 4.425 0.925 ;
        RECT  3.360 0.855 4.355 0.925 ;
        RECT  3.945 0.520 4.020 0.640 ;
        RECT  3.875 0.190 3.945 0.785 ;
        RECT  3.500 0.715 3.875 0.785 ;
        RECT  3.740 0.995 3.860 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.785 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.255 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.685 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.755 ;
        RECT  2.100 0.685 2.760 0.755 ;
        RECT  2.620 0.205 2.690 0.470 ;
        RECT  2.505 0.540 2.680 0.610 ;
        RECT  2.300 0.400 2.620 0.470 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.455 0.540 2.505 0.615 ;
        RECT  1.945 0.545 2.455 0.615 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.125 0.840 2.240 0.910 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  2.055 0.840 2.125 0.960 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.960 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.740 0.195 1.735 0.265 ;
        RECT  1.660 0.545 1.720 0.615 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.920 0.490 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFNCND0BWP

MACRO SDFNCND1BWP
    CLASS CORE ;
    FOREIGN SDFNCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.585 1.045 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.735 4.515 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 0.715 4.220 0.785 ;
        RECT  4.090 0.185 4.185 0.785 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0330 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.355 3.745 0.640 ;
        RECT  3.605 0.520 3.665 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 -0.115 4.620 0.115 ;
        RECT  4.300 -0.115 4.380 0.445 ;
        RECT  3.535 -0.115 4.300 0.115 ;
        RECT  3.465 -0.115 3.535 0.440 ;
        RECT  2.550 -0.115 3.465 0.115 ;
        RECT  2.480 -0.115 2.550 0.320 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 1.005 4.400 1.375 ;
        RECT  3.620 1.145 4.280 1.375 ;
        RECT  3.500 1.135 3.620 1.375 ;
        RECT  2.660 1.145 3.500 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.410 0.520 4.440 0.640 ;
        RECT  4.340 0.520 4.410 0.925 ;
        RECT  3.360 0.855 4.340 0.925 ;
        RECT  3.945 0.520 4.020 0.640 ;
        RECT  3.875 0.190 3.945 0.785 ;
        RECT  3.500 0.715 3.875 0.785 ;
        RECT  3.740 0.995 3.860 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.785 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.255 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.685 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.755 ;
        RECT  2.100 0.685 2.760 0.755 ;
        RECT  2.620 0.205 2.690 0.470 ;
        RECT  2.505 0.540 2.680 0.610 ;
        RECT  2.300 0.400 2.620 0.470 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.455 0.540 2.505 0.615 ;
        RECT  1.945 0.545 2.455 0.615 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.125 0.840 2.240 0.910 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  2.055 0.840 2.125 0.960 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.960 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.660 0.545 1.720 0.615 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCND1BWP

MACRO SDFNCND2BWP
    CLASS CORE ;
    FOREIGN SDFNCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.945 0.355 5.005 0.805 ;
        RECT  4.935 0.185 4.945 1.035 ;
        RECT  4.875 0.185 4.935 0.465 ;
        RECT  4.875 0.735 4.935 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.590 0.780 ;
        RECT  4.495 0.185 4.515 0.485 ;
        RECT  4.470 0.710 4.515 0.780 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.580 0.535 3.675 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.130 0.300 ;
        RECT  4.755 -0.115 5.050 0.115 ;
        RECT  4.685 -0.115 4.755 0.465 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.275 ;
        RECT  3.555 -0.115 4.280 0.115 ;
        RECT  3.485 -0.115 3.555 0.400 ;
        RECT  2.550 -0.115 3.485 0.115 ;
        RECT  2.480 -0.115 2.550 0.320 ;
        RECT  1.440 -0.115 2.480 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.145 5.180 1.375 ;
        RECT  5.050 0.895 5.130 1.375 ;
        RECT  4.780 1.145 5.050 1.375 ;
        RECT  4.660 0.995 4.780 1.375 ;
        RECT  4.410 1.145 4.660 1.375 ;
        RECT  4.290 0.995 4.410 1.375 ;
        RECT  2.660 1.145 4.290 1.375 ;
        RECT  2.540 1.060 2.660 1.375 ;
        RECT  1.400 1.145 2.540 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.805 0.545 4.860 0.615 ;
        RECT  4.735 0.545 4.805 0.925 ;
        RECT  3.360 0.855 4.735 0.925 ;
        RECT  4.375 0.520 4.430 0.640 ;
        RECT  4.305 0.350 4.375 0.780 ;
        RECT  3.840 0.350 4.305 0.420 ;
        RECT  3.500 0.710 4.305 0.780 ;
        RECT  3.740 0.995 3.870 1.075 ;
        RECT  3.160 0.995 3.740 1.065 ;
        RECT  3.430 0.520 3.500 0.780 ;
        RECT  3.290 0.320 3.360 0.925 ;
        RECT  3.235 0.320 3.290 0.440 ;
        RECT  3.165 0.670 3.215 0.895 ;
        RECT  3.145 0.205 3.165 0.895 ;
        RECT  3.090 0.975 3.160 1.065 ;
        RECT  3.095 0.205 3.145 0.740 ;
        RECT  2.690 0.205 3.095 0.275 ;
        RECT  3.025 0.975 3.090 1.045 ;
        RECT  2.955 0.360 3.025 1.045 ;
        RECT  2.830 0.685 2.885 1.040 ;
        RECT  2.815 0.360 2.830 1.040 ;
        RECT  2.760 0.360 2.815 0.755 ;
        RECT  2.100 0.685 2.760 0.755 ;
        RECT  2.620 0.205 2.690 0.470 ;
        RECT  2.505 0.540 2.670 0.610 ;
        RECT  2.300 0.400 2.620 0.470 ;
        RECT  2.300 0.830 2.510 0.900 ;
        RECT  2.455 0.540 2.505 0.615 ;
        RECT  1.945 0.545 2.455 0.615 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.240 0.830 2.300 0.910 ;
        RECT  2.125 0.840 2.240 0.910 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  2.055 0.840 2.125 0.960 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.960 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.660 0.545 1.720 0.615 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCND2BWP

MACRO SDFNCND4BWP
    CLASS CORE ;
    FOREIGN SDFNCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.185 5.925 0.465 ;
        RECT  5.915 0.775 5.925 1.065 ;
        RECT  5.855 0.185 5.915 1.065 ;
        RECT  5.705 0.355 5.855 0.905 ;
        RECT  5.565 0.355 5.705 0.465 ;
        RECT  5.565 0.775 5.705 0.905 ;
        RECT  5.495 0.185 5.565 0.465 ;
        RECT  5.495 0.775 5.565 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.705 5.230 0.795 ;
        RECT  5.135 0.185 5.205 0.485 ;
        RECT  5.075 0.355 5.135 0.485 ;
        RECT  4.865 0.355 5.075 0.795 ;
        RECT  4.845 0.355 4.865 0.485 ;
        RECT  4.750 0.705 4.865 0.795 ;
        RECT  4.775 0.185 4.845 0.485 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0532 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.535 0.495 3.675 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 -0.115 6.160 0.115 ;
        RECT  6.035 -0.115 6.105 0.465 ;
        RECT  5.770 -0.115 6.035 0.115 ;
        RECT  5.650 -0.115 5.770 0.275 ;
        RECT  5.385 -0.115 5.650 0.115 ;
        RECT  5.315 -0.115 5.385 0.465 ;
        RECT  5.050 -0.115 5.315 0.115 ;
        RECT  4.930 -0.115 5.050 0.275 ;
        RECT  4.665 -0.115 4.930 0.115 ;
        RECT  4.595 -0.115 4.665 0.310 ;
        RECT  4.340 -0.115 4.595 0.115 ;
        RECT  4.220 -0.115 4.340 0.145 ;
        RECT  3.325 -0.115 4.220 0.115 ;
        RECT  3.255 -0.115 3.325 0.250 ;
        RECT  2.570 -0.115 3.255 0.115 ;
        RECT  2.500 -0.115 2.570 0.320 ;
        RECT  1.480 -0.115 2.500 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  1.130 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.130 0.135 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 1.145 6.160 1.375 ;
        RECT  6.035 0.675 6.105 1.375 ;
        RECT  5.745 1.145 6.035 1.375 ;
        RECT  5.675 0.975 5.745 1.375 ;
        RECT  5.410 1.145 5.675 1.375 ;
        RECT  5.290 1.005 5.410 1.375 ;
        RECT  5.050 1.145 5.290 1.375 ;
        RECT  4.930 1.005 5.050 1.375 ;
        RECT  4.690 1.145 4.930 1.375 ;
        RECT  4.570 1.005 4.690 1.375 ;
        RECT  4.330 1.145 4.570 1.375 ;
        RECT  4.210 1.005 4.330 1.375 ;
        RECT  2.680 1.145 4.210 1.375 ;
        RECT  2.560 1.055 2.680 1.375 ;
        RECT  1.440 1.145 2.560 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.355 5.635 0.465 ;
        RECT  5.565 0.775 5.635 0.905 ;
        RECT  5.495 0.185 5.565 0.465 ;
        RECT  5.495 0.775 5.565 1.065 ;
        RECT  5.145 0.705 5.230 0.795 ;
        RECT  5.145 0.185 5.205 0.485 ;
        RECT  4.775 0.185 4.795 0.485 ;
        RECT  4.750 0.705 4.795 0.795 ;
        RECT  5.400 0.545 5.540 0.615 ;
        RECT  5.330 0.545 5.400 0.935 ;
        RECT  4.680 0.865 5.330 0.935 ;
        RECT  4.610 0.395 4.680 0.935 ;
        RECT  4.485 0.395 4.610 0.465 ;
        RECT  4.485 0.865 4.610 0.935 ;
        RECT  4.415 0.185 4.485 0.465 ;
        RECT  4.415 0.735 4.485 1.035 ;
        RECT  4.150 0.545 4.460 0.615 ;
        RECT  4.150 0.260 4.415 0.330 ;
        RECT  3.270 0.855 4.415 0.925 ;
        RECT  4.080 0.205 4.150 0.330 ;
        RECT  4.080 0.400 4.150 0.780 ;
        RECT  3.595 0.205 4.080 0.275 ;
        RECT  3.820 0.400 4.080 0.470 ;
        RECT  3.455 0.710 4.080 0.780 ;
        RECT  3.720 0.995 3.850 1.075 ;
        RECT  3.180 0.995 3.720 1.065 ;
        RECT  3.525 0.205 3.595 0.400 ;
        RECT  3.325 0.330 3.525 0.400 ;
        RECT  3.385 0.520 3.455 0.780 ;
        RECT  3.255 0.330 3.325 0.460 ;
        RECT  3.185 0.685 3.290 0.755 ;
        RECT  3.115 0.205 3.185 0.755 ;
        RECT  3.110 0.965 3.180 1.065 ;
        RECT  2.710 0.205 3.115 0.275 ;
        RECT  3.045 0.965 3.110 1.035 ;
        RECT  2.975 0.360 3.045 1.035 ;
        RECT  2.850 0.685 2.905 1.040 ;
        RECT  2.835 0.360 2.850 1.040 ;
        RECT  2.780 0.360 2.835 0.755 ;
        RECT  2.120 0.685 2.780 0.755 ;
        RECT  2.640 0.205 2.710 0.470 ;
        RECT  2.525 0.540 2.690 0.610 ;
        RECT  2.320 0.400 2.640 0.470 ;
        RECT  2.320 0.830 2.530 0.900 ;
        RECT  2.475 0.540 2.525 0.615 ;
        RECT  1.965 0.545 2.475 0.615 ;
        RECT  2.225 0.375 2.320 0.470 ;
        RECT  2.260 0.830 2.320 0.910 ;
        RECT  2.145 0.840 2.260 0.910 ;
        RECT  2.040 0.375 2.225 0.445 ;
        RECT  2.075 0.840 2.145 0.960 ;
        RECT  1.965 0.225 2.060 0.295 ;
        RECT  1.895 0.225 1.965 0.960 ;
        RECT  1.755 0.205 1.825 0.430 ;
        RECT  0.685 0.985 1.810 1.055 ;
        RECT  0.610 0.205 1.755 0.275 ;
        RECT  1.680 0.545 1.740 0.615 ;
        RECT  1.610 0.350 1.680 0.905 ;
        RECT  1.540 0.350 1.610 0.420 ;
        RECT  1.510 0.835 1.610 0.905 ;
        RECT  1.410 0.520 1.530 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCND4BWP

MACRO SDFNCSND0BWP
    CLASS CORE ;
    FOREIGN SDFNCSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.760 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.195 5.005 1.045 ;
        RECT  4.915 0.195 4.935 0.315 ;
        RECT  4.915 0.910 4.935 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.695 0.775 4.730 1.045 ;
        RECT  4.625 0.350 4.695 1.045 ;
        RECT  4.535 0.350 4.625 0.470 ;
        RECT  4.540 0.920 4.625 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.495 4.165 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.140 ;
        RECT  4.070 -0.115 4.700 0.115 ;
        RECT  3.950 -0.115 4.070 0.275 ;
        RECT  2.560 -0.115 3.950 0.115 ;
        RECT  2.490 -0.115 2.560 0.320 ;
        RECT  1.440 -0.115 2.490 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 1.120 4.820 1.375 ;
        RECT  4.450 1.145 4.700 1.375 ;
        RECT  4.330 1.120 4.450 1.375 ;
        RECT  4.040 1.145 4.330 1.375 ;
        RECT  3.920 1.130 4.040 1.375 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 0.990 3.690 1.375 ;
        RECT  2.900 1.145 3.570 1.375 ;
        RECT  2.780 1.120 2.900 1.375 ;
        RECT  2.380 1.145 2.780 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.835 0.520 4.860 0.640 ;
        RECT  4.765 0.210 4.835 0.640 ;
        RECT  4.220 0.210 4.765 0.280 ;
        RECT  4.460 0.545 4.540 0.615 ;
        RECT  4.390 0.355 4.460 1.050 ;
        RECT  4.320 0.355 4.390 0.425 ;
        RECT  3.820 0.975 4.390 1.050 ;
        RECT  4.245 0.520 4.315 0.905 ;
        RECT  3.305 0.835 4.245 0.905 ;
        RECT  4.150 0.210 4.220 0.425 ;
        RECT  3.450 0.355 4.150 0.425 ;
        RECT  3.450 0.695 3.870 0.765 ;
        RECT  2.700 0.205 3.470 0.275 ;
        RECT  3.380 0.355 3.450 0.765 ;
        RECT  3.250 0.375 3.380 0.445 ;
        RECT  3.235 0.630 3.305 0.905 ;
        RECT  3.145 0.630 3.235 0.700 ;
        RECT  3.095 0.980 3.230 1.050 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  3.025 0.970 3.095 1.050 ;
        RECT  2.965 0.830 3.090 0.900 ;
        RECT  2.700 0.970 3.025 1.040 ;
        RECT  2.895 0.350 2.965 0.900 ;
        RECT  2.685 0.830 2.895 0.900 ;
        RECT  1.945 0.545 2.740 0.615 ;
        RECT  2.630 0.205 2.700 0.470 ;
        RECT  2.630 0.970 2.700 1.065 ;
        RECT  2.615 0.685 2.685 0.900 ;
        RECT  2.300 0.400 2.630 0.470 ;
        RECT  2.080 0.995 2.630 1.065 ;
        RECT  2.160 0.685 2.615 0.755 ;
        RECT  2.050 0.840 2.530 0.910 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  1.960 0.995 2.080 1.075 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.915 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.740 0.195 1.735 0.265 ;
        RECT  1.660 0.535 1.720 0.605 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.920 0.490 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFNCSND0BWP

MACRO SDFNCSND1BWP
    CLASS CORE ;
    FOREIGN SDFNCSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.760 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.045 ;
        RECT  4.915 0.185 4.935 0.465 ;
        RECT  4.915 0.750 4.935 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.695 0.775 4.730 1.045 ;
        RECT  4.625 0.350 4.695 1.045 ;
        RECT  4.535 0.350 4.625 0.470 ;
        RECT  4.540 0.775 4.625 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 0.495 4.165 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.140 ;
        RECT  4.070 -0.115 4.700 0.115 ;
        RECT  3.950 -0.115 4.070 0.275 ;
        RECT  2.560 -0.115 3.950 0.115 ;
        RECT  2.490 -0.115 2.560 0.320 ;
        RECT  1.440 -0.115 2.490 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 1.120 4.820 1.375 ;
        RECT  4.450 1.145 4.700 1.375 ;
        RECT  4.330 1.120 4.450 1.375 ;
        RECT  4.040 1.145 4.330 1.375 ;
        RECT  3.920 1.130 4.040 1.375 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 0.990 3.690 1.375 ;
        RECT  2.900 1.145 3.570 1.375 ;
        RECT  2.780 1.120 2.900 1.375 ;
        RECT  2.380 1.145 2.780 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.835 0.520 4.860 0.640 ;
        RECT  4.765 0.210 4.835 0.640 ;
        RECT  4.220 0.210 4.765 0.280 ;
        RECT  4.460 0.545 4.540 0.615 ;
        RECT  4.390 0.355 4.460 1.050 ;
        RECT  4.320 0.355 4.390 0.425 ;
        RECT  3.820 0.975 4.390 1.050 ;
        RECT  4.245 0.520 4.315 0.905 ;
        RECT  3.305 0.835 4.245 0.905 ;
        RECT  4.150 0.210 4.220 0.425 ;
        RECT  3.450 0.355 4.150 0.425 ;
        RECT  3.450 0.695 3.870 0.765 ;
        RECT  2.700 0.205 3.470 0.275 ;
        RECT  3.380 0.355 3.450 0.765 ;
        RECT  3.250 0.375 3.380 0.445 ;
        RECT  3.235 0.630 3.305 0.905 ;
        RECT  3.145 0.630 3.235 0.700 ;
        RECT  3.095 0.980 3.230 1.050 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  3.025 0.970 3.095 1.050 ;
        RECT  2.965 0.830 3.090 0.900 ;
        RECT  2.700 0.970 3.025 1.040 ;
        RECT  2.895 0.350 2.965 0.900 ;
        RECT  2.685 0.830 2.895 0.900 ;
        RECT  1.945 0.545 2.740 0.615 ;
        RECT  2.630 0.205 2.700 0.470 ;
        RECT  2.630 0.970 2.700 1.065 ;
        RECT  2.615 0.685 2.685 0.900 ;
        RECT  2.300 0.400 2.630 0.470 ;
        RECT  2.080 0.995 2.630 1.065 ;
        RECT  2.160 0.685 2.615 0.755 ;
        RECT  2.050 0.840 2.530 0.910 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  1.960 0.995 2.080 1.075 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.915 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.660 0.535 1.720 0.605 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCSND1BWP

MACRO SDFNCSND2BWP
    CLASS CORE ;
    FOREIGN SDFNCSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.745 0.625 ;
        RECT  3.600 0.540 3.675 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.355 5.145 0.810 ;
        RECT  5.075 0.185 5.085 1.040 ;
        RECT  5.015 0.185 5.075 0.465 ;
        RECT  5.015 0.740 5.075 1.040 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.690 0.350 4.760 1.045 ;
        RECT  4.620 0.350 4.690 0.450 ;
        RECT  4.655 0.735 4.690 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.495 4.165 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.300 ;
        RECT  4.920 -0.115 5.190 0.115 ;
        RECT  4.800 -0.115 4.920 0.140 ;
        RECT  4.540 -0.115 4.800 0.115 ;
        RECT  4.420 -0.115 4.540 0.140 ;
        RECT  4.010 -0.115 4.420 0.115 ;
        RECT  3.890 -0.115 4.010 0.275 ;
        RECT  2.555 -0.115 3.890 0.115 ;
        RECT  2.485 -0.115 2.555 0.320 ;
        RECT  1.440 -0.115 2.485 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.265 1.145 5.320 1.375 ;
        RECT  5.195 0.905 5.265 1.375 ;
        RECT  4.905 1.145 5.195 1.375 ;
        RECT  4.835 0.745 4.905 1.375 ;
        RECT  4.545 1.145 4.835 1.375 ;
        RECT  4.475 0.980 4.545 1.375 ;
        RECT  4.390 1.145 4.475 1.375 ;
        RECT  4.270 0.980 4.390 1.375 ;
        RECT  4.000 1.145 4.270 1.375 ;
        RECT  3.880 1.130 4.000 1.375 ;
        RECT  3.640 1.145 3.880 1.375 ;
        RECT  3.520 0.990 3.640 1.375 ;
        RECT  2.360 1.145 3.520 1.375 ;
        RECT  2.240 1.135 2.360 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.910 0.545 5.000 0.615 ;
        RECT  4.840 0.210 4.910 0.615 ;
        RECT  4.170 0.210 4.840 0.280 ;
        RECT  4.525 0.520 4.620 0.640 ;
        RECT  4.455 0.350 4.525 0.905 ;
        RECT  4.250 0.350 4.455 0.420 ;
        RECT  4.185 0.835 4.455 0.905 ;
        RECT  4.305 0.520 4.375 0.765 ;
        RECT  4.045 0.695 4.305 0.765 ;
        RECT  4.115 0.835 4.185 1.045 ;
        RECT  4.100 0.210 4.170 0.425 ;
        RECT  3.780 0.975 4.115 1.045 ;
        RECT  3.885 0.355 4.100 0.425 ;
        RECT  3.975 0.695 4.045 0.905 ;
        RECT  3.265 0.835 3.975 0.905 ;
        RECT  3.815 0.355 3.885 0.765 ;
        RECT  3.410 0.695 3.815 0.765 ;
        RECT  3.530 0.305 3.605 0.445 ;
        RECT  3.410 0.375 3.530 0.445 ;
        RECT  2.700 0.205 3.440 0.275 ;
        RECT  3.340 0.375 3.410 0.765 ;
        RECT  3.210 0.375 3.340 0.445 ;
        RECT  3.195 0.630 3.265 0.905 ;
        RECT  3.110 0.985 3.230 1.065 ;
        RECT  3.125 0.630 3.195 0.700 ;
        RECT  3.055 0.350 3.125 0.700 ;
        RECT  2.945 0.825 3.110 0.895 ;
        RECT  2.080 0.995 3.110 1.065 ;
        RECT  2.875 0.350 2.945 0.895 ;
        RECT  2.665 0.825 2.875 0.895 ;
        RECT  2.630 0.205 2.700 0.470 ;
        RECT  1.945 0.545 2.700 0.615 ;
        RECT  2.595 0.685 2.665 0.925 ;
        RECT  2.300 0.400 2.630 0.470 ;
        RECT  2.140 0.685 2.595 0.755 ;
        RECT  2.030 0.840 2.510 0.910 ;
        RECT  2.205 0.375 2.300 0.470 ;
        RECT  2.020 0.375 2.205 0.445 ;
        RECT  1.960 0.995 2.080 1.075 ;
        RECT  1.945 0.225 2.040 0.295 ;
        RECT  1.875 0.225 1.945 0.915 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.660 0.535 1.720 0.605 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.940 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.820 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCSND2BWP

MACRO SDFNCSND4BWP
    CLASS CORE ;
    FOREIGN SDFNCSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0324 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.745 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.185 6.065 0.465 ;
        RECT  6.055 0.775 6.065 1.055 ;
        RECT  5.995 0.185 6.055 1.055 ;
        RECT  5.845 0.355 5.995 0.905 ;
        RECT  5.705 0.355 5.845 0.465 ;
        RECT  5.705 0.775 5.845 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.775 5.705 1.055 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.350 5.350 0.470 ;
        RECT  5.255 0.775 5.325 1.055 ;
        RECT  5.215 0.775 5.255 0.905 ;
        RECT  5.005 0.350 5.215 0.905 ;
        RECT  4.880 0.350 5.005 0.470 ;
        RECT  4.985 0.775 5.005 0.905 ;
        RECT  4.895 0.775 4.985 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.0592 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.585 0.495 4.670 0.640 ;
        RECT  4.515 0.495 4.585 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 -0.115 6.300 0.115 ;
        RECT  6.175 -0.115 6.245 0.465 ;
        RECT  5.885 -0.115 6.175 0.115 ;
        RECT  5.815 -0.115 5.885 0.280 ;
        RECT  5.540 -0.115 5.815 0.115 ;
        RECT  5.420 -0.115 5.540 0.140 ;
        RECT  5.160 -0.115 5.420 0.115 ;
        RECT  5.040 -0.115 5.160 0.140 ;
        RECT  4.780 -0.115 5.040 0.115 ;
        RECT  4.660 -0.115 4.780 0.140 ;
        RECT  4.015 -0.115 4.660 0.115 ;
        RECT  3.945 -0.115 4.015 0.270 ;
        RECT  2.575 -0.115 3.945 0.115 ;
        RECT  2.505 -0.115 2.575 0.320 ;
        RECT  1.480 -0.115 2.505 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.245 1.145 6.300 1.375 ;
        RECT  6.175 0.675 6.245 1.375 ;
        RECT  5.885 1.145 6.175 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  5.515 1.145 5.815 1.375 ;
        RECT  5.445 0.745 5.515 1.375 ;
        RECT  5.150 1.145 5.445 1.375 ;
        RECT  5.070 0.975 5.150 1.375 ;
        RECT  4.810 1.145 5.070 1.375 ;
        RECT  4.690 1.005 4.810 1.375 ;
        RECT  4.450 1.145 4.690 1.375 ;
        RECT  4.330 1.005 4.450 1.375 ;
        RECT  4.070 1.145 4.330 1.375 ;
        RECT  3.950 1.005 4.070 1.375 ;
        RECT  3.660 1.145 3.950 1.375 ;
        RECT  3.540 1.010 3.660 1.375 ;
        RECT  2.920 1.145 3.540 1.375 ;
        RECT  2.800 1.135 2.920 1.375 ;
        RECT  2.380 1.145 2.800 1.375 ;
        RECT  2.260 1.135 2.380 1.375 ;
        RECT  1.440 1.145 2.260 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.355 5.775 0.465 ;
        RECT  5.705 0.775 5.775 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.775 5.705 1.055 ;
        RECT  5.285 0.350 5.350 0.470 ;
        RECT  5.285 0.775 5.325 1.055 ;
        RECT  4.880 0.350 4.935 0.470 ;
        RECT  4.895 0.775 4.935 1.065 ;
        RECT  5.530 0.545 5.670 0.615 ;
        RECT  5.460 0.210 5.530 0.615 ;
        RECT  4.165 0.210 5.460 0.280 ;
        RECT  4.810 0.545 4.910 0.615 ;
        RECT  4.740 0.350 4.810 0.915 ;
        RECT  4.305 0.350 4.740 0.420 ;
        RECT  4.605 0.845 4.740 0.915 ;
        RECT  4.535 0.845 4.605 1.075 ;
        RECT  4.150 0.845 4.535 0.915 ;
        RECT  4.375 0.520 4.445 0.755 ;
        RECT  4.060 0.685 4.375 0.755 ;
        RECT  4.235 0.350 4.305 0.615 ;
        RECT  3.840 0.545 4.235 0.615 ;
        RECT  4.095 0.210 4.165 0.425 ;
        RECT  3.430 0.355 4.095 0.425 ;
        RECT  3.990 0.685 4.060 0.915 ;
        RECT  3.285 0.845 3.990 0.915 ;
        RECT  3.430 0.700 3.860 0.770 ;
        RECT  2.720 0.205 3.460 0.275 ;
        RECT  3.360 0.355 3.430 0.770 ;
        RECT  3.230 0.375 3.360 0.445 ;
        RECT  3.215 0.630 3.285 0.915 ;
        RECT  3.130 0.985 3.250 1.065 ;
        RECT  3.145 0.630 3.215 0.700 ;
        RECT  3.075 0.350 3.145 0.700 ;
        RECT  2.965 0.825 3.130 0.895 ;
        RECT  2.100 0.995 3.130 1.065 ;
        RECT  2.895 0.350 2.965 0.895 ;
        RECT  2.685 0.825 2.895 0.895 ;
        RECT  2.650 0.205 2.720 0.470 ;
        RECT  1.965 0.545 2.720 0.615 ;
        RECT  2.615 0.685 2.685 0.925 ;
        RECT  2.320 0.400 2.650 0.470 ;
        RECT  2.160 0.685 2.615 0.755 ;
        RECT  2.050 0.840 2.530 0.910 ;
        RECT  2.225 0.375 2.320 0.470 ;
        RECT  2.040 0.375 2.225 0.445 ;
        RECT  1.980 0.995 2.100 1.075 ;
        RECT  1.965 0.225 2.060 0.295 ;
        RECT  1.895 0.225 1.965 0.915 ;
        RECT  1.755 0.205 1.825 0.430 ;
        RECT  0.685 0.985 1.810 1.055 ;
        RECT  0.610 0.205 1.755 0.275 ;
        RECT  1.680 0.545 1.740 0.615 ;
        RECT  1.610 0.350 1.680 0.905 ;
        RECT  1.540 0.350 1.610 0.420 ;
        RECT  1.510 0.835 1.610 0.905 ;
        RECT  1.410 0.520 1.530 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.820 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNCSND4BWP

MACRO SDFND0BWP
    CLASS CORE ;
    FOREIGN SDFND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.350 4.025 0.905 ;
        RECT  3.935 0.350 3.955 0.470 ;
        RECT  3.935 0.710 3.955 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.350 3.410 0.420 ;
        RECT  3.325 0.790 3.385 0.910 ;
        RECT  3.255 0.350 3.325 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.700 -0.115 3.820 0.140 ;
        RECT  3.200 -0.115 3.700 0.115 ;
        RECT  3.080 -0.115 3.200 0.130 ;
        RECT  2.360 -0.115 3.080 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 1.145 4.060 1.375 ;
        RECT  3.700 1.130 3.820 1.375 ;
        RECT  3.240 1.145 3.700 1.375 ;
        RECT  3.120 1.130 3.240 1.375 ;
        RECT  2.380 1.145 3.120 1.375 ;
        RECT  2.260 0.875 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.885 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.075 0.210 3.790 0.280 ;
        RECT  3.650 0.520 3.720 1.060 ;
        RECT  3.630 0.520 3.650 0.640 ;
        RECT  2.765 0.990 3.650 1.060 ;
        RECT  3.560 0.350 3.610 0.420 ;
        RECT  3.560 0.790 3.580 0.910 ;
        RECT  3.490 0.350 3.560 0.910 ;
        RECT  3.395 0.520 3.490 0.640 ;
        RECT  3.005 0.210 3.075 0.920 ;
        RECT  2.940 0.315 3.005 0.415 ;
        RECT  2.910 0.850 3.005 0.920 ;
        RECT  2.870 0.500 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.570 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.180 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  1.985 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  2.110 0.185 2.180 0.265 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.945 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.945 0.995 ;
        RECT  1.875 0.510 1.915 0.995 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.740 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFND0BWP

MACRO SDFND1BWP
    CLASS CORE ;
    FOREIGN SDFND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.045 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.735 3.955 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.350 3.410 0.420 ;
        RECT  3.325 0.790 3.385 0.910 ;
        RECT  3.255 0.350 3.325 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0150 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 -0.115 4.060 0.115 ;
        RECT  3.700 -0.115 3.820 0.140 ;
        RECT  3.200 -0.115 3.700 0.115 ;
        RECT  3.080 -0.115 3.200 0.130 ;
        RECT  2.360 -0.115 3.080 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.820 1.145 4.060 1.375 ;
        RECT  3.700 1.130 3.820 1.375 ;
        RECT  3.220 1.145 3.700 1.375 ;
        RECT  3.100 1.130 3.220 1.375 ;
        RECT  2.380 1.145 3.100 1.375 ;
        RECT  2.260 0.875 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.860 0.520 3.885 0.640 ;
        RECT  3.790 0.210 3.860 0.640 ;
        RECT  3.075 0.210 3.790 0.280 ;
        RECT  3.650 0.520 3.720 1.060 ;
        RECT  3.630 0.520 3.650 0.640 ;
        RECT  2.765 0.990 3.650 1.060 ;
        RECT  3.560 0.350 3.610 0.420 ;
        RECT  3.560 0.790 3.580 0.910 ;
        RECT  3.490 0.350 3.560 0.910 ;
        RECT  3.395 0.520 3.490 0.640 ;
        RECT  3.005 0.210 3.075 0.920 ;
        RECT  2.940 0.315 3.005 0.415 ;
        RECT  2.910 0.850 3.005 0.920 ;
        RECT  2.870 0.500 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.570 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.180 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  1.985 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  2.110 0.185 2.180 0.265 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.945 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.945 0.995 ;
        RECT  1.875 0.510 1.915 0.995 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFND1BWP

MACRO SDFND2BWP
    CLASS CORE ;
    FOREIGN SDFND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.355 4.305 0.805 ;
        RECT  4.235 0.185 4.245 1.035 ;
        RECT  4.175 0.185 4.235 0.465 ;
        RECT  4.175 0.735 4.235 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.350 3.885 0.910 ;
        RECT  3.795 0.350 3.815 0.470 ;
        RECT  3.795 0.770 3.815 0.910 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0150 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.300 ;
        RECT  4.080 -0.115 4.350 0.115 ;
        RECT  3.960 -0.115 4.080 0.140 ;
        RECT  3.650 -0.115 3.960 0.115 ;
        RECT  3.530 -0.115 3.650 0.140 ;
        RECT  3.260 -0.115 3.530 0.115 ;
        RECT  3.140 -0.115 3.260 0.140 ;
        RECT  2.360 -0.115 3.140 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.905 4.430 1.375 ;
        RECT  4.080 1.145 4.350 1.375 ;
        RECT  3.960 1.120 4.080 1.375 ;
        RECT  3.650 1.145 3.960 1.375 ;
        RECT  3.530 1.120 3.650 1.375 ;
        RECT  3.280 1.145 3.530 1.375 ;
        RECT  3.160 1.120 3.280 1.375 ;
        RECT  2.380 1.145 3.160 1.375 ;
        RECT  2.260 0.875 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.520 4.130 0.640 ;
        RECT  4.000 0.210 4.070 1.050 ;
        RECT  3.025 0.210 4.000 0.280 ;
        RECT  3.070 0.980 4.000 1.050 ;
        RECT  3.680 0.520 3.745 0.640 ;
        RECT  3.610 0.365 3.680 0.830 ;
        RECT  3.165 0.365 3.610 0.435 ;
        RECT  3.445 0.760 3.610 0.830 ;
        RECT  3.375 0.760 3.445 0.900 ;
        RECT  3.305 0.545 3.400 0.615 ;
        RECT  3.235 0.545 3.305 0.910 ;
        RECT  2.765 0.840 3.235 0.910 ;
        RECT  3.095 0.365 3.165 0.615 ;
        RECT  3.040 0.545 3.095 0.615 ;
        RECT  2.950 0.980 3.070 1.075 ;
        RECT  2.955 0.185 3.025 0.465 ;
        RECT  2.870 0.580 2.935 0.770 ;
        RECT  2.865 0.195 2.870 0.770 ;
        RECT  2.800 0.195 2.865 0.650 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.180 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  1.985 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  2.110 0.185 2.180 0.265 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.945 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.945 0.995 ;
        RECT  1.875 0.510 1.915 0.995 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFND2BWP

MACRO SDFND4BWP
    CLASS CORE ;
    FOREIGN SDFND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.775 4.945 1.065 ;
        RECT  4.795 0.355 4.875 0.465 ;
        RECT  4.795 0.775 4.875 0.905 ;
        RECT  4.585 0.355 4.795 0.905 ;
        RECT  4.565 0.355 4.585 0.465 ;
        RECT  4.495 0.775 4.585 1.075 ;
        RECT  4.495 0.185 4.565 0.465 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.710 4.230 0.800 ;
        RECT  4.095 0.355 4.210 0.445 ;
        RECT  3.885 0.355 4.095 0.800 ;
        RECT  3.710 0.355 3.885 0.445 ;
        RECT  3.750 0.710 3.885 0.800 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.055 -0.115 5.125 0.465 ;
        RECT  4.755 -0.115 5.055 0.115 ;
        RECT  4.685 -0.115 4.755 0.285 ;
        RECT  4.400 -0.115 4.685 0.115 ;
        RECT  4.280 -0.115 4.400 0.145 ;
        RECT  4.020 -0.115 4.280 0.115 ;
        RECT  3.900 -0.115 4.020 0.145 ;
        RECT  3.640 -0.115 3.900 0.115 ;
        RECT  3.520 -0.115 3.640 0.145 ;
        RECT  3.260 -0.115 3.520 0.115 ;
        RECT  3.140 -0.115 3.260 0.145 ;
        RECT  2.380 -0.115 3.140 0.115 ;
        RECT  2.260 -0.115 2.380 0.125 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.055 0.685 5.125 1.375 ;
        RECT  4.755 1.145 5.055 1.375 ;
        RECT  4.685 0.975 4.755 1.375 ;
        RECT  4.410 1.145 4.685 1.375 ;
        RECT  4.290 1.010 4.410 1.375 ;
        RECT  4.050 1.145 4.290 1.375 ;
        RECT  3.930 1.010 4.050 1.375 ;
        RECT  3.680 1.145 3.930 1.375 ;
        RECT  3.560 1.010 3.680 1.375 ;
        RECT  3.300 1.145 3.560 1.375 ;
        RECT  3.180 1.130 3.300 1.375 ;
        RECT  2.400 1.145 3.180 1.375 ;
        RECT  2.280 0.870 2.400 1.375 ;
        RECT  1.440 1.145 2.280 1.375 ;
        RECT  1.320 1.120 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.120 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.875 0.185 4.945 0.465 ;
        RECT  4.875 0.775 4.945 1.065 ;
        RECT  4.865 0.355 4.875 0.465 ;
        RECT  4.865 0.775 4.875 0.905 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.775 4.515 1.075 ;
        RECT  4.165 0.710 4.230 0.800 ;
        RECT  4.165 0.355 4.210 0.445 ;
        RECT  3.710 0.355 3.815 0.445 ;
        RECT  3.750 0.710 3.815 0.800 ;
        RECT  4.370 0.545 4.490 0.615 ;
        RECT  4.300 0.215 4.370 0.940 ;
        RECT  3.030 0.215 4.300 0.285 ;
        RECT  3.475 0.870 4.300 0.940 ;
        RECT  3.600 0.545 3.780 0.615 ;
        RECT  3.530 0.365 3.600 0.800 ;
        RECT  3.170 0.365 3.530 0.435 ;
        RECT  3.380 0.700 3.530 0.800 ;
        RECT  3.405 0.870 3.475 1.060 ;
        RECT  3.310 0.545 3.450 0.615 ;
        RECT  2.920 0.990 3.405 1.060 ;
        RECT  3.240 0.545 3.310 0.920 ;
        RECT  2.795 0.850 3.240 0.920 ;
        RECT  3.100 0.365 3.170 0.630 ;
        RECT  3.070 0.530 3.100 0.630 ;
        RECT  2.960 0.215 3.030 0.425 ;
        RECT  2.890 0.710 3.000 0.780 ;
        RECT  2.820 0.195 2.890 0.780 ;
        RECT  2.700 0.195 2.820 0.265 ;
        RECT  2.750 0.850 2.795 1.070 ;
        RECT  2.725 0.350 2.750 1.070 ;
        RECT  2.680 0.350 2.725 0.920 ;
        RECT  2.580 0.185 2.700 0.265 ;
        RECT  2.540 0.355 2.610 1.040 ;
        RECT  2.180 0.195 2.580 0.265 ;
        RECT  2.470 0.355 2.540 0.425 ;
        RECT  2.535 0.730 2.540 1.040 ;
        RECT  2.275 0.730 2.535 0.800 ;
        RECT  2.400 0.510 2.470 0.640 ;
        RECT  2.005 0.510 2.400 0.580 ;
        RECT  2.205 0.650 2.275 0.800 ;
        RECT  2.110 0.185 2.180 0.265 ;
        RECT  2.020 0.185 2.110 0.255 ;
        RECT  1.965 0.325 2.005 0.580 ;
        RECT  1.935 0.325 1.965 0.990 ;
        RECT  1.895 0.510 1.935 0.990 ;
        RECT  1.755 0.200 1.825 0.430 ;
        RECT  0.685 0.980 1.815 1.050 ;
        RECT  1.680 0.565 1.810 0.635 ;
        RECT  0.610 0.200 1.755 0.270 ;
        RECT  1.610 0.340 1.680 0.910 ;
        RECT  1.540 0.340 1.610 0.410 ;
        RECT  1.510 0.840 1.610 0.910 ;
        RECT  1.410 0.520 1.530 0.640 ;
        RECT  1.340 0.340 1.410 0.910 ;
        RECT  1.170 0.340 1.340 0.410 ;
        RECT  1.120 0.840 1.340 0.910 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.840 0.900 0.910 ;
        RECT  0.760 0.350 0.830 0.910 ;
        RECT  0.615 0.790 0.685 1.050 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFND4BWP

MACRO SDFNSND0BWP
    CLASS CORE ;
    FOREIGN SDFNSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.195 4.585 0.905 ;
        RECT  4.495 0.195 4.515 0.315 ;
        RECT  4.495 0.755 4.515 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.210 0.350 4.280 0.775 ;
        RECT  4.095 0.350 4.210 0.470 ;
        RECT  4.185 0.695 4.210 0.775 ;
        RECT  4.095 0.695 4.185 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  2.380 -0.115 4.280 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.845 4.400 1.375 ;
        RECT  3.820 1.145 4.280 1.375 ;
        RECT  3.700 1.135 3.820 1.375 ;
        RECT  3.460 1.145 3.700 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.240 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.640 ;
        RECT  4.355 0.210 4.425 0.640 ;
        RECT  3.450 0.210 4.355 0.280 ;
        RECT  4.010 0.545 4.130 0.615 ;
        RECT  3.940 0.350 4.010 1.045 ;
        RECT  3.600 0.975 3.940 1.045 ;
        RECT  3.800 0.520 3.870 0.905 ;
        RECT  3.085 0.835 3.800 0.905 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.180 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.905 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.160 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.235 0.710 2.675 0.780 ;
        RECT  2.385 0.510 2.455 0.640 ;
        RECT  1.985 0.510 2.385 0.580 ;
        RECT  2.165 0.650 2.235 0.780 ;
        RECT  2.110 0.185 2.180 0.275 ;
        RECT  2.090 0.850 2.160 1.075 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.980 1.005 2.090 1.075 ;
        RECT  1.965 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.965 0.930 ;
        RECT  1.895 0.510 1.915 0.930 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.740 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.905 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.835 1.590 0.905 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.905 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.835 1.340 0.905 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFNSND0BWP

MACRO SDFNSND1BWP
    CLASS CORE ;
    FOREIGN SDFNSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.585 1.045 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.730 4.515 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.210 0.350 4.280 0.775 ;
        RECT  4.095 0.350 4.210 0.470 ;
        RECT  4.185 0.695 4.210 0.775 ;
        RECT  4.095 0.695 4.185 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  2.380 -0.115 4.280 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.375 1.145 4.620 1.375 ;
        RECT  4.305 0.895 4.375 1.375 ;
        RECT  3.820 1.145 4.305 1.375 ;
        RECT  3.700 1.135 3.820 1.375 ;
        RECT  3.460 1.145 3.700 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.240 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.640 ;
        RECT  4.355 0.210 4.425 0.640 ;
        RECT  3.450 0.210 4.355 0.280 ;
        RECT  4.010 0.545 4.130 0.615 ;
        RECT  3.940 0.350 4.010 1.045 ;
        RECT  3.600 0.975 3.940 1.045 ;
        RECT  3.800 0.520 3.870 0.905 ;
        RECT  3.085 0.835 3.800 0.905 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.180 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.905 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.160 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.235 0.710 2.675 0.780 ;
        RECT  2.385 0.510 2.455 0.640 ;
        RECT  1.985 0.510 2.385 0.580 ;
        RECT  2.165 0.650 2.235 0.780 ;
        RECT  2.110 0.185 2.180 0.275 ;
        RECT  2.090 0.850 2.160 1.075 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.980 1.005 2.090 1.075 ;
        RECT  1.965 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.965 0.930 ;
        RECT  1.895 0.510 1.915 0.930 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.915 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.845 1.590 0.915 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNSND1BWP

MACRO SDFNSND2BWP
    CLASS CORE ;
    FOREIGN SDFNSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.805 0.355 4.865 0.815 ;
        RECT  4.795 0.185 4.805 1.035 ;
        RECT  4.735 0.185 4.795 0.465 ;
        RECT  4.735 0.745 4.795 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.350 4.445 1.045 ;
        RECT  4.360 0.350 4.375 0.480 ;
        RECT  4.355 0.745 4.375 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.300 ;
        RECT  4.640 -0.115 4.910 0.115 ;
        RECT  4.520 -0.115 4.640 0.140 ;
        RECT  4.250 -0.115 4.520 0.115 ;
        RECT  4.130 -0.115 4.250 0.140 ;
        RECT  3.850 -0.115 4.130 0.115 ;
        RECT  3.730 -0.115 3.850 0.140 ;
        RECT  2.380 -0.115 3.730 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.905 4.990 1.375 ;
        RECT  4.615 1.145 4.910 1.375 ;
        RECT  4.545 0.735 4.615 1.375 ;
        RECT  4.250 1.145 4.545 1.375 ;
        RECT  4.130 1.120 4.250 1.375 ;
        RECT  3.865 1.145 4.130 1.375 ;
        RECT  3.795 0.980 3.865 1.375 ;
        RECT  3.460 1.145 3.795 1.375 ;
        RECT  3.340 1.015 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.240 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.240 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.630 0.545 4.720 0.615 ;
        RECT  4.560 0.210 4.630 0.615 ;
        RECT  3.450 0.210 4.560 0.280 ;
        RECT  4.230 0.520 4.300 0.640 ;
        RECT  4.160 0.365 4.230 1.050 ;
        RECT  3.765 0.365 4.160 0.435 ;
        RECT  3.950 0.980 4.160 1.050 ;
        RECT  3.905 0.520 3.975 0.910 ;
        RECT  3.085 0.840 3.905 0.910 ;
        RECT  3.695 0.365 3.765 0.640 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.180 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.910 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.160 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.235 0.710 2.675 0.780 ;
        RECT  2.385 0.510 2.455 0.640 ;
        RECT  1.985 0.510 2.385 0.580 ;
        RECT  2.165 0.650 2.235 0.780 ;
        RECT  2.110 0.185 2.180 0.275 ;
        RECT  2.090 0.850 2.160 1.075 ;
        RECT  2.000 0.185 2.110 0.255 ;
        RECT  1.980 1.005 2.090 1.075 ;
        RECT  1.965 0.325 1.985 0.580 ;
        RECT  1.915 0.325 1.965 0.930 ;
        RECT  1.895 0.510 1.915 0.930 ;
        RECT  1.735 0.195 1.805 0.430 ;
        RECT  1.660 0.565 1.790 0.635 ;
        RECT  0.685 0.985 1.790 1.055 ;
        RECT  0.610 0.195 1.735 0.265 ;
        RECT  1.590 0.350 1.660 0.915 ;
        RECT  1.520 0.350 1.590 0.420 ;
        RECT  1.490 0.845 1.590 0.915 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNSND2BWP

MACRO SDFNSND4BWP
    CLASS CORE ;
    FOREIGN SDFNSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.640 ;
        RECT  3.470 0.520 3.535 0.640 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.185 5.505 0.465 ;
        RECT  5.495 0.765 5.505 1.065 ;
        RECT  5.435 0.185 5.495 1.065 ;
        RECT  5.285 0.355 5.435 0.905 ;
        RECT  5.145 0.355 5.285 0.465 ;
        RECT  5.145 0.765 5.285 0.905 ;
        RECT  5.075 0.185 5.145 0.465 ;
        RECT  5.075 0.765 5.145 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.355 4.790 0.455 ;
        RECT  4.695 0.765 4.765 1.065 ;
        RECT  4.655 0.765 4.695 0.905 ;
        RECT  4.445 0.355 4.655 0.905 ;
        RECT  4.290 0.355 4.445 0.455 ;
        RECT  4.385 0.765 4.445 0.905 ;
        RECT  4.315 0.765 4.385 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.465 ;
        RECT  5.350 -0.115 5.610 0.115 ;
        RECT  5.230 -0.115 5.350 0.275 ;
        RECT  4.980 -0.115 5.230 0.115 ;
        RECT  4.860 -0.115 4.980 0.140 ;
        RECT  4.600 -0.115 4.860 0.115 ;
        RECT  4.480 -0.115 4.600 0.140 ;
        RECT  4.220 -0.115 4.480 0.115 ;
        RECT  4.100 -0.115 4.220 0.140 ;
        RECT  3.840 -0.115 4.100 0.115 ;
        RECT  3.720 -0.115 3.840 0.140 ;
        RECT  2.380 -0.115 3.720 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.135 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.685 5.690 1.375 ;
        RECT  5.325 1.145 5.610 1.375 ;
        RECT  5.255 0.975 5.325 1.375 ;
        RECT  4.945 1.145 5.255 1.375 ;
        RECT  4.875 0.745 4.945 1.375 ;
        RECT  4.590 1.145 4.875 1.375 ;
        RECT  4.490 0.985 4.590 1.375 ;
        RECT  4.220 1.145 4.490 1.375 ;
        RECT  4.100 1.110 4.220 1.375 ;
        RECT  3.850 1.145 4.100 1.375 ;
        RECT  3.730 1.005 3.850 1.375 ;
        RECT  3.490 1.145 3.730 1.375 ;
        RECT  3.370 1.005 3.490 1.375 ;
        RECT  2.750 1.145 3.370 1.375 ;
        RECT  2.630 0.990 2.750 1.375 ;
        RECT  2.390 1.145 2.630 1.375 ;
        RECT  2.260 1.005 2.390 1.375 ;
        RECT  1.440 1.145 2.260 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.145 0.355 5.215 0.465 ;
        RECT  5.145 0.765 5.215 0.905 ;
        RECT  5.075 0.185 5.145 0.465 ;
        RECT  5.075 0.765 5.145 1.065 ;
        RECT  4.725 0.355 4.790 0.455 ;
        RECT  4.725 0.765 4.765 1.065 ;
        RECT  4.290 0.355 4.375 0.455 ;
        RECT  4.315 0.765 4.375 1.065 ;
        RECT  4.950 0.545 5.110 0.615 ;
        RECT  4.880 0.210 4.950 0.615 ;
        RECT  3.450 0.210 4.880 0.280 ;
        RECT  4.200 0.545 4.325 0.615 ;
        RECT  4.130 0.365 4.200 0.990 ;
        RECT  3.755 0.365 4.130 0.435 ;
        RECT  3.920 0.890 4.130 0.990 ;
        RECT  3.935 0.520 4.005 0.810 ;
        RECT  3.820 0.740 3.935 0.810 ;
        RECT  3.750 0.740 3.820 0.935 ;
        RECT  3.685 0.365 3.755 0.640 ;
        RECT  3.085 0.865 3.750 0.935 ;
        RECT  3.230 0.720 3.670 0.790 ;
        RECT  3.330 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.330 0.425 ;
        RECT  2.200 0.205 3.260 0.275 ;
        RECT  3.160 0.355 3.230 0.790 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.935 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.835 0.850 2.905 1.060 ;
        RECT  2.180 0.850 2.835 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.255 0.710 2.675 0.780 ;
        RECT  2.405 0.510 2.475 0.640 ;
        RECT  2.005 0.510 2.405 0.580 ;
        RECT  2.185 0.650 2.255 0.780 ;
        RECT  2.130 0.185 2.200 0.275 ;
        RECT  2.110 0.850 2.180 1.075 ;
        RECT  2.020 0.185 2.130 0.255 ;
        RECT  2.000 1.005 2.110 1.075 ;
        RECT  1.985 0.325 2.005 0.580 ;
        RECT  1.935 0.325 1.985 0.930 ;
        RECT  1.915 0.510 1.935 0.930 ;
        RECT  1.755 0.205 1.825 0.430 ;
        RECT  1.680 0.565 1.810 0.635 ;
        RECT  0.685 0.985 1.810 1.055 ;
        RECT  0.610 0.205 1.755 0.275 ;
        RECT  1.610 0.350 1.680 0.915 ;
        RECT  1.540 0.350 1.610 0.420 ;
        RECT  1.510 0.845 1.610 0.915 ;
        RECT  1.410 0.520 1.530 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFNSND4BWP

MACRO SDFQD0BWP
    CLASS CORE ;
    FOREIGN SDFQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.195 3.745 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.635 0.945 0.905 ;
        RECT  0.805 0.635 0.875 0.765 ;
        RECT  0.735 0.570 0.805 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.520 1.175 0.705 ;
        RECT  1.085 0.635 1.105 0.705 ;
        RECT  1.015 0.635 1.085 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 -0.115 3.780 0.115 ;
        RECT  3.475 -0.115 3.545 0.295 ;
        RECT  3.220 -0.115 3.475 0.115 ;
        RECT  3.100 -0.115 3.220 0.145 ;
        RECT  2.440 -0.115 3.100 0.115 ;
        RECT  2.315 -0.115 2.440 0.120 ;
        RECT  1.670 -0.115 2.315 0.115 ;
        RECT  1.550 -0.115 1.670 0.300 ;
        RECT  1.070 -0.115 1.550 0.115 ;
        RECT  0.950 -0.115 1.070 0.240 ;
        RECT  0.340 -0.115 0.950 0.115 ;
        RECT  0.210 -0.115 0.340 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.145 3.780 1.375 ;
        RECT  3.450 1.005 3.570 1.375 ;
        RECT  3.240 1.145 3.450 1.375 ;
        RECT  3.120 1.135 3.240 1.375 ;
        RECT  2.460 1.145 3.120 1.375 ;
        RECT  2.340 0.860 2.460 1.375 ;
        RECT  1.700 1.145 2.340 1.375 ;
        RECT  1.580 1.040 1.700 1.375 ;
        RECT  1.120 1.145 1.580 1.375 ;
        RECT  1.000 1.125 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.210 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.515 0.375 3.585 0.935 ;
        RECT  3.115 0.375 3.515 0.445 ;
        RECT  3.270 0.865 3.515 0.935 ;
        RECT  3.365 0.520 3.435 0.790 ;
        RECT  3.125 0.720 3.365 0.790 ;
        RECT  3.055 0.720 3.125 1.060 ;
        RECT  3.045 0.375 3.115 0.640 ;
        RECT  2.780 0.990 3.055 1.060 ;
        RECT  2.885 0.200 2.955 0.920 ;
        RECT  2.760 0.200 2.885 0.270 ;
        RECT  2.855 0.800 2.885 0.920 ;
        RECT  2.780 0.350 2.805 0.470 ;
        RECT  2.710 0.350 2.780 1.060 ;
        RECT  2.640 0.185 2.760 0.270 ;
        RECT  1.820 0.200 2.640 0.270 ;
        RECT  2.560 0.350 2.630 1.065 ;
        RECT  2.555 0.720 2.560 1.065 ;
        RECT  2.315 0.720 2.555 0.790 ;
        RECT  2.420 0.350 2.490 0.640 ;
        RECT  2.065 0.350 2.420 0.420 ;
        RECT  2.245 0.520 2.315 0.790 ;
        RECT  1.995 0.350 2.065 0.950 ;
        RECT  1.750 0.200 1.820 0.440 ;
        RECT  1.705 0.520 1.775 0.965 ;
        RECT  1.630 0.370 1.750 0.440 ;
        RECT  1.480 0.895 1.705 0.965 ;
        RECT  1.560 0.370 1.630 0.825 ;
        RECT  1.465 0.370 1.560 0.440 ;
        RECT  1.395 0.705 1.560 0.825 ;
        RECT  1.320 0.545 1.490 0.615 ;
        RECT  1.410 0.895 1.480 1.055 ;
        RECT  1.395 0.235 1.465 0.440 ;
        RECT  0.795 0.985 1.410 1.055 ;
        RECT  1.250 0.315 1.320 0.905 ;
        RECT  1.190 0.315 1.250 0.385 ;
        RECT  1.180 0.835 1.250 0.905 ;
        RECT  0.915 0.310 0.985 0.560 ;
        RECT  0.840 0.310 0.915 0.380 ;
        RECT  0.770 0.195 0.840 0.380 ;
        RECT  0.725 0.835 0.795 1.055 ;
        RECT  0.525 0.195 0.770 0.265 ;
        RECT  0.665 0.835 0.725 0.905 ;
        RECT  0.665 0.335 0.685 0.455 ;
        RECT  0.595 0.335 0.665 0.905 ;
        RECT  0.525 0.985 0.625 1.055 ;
        RECT  0.455 0.195 0.525 1.055 ;
        RECT  0.125 0.355 0.455 0.425 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFQD0BWP

MACRO SDFQD1BWP
    CLASS CORE ;
    FOREIGN SDFQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.195 3.745 1.070 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 -0.115 3.780 0.115 ;
        RECT  3.475 -0.115 3.545 0.315 ;
        RECT  3.185 -0.115 3.475 0.115 ;
        RECT  3.115 -0.115 3.185 0.315 ;
        RECT  2.360 -0.115 3.115 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 1.145 3.780 1.375 ;
        RECT  3.475 0.895 3.545 1.375 ;
        RECT  3.180 1.145 3.475 1.375 ;
        RECT  3.060 1.130 3.180 1.375 ;
        RECT  2.380 1.145 3.060 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.435 0.395 3.505 0.810 ;
        RECT  3.365 0.395 3.435 0.465 ;
        RECT  3.365 0.740 3.435 0.810 ;
        RECT  3.295 0.185 3.365 0.465 ;
        RECT  3.295 0.740 3.365 1.025 ;
        RECT  3.225 0.545 3.320 0.615 ;
        RECT  3.075 0.395 3.295 0.465 ;
        RECT  3.155 0.545 3.225 0.930 ;
        RECT  2.765 0.860 3.155 0.930 ;
        RECT  3.005 0.395 3.075 0.600 ;
        RECT  2.865 0.195 2.935 0.780 ;
        RECT  2.680 0.195 2.865 0.265 ;
        RECT  2.695 0.350 2.765 1.060 ;
        RECT  2.660 0.350 2.695 0.470 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQD1BWP

MACRO SDFQD2BWP
    CLASS CORE ;
    FOREIGN SDFQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.685 0.355 3.745 0.805 ;
        RECT  3.675 0.185 3.685 1.035 ;
        RECT  3.615 0.185 3.675 0.465 ;
        RECT  3.615 0.735 3.675 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.300 ;
        RECT  3.505 -0.115 3.790 0.115 ;
        RECT  3.435 -0.115 3.505 0.465 ;
        RECT  3.170 -0.115 3.435 0.115 ;
        RECT  3.050 -0.115 3.170 0.280 ;
        RECT  2.360 -0.115 3.050 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.925 3.870 1.375 ;
        RECT  3.505 1.145 3.790 1.375 ;
        RECT  3.435 0.735 3.505 1.375 ;
        RECT  3.160 1.145 3.435 1.375 ;
        RECT  3.040 1.130 3.160 1.375 ;
        RECT  2.380 1.145 3.040 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.360 0.545 3.600 0.615 ;
        RECT  3.325 0.370 3.360 1.035 ;
        RECT  3.290 0.185 3.325 1.035 ;
        RECT  3.255 0.185 3.290 0.440 ;
        RECT  3.255 0.735 3.290 1.035 ;
        RECT  3.015 0.370 3.255 0.440 ;
        RECT  3.180 0.520 3.215 0.640 ;
        RECT  3.110 0.520 3.180 1.060 ;
        RECT  2.730 0.990 3.110 1.060 ;
        RECT  2.945 0.370 3.015 0.640 ;
        RECT  2.800 0.195 2.870 0.910 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.660 0.350 2.730 1.060 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.565 0.355 2.590 0.800 ;
        RECT  2.520 0.355 2.565 1.050 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.495 0.730 2.520 1.050 ;
        RECT  2.255 0.730 2.495 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.865 1.790 0.935 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.865 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQD2BWP

MACRO SDFQD4BWP
    CLASS CORE ;
    FOREIGN SDFQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.105 0.465 ;
        RECT  4.095 0.765 4.105 1.065 ;
        RECT  4.035 0.185 4.095 1.065 ;
        RECT  3.885 0.355 4.035 0.905 ;
        RECT  3.745 0.355 3.885 0.465 ;
        RECT  3.745 0.765 3.885 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.115 4.340 0.115 ;
        RECT  4.215 -0.115 4.285 0.465 ;
        RECT  3.950 -0.115 4.215 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.565 -0.115 3.830 0.115 ;
        RECT  3.495 -0.115 3.565 0.465 ;
        RECT  3.230 -0.115 3.495 0.115 ;
        RECT  3.110 -0.115 3.230 0.280 ;
        RECT  2.380 -0.115 3.110 0.115 ;
        RECT  2.260 -0.115 2.380 0.125 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 1.145 4.340 1.375 ;
        RECT  4.215 0.675 4.285 1.375 ;
        RECT  3.925 1.145 4.215 1.375 ;
        RECT  3.855 0.975 3.925 1.375 ;
        RECT  3.565 1.145 3.855 1.375 ;
        RECT  3.495 0.735 3.565 1.375 ;
        RECT  3.195 1.145 3.495 1.375 ;
        RECT  3.125 0.970 3.195 1.375 ;
        RECT  2.400 1.145 3.125 1.375 ;
        RECT  2.280 0.870 2.400 1.375 ;
        RECT  1.440 1.145 2.280 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.355 3.815 0.465 ;
        RECT  3.745 0.765 3.815 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        RECT  3.420 0.545 3.710 0.615 ;
        RECT  3.385 0.370 3.420 1.035 ;
        RECT  3.350 0.185 3.385 1.035 ;
        RECT  3.315 0.185 3.350 0.440 ;
        RECT  3.315 0.735 3.350 1.035 ;
        RECT  3.075 0.370 3.315 0.440 ;
        RECT  3.220 0.520 3.275 0.640 ;
        RECT  3.150 0.520 3.220 0.890 ;
        RECT  3.045 0.820 3.150 0.890 ;
        RECT  3.005 0.370 3.075 0.640 ;
        RECT  2.975 0.820 3.045 1.060 ;
        RECT  2.750 0.990 2.975 1.060 ;
        RECT  2.825 0.195 2.895 0.910 ;
        RECT  2.700 0.195 2.825 0.265 ;
        RECT  2.680 0.350 2.750 1.060 ;
        RECT  2.580 0.185 2.700 0.265 ;
        RECT  2.540 0.355 2.610 1.060 ;
        RECT  2.040 0.195 2.580 0.265 ;
        RECT  2.470 0.355 2.540 0.425 ;
        RECT  2.535 0.730 2.540 1.060 ;
        RECT  2.275 0.730 2.535 0.800 ;
        RECT  2.400 0.510 2.470 0.640 ;
        RECT  2.025 0.510 2.400 0.580 ;
        RECT  2.205 0.650 2.275 0.800 ;
        RECT  1.965 0.350 2.025 0.580 ;
        RECT  1.955 0.350 1.965 0.950 ;
        RECT  1.895 0.510 1.955 0.950 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.655 0.350 1.725 0.795 ;
        RECT  1.540 0.350 1.655 0.420 ;
        RECT  1.510 0.725 1.655 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQD4BWP

MACRO SDFQND0BWP
    CLASS CORE ;
    FOREIGN SDFQND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNAGATEAREA 0.0096 ;
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.215 3.465 1.045 ;
        RECT  3.375 0.215 3.395 0.450 ;
        RECT  3.375 0.735 3.395 1.045 ;
        RECT  3.135 0.380 3.375 0.450 ;
        RECT  3.065 0.380 3.135 0.640 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 -0.115 3.500 0.115 ;
        RECT  3.195 -0.115 3.265 0.305 ;
        RECT  2.360 -0.115 3.195 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.145 3.500 1.375 ;
        RECT  3.140 1.130 3.260 1.375 ;
        RECT  2.380 1.145 3.140 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.305 0.520 3.325 0.640 ;
        RECT  3.235 0.520 3.305 1.060 ;
        RECT  2.765 0.990 3.235 1.060 ;
        RECT  2.875 0.195 2.945 0.840 ;
        RECT  2.680 0.195 2.875 0.265 ;
        RECT  2.730 0.730 2.765 1.060 ;
        RECT  2.695 0.350 2.730 1.060 ;
        RECT  2.660 0.350 2.695 0.800 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.480 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFQND0BWP

MACRO SDFQND1BWP
    CLASS CORE ;
    FOREIGN SDFQND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.195 3.745 1.070 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 -0.115 3.780 0.115 ;
        RECT  3.450 -0.115 3.570 0.280 ;
        RECT  3.175 -0.115 3.450 0.115 ;
        RECT  3.105 -0.115 3.175 0.285 ;
        RECT  2.360 -0.115 3.105 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 1.145 3.780 1.375 ;
        RECT  3.475 0.895 3.545 1.375 ;
        RECT  3.220 1.145 3.475 1.375 ;
        RECT  3.100 1.125 3.220 1.375 ;
        RECT  2.380 1.145 3.100 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.435 0.355 3.505 0.810 ;
        RECT  3.075 0.355 3.435 0.425 ;
        RECT  3.365 0.740 3.435 0.810 ;
        RECT  3.295 0.740 3.365 0.950 ;
        RECT  3.225 0.545 3.340 0.615 ;
        RECT  3.155 0.545 3.225 0.930 ;
        RECT  2.765 0.860 3.155 0.930 ;
        RECT  3.005 0.355 3.075 0.600 ;
        RECT  2.865 0.195 2.935 0.780 ;
        RECT  2.680 0.195 2.865 0.265 ;
        RECT  2.695 0.350 2.765 1.060 ;
        RECT  2.660 0.350 2.695 0.470 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.520 0.355 2.590 1.060 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.515 0.730 2.520 1.060 ;
        RECT  2.255 0.730 2.515 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQND1BWP

MACRO SDFQND2BWP
    CLASS CORE ;
    FOREIGN SDFQND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.685 0.355 3.745 0.805 ;
        RECT  3.675 0.185 3.685 1.035 ;
        RECT  3.615 0.185 3.675 0.465 ;
        RECT  3.615 0.735 3.675 1.035 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.300 ;
        RECT  3.505 -0.115 3.790 0.115 ;
        RECT  3.435 -0.115 3.505 0.465 ;
        RECT  3.135 -0.115 3.435 0.115 ;
        RECT  3.065 -0.115 3.135 0.285 ;
        RECT  2.360 -0.115 3.065 0.115 ;
        RECT  2.240 -0.115 2.360 0.125 ;
        RECT  1.440 -0.115 2.240 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.925 3.870 1.375 ;
        RECT  3.505 1.145 3.790 1.375 ;
        RECT  3.435 0.675 3.505 1.375 ;
        RECT  3.160 1.145 3.435 1.375 ;
        RECT  3.040 1.130 3.160 1.375 ;
        RECT  2.380 1.145 3.040 1.375 ;
        RECT  2.260 0.870 2.380 1.375 ;
        RECT  1.400 1.145 2.260 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.290 0.355 3.360 1.070 ;
        RECT  3.015 0.355 3.290 0.425 ;
        RECT  3.255 0.950 3.290 1.070 ;
        RECT  3.180 0.520 3.215 0.640 ;
        RECT  3.110 0.520 3.180 1.060 ;
        RECT  2.730 0.990 3.110 1.060 ;
        RECT  2.945 0.355 3.015 0.640 ;
        RECT  2.800 0.195 2.870 0.910 ;
        RECT  2.680 0.195 2.800 0.265 ;
        RECT  2.660 0.350 2.730 1.060 ;
        RECT  2.560 0.185 2.680 0.265 ;
        RECT  2.565 0.355 2.590 0.800 ;
        RECT  2.520 0.355 2.565 1.050 ;
        RECT  2.020 0.195 2.560 0.265 ;
        RECT  2.450 0.355 2.520 0.425 ;
        RECT  2.495 0.730 2.520 1.050 ;
        RECT  2.255 0.730 2.495 0.800 ;
        RECT  2.380 0.510 2.450 0.640 ;
        RECT  2.005 0.510 2.380 0.580 ;
        RECT  2.185 0.650 2.255 0.800 ;
        RECT  1.945 0.350 2.005 0.580 ;
        RECT  1.935 0.350 1.945 0.950 ;
        RECT  1.875 0.510 1.935 0.950 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.610 0.875 1.790 0.945 ;
        RECT  1.635 0.350 1.705 0.795 ;
        RECT  1.520 0.350 1.635 0.420 ;
        RECT  1.490 0.725 1.635 0.795 ;
        RECT  1.540 0.875 1.610 1.055 ;
        RECT  0.685 0.985 1.540 1.055 ;
        RECT  1.410 0.520 1.515 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQND2BWP

MACRO SDFQND4BWP
    CLASS CORE ;
    FOREIGN SDFQND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.105 0.465 ;
        RECT  4.095 0.765 4.105 1.065 ;
        RECT  4.035 0.185 4.095 1.065 ;
        RECT  3.885 0.355 4.035 0.905 ;
        RECT  3.745 0.355 3.885 0.465 ;
        RECT  3.745 0.765 3.885 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.465 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.275 ;
        RECT  3.565 -0.115 3.830 0.115 ;
        RECT  3.495 -0.115 3.565 0.465 ;
        RECT  3.195 -0.115 3.495 0.115 ;
        RECT  3.125 -0.115 3.195 0.305 ;
        RECT  2.380 -0.115 3.125 0.115 ;
        RECT  2.260 -0.115 2.380 0.125 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.685 4.290 1.375 ;
        RECT  3.925 1.145 4.210 1.375 ;
        RECT  3.855 0.975 3.925 1.375 ;
        RECT  3.565 1.145 3.855 1.375 ;
        RECT  3.495 0.675 3.565 1.375 ;
        RECT  3.195 1.145 3.495 1.375 ;
        RECT  3.125 0.950 3.195 1.375 ;
        RECT  2.400 1.145 3.125 1.375 ;
        RECT  2.280 0.870 2.400 1.375 ;
        RECT  1.440 1.145 2.280 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.355 3.815 0.465 ;
        RECT  3.745 0.765 3.815 0.905 ;
        RECT  3.675 0.185 3.745 0.465 ;
        RECT  3.675 0.765 3.745 1.065 ;
        RECT  3.355 0.375 3.425 1.045 ;
        RECT  3.075 0.375 3.355 0.445 ;
        RECT  3.290 0.975 3.355 1.045 ;
        RECT  3.205 0.520 3.275 0.870 ;
        RECT  3.045 0.800 3.205 0.870 ;
        RECT  3.005 0.375 3.075 0.640 ;
        RECT  2.975 0.800 3.045 1.060 ;
        RECT  2.750 0.990 2.975 1.060 ;
        RECT  2.825 0.195 2.895 0.910 ;
        RECT  2.700 0.195 2.825 0.265 ;
        RECT  2.680 0.350 2.750 1.060 ;
        RECT  2.580 0.185 2.700 0.265 ;
        RECT  2.540 0.355 2.610 1.060 ;
        RECT  2.040 0.195 2.580 0.265 ;
        RECT  2.470 0.355 2.540 0.425 ;
        RECT  2.535 0.730 2.540 1.060 ;
        RECT  2.275 0.730 2.535 0.800 ;
        RECT  2.400 0.510 2.470 0.640 ;
        RECT  2.025 0.510 2.400 0.580 ;
        RECT  2.205 0.650 2.275 0.800 ;
        RECT  1.965 0.350 2.025 0.580 ;
        RECT  1.955 0.350 1.965 0.950 ;
        RECT  1.895 0.510 1.955 0.950 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.655 0.350 1.725 0.795 ;
        RECT  1.540 0.350 1.655 0.420 ;
        RECT  1.510 0.725 1.655 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFQND4BWP

MACRO SDFSND0BWP
    CLASS CORE ;
    FOREIGN SDFSND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.490 0.500 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.195 4.585 0.905 ;
        RECT  4.495 0.195 4.515 0.315 ;
        RECT  4.495 0.755 4.515 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.210 0.350 4.280 0.775 ;
        RECT  4.095 0.350 4.210 0.470 ;
        RECT  4.185 0.695 4.210 0.775 ;
        RECT  4.095 0.695 4.185 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  3.840 -0.115 4.280 0.115 ;
        RECT  3.720 -0.115 3.840 0.140 ;
        RECT  2.380 -0.115 3.720 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.845 4.400 1.375 ;
        RECT  3.820 1.145 4.280 1.375 ;
        RECT  3.700 1.135 3.820 1.375 ;
        RECT  3.460 1.145 3.700 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.640 ;
        RECT  4.355 0.210 4.425 0.640 ;
        RECT  3.450 0.210 4.355 0.280 ;
        RECT  4.010 0.545 4.130 0.615 ;
        RECT  3.940 0.350 4.010 1.045 ;
        RECT  3.600 0.975 3.940 1.045 ;
        RECT  3.800 0.520 3.870 0.905 ;
        RECT  3.085 0.835 3.800 0.905 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.905 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFSND0BWP

MACRO SDFSND1BWP
    CLASS CORE ;
    FOREIGN SDFSND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.185 4.585 1.045 ;
        RECT  4.495 0.185 4.515 0.465 ;
        RECT  4.495 0.730 4.515 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.210 0.350 4.280 0.775 ;
        RECT  4.095 0.350 4.210 0.470 ;
        RECT  4.185 0.695 4.210 0.775 ;
        RECT  4.095 0.695 4.185 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.280 -0.115 4.400 0.140 ;
        RECT  3.840 -0.115 4.280 0.115 ;
        RECT  3.720 -0.115 3.840 0.140 ;
        RECT  2.380 -0.115 3.720 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.375 1.145 4.620 1.375 ;
        RECT  4.305 0.895 4.375 1.375 ;
        RECT  3.820 1.145 4.305 1.375 ;
        RECT  3.700 1.135 3.820 1.375 ;
        RECT  3.460 1.145 3.700 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.520 4.445 0.640 ;
        RECT  4.355 0.210 4.425 0.640 ;
        RECT  3.450 0.210 4.355 0.280 ;
        RECT  4.010 0.545 4.130 0.615 ;
        RECT  3.940 0.350 4.010 1.045 ;
        RECT  3.600 0.975 3.940 1.045 ;
        RECT  3.800 0.520 3.870 0.905 ;
        RECT  3.085 0.835 3.800 0.905 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.905 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSND1BWP

MACRO SDFSND2BWP
    CLASS CORE ;
    FOREIGN SDFSND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.805 0.355 4.865 0.815 ;
        RECT  4.795 0.185 4.805 1.035 ;
        RECT  4.735 0.185 4.795 0.465 ;
        RECT  4.735 0.745 4.795 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.350 4.445 1.045 ;
        RECT  4.360 0.350 4.375 0.480 ;
        RECT  4.355 0.745 4.375 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.300 ;
        RECT  4.640 -0.115 4.910 0.115 ;
        RECT  4.520 -0.115 4.640 0.140 ;
        RECT  4.250 -0.115 4.520 0.115 ;
        RECT  4.130 -0.115 4.250 0.140 ;
        RECT  3.850 -0.115 4.130 0.115 ;
        RECT  3.730 -0.115 3.850 0.140 ;
        RECT  2.380 -0.115 3.730 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.905 4.990 1.375 ;
        RECT  4.615 1.145 4.910 1.375 ;
        RECT  4.545 0.735 4.615 1.375 ;
        RECT  4.250 1.145 4.545 1.375 ;
        RECT  4.130 1.120 4.250 1.375 ;
        RECT  3.865 1.145 4.130 1.375 ;
        RECT  3.795 0.980 3.865 1.375 ;
        RECT  3.460 1.145 3.795 1.375 ;
        RECT  3.340 1.015 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.630 0.545 4.720 0.615 ;
        RECT  4.560 0.210 4.630 0.615 ;
        RECT  3.450 0.210 4.560 0.280 ;
        RECT  4.230 0.520 4.300 0.640 ;
        RECT  4.160 0.365 4.230 1.050 ;
        RECT  3.765 0.365 4.160 0.435 ;
        RECT  3.950 0.980 4.160 1.050 ;
        RECT  3.905 0.520 3.975 0.910 ;
        RECT  3.085 0.840 3.905 0.910 ;
        RECT  3.695 0.365 3.765 0.640 ;
        RECT  3.230 0.695 3.650 0.765 ;
        RECT  3.380 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.380 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.160 0.355 3.230 0.765 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.910 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSND2BWP

MACRO SDFSND4BWP
    CLASS CORE ;
    FOREIGN SDFSND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.640 ;
        RECT  3.470 0.520 3.535 0.640 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.185 5.505 0.465 ;
        RECT  5.495 0.765 5.505 1.065 ;
        RECT  5.435 0.185 5.495 1.065 ;
        RECT  5.285 0.355 5.435 0.905 ;
        RECT  5.145 0.355 5.285 0.465 ;
        RECT  5.145 0.765 5.285 0.905 ;
        RECT  5.075 0.185 5.145 0.465 ;
        RECT  5.075 0.765 5.145 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.355 4.790 0.455 ;
        RECT  4.695 0.765 4.765 1.065 ;
        RECT  4.655 0.765 4.695 0.905 ;
        RECT  4.445 0.355 4.655 0.905 ;
        RECT  4.290 0.355 4.445 0.455 ;
        RECT  4.385 0.765 4.445 0.905 ;
        RECT  4.315 0.765 4.385 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.465 ;
        RECT  5.350 -0.115 5.610 0.115 ;
        RECT  5.230 -0.115 5.350 0.275 ;
        RECT  4.980 -0.115 5.230 0.115 ;
        RECT  4.860 -0.115 4.980 0.140 ;
        RECT  4.600 -0.115 4.860 0.115 ;
        RECT  4.480 -0.115 4.600 0.140 ;
        RECT  4.220 -0.115 4.480 0.115 ;
        RECT  4.100 -0.115 4.220 0.140 ;
        RECT  3.840 -0.115 4.100 0.115 ;
        RECT  3.720 -0.115 3.840 0.140 ;
        RECT  2.380 -0.115 3.720 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.480 -0.115 2.260 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.685 5.690 1.375 ;
        RECT  5.325 1.145 5.610 1.375 ;
        RECT  5.255 0.975 5.325 1.375 ;
        RECT  4.945 1.145 5.255 1.375 ;
        RECT  4.875 0.745 4.945 1.375 ;
        RECT  4.590 1.145 4.875 1.375 ;
        RECT  4.490 0.985 4.590 1.375 ;
        RECT  4.220 1.145 4.490 1.375 ;
        RECT  4.100 1.110 4.220 1.375 ;
        RECT  3.850 1.145 4.100 1.375 ;
        RECT  3.730 1.005 3.850 1.375 ;
        RECT  3.490 1.145 3.730 1.375 ;
        RECT  3.370 1.005 3.490 1.375 ;
        RECT  2.730 1.145 3.370 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.440 1.145 2.250 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.145 0.355 5.215 0.465 ;
        RECT  5.145 0.765 5.215 0.905 ;
        RECT  5.075 0.185 5.145 0.465 ;
        RECT  5.075 0.765 5.145 1.065 ;
        RECT  4.725 0.355 4.790 0.455 ;
        RECT  4.725 0.765 4.765 1.065 ;
        RECT  4.290 0.355 4.375 0.455 ;
        RECT  4.315 0.765 4.375 1.065 ;
        RECT  4.950 0.545 5.110 0.615 ;
        RECT  4.880 0.210 4.950 0.615 ;
        RECT  3.450 0.210 4.880 0.280 ;
        RECT  4.200 0.545 4.325 0.615 ;
        RECT  4.130 0.365 4.200 0.990 ;
        RECT  3.755 0.365 4.130 0.435 ;
        RECT  3.920 0.890 4.130 0.990 ;
        RECT  3.935 0.520 4.005 0.810 ;
        RECT  3.820 0.740 3.935 0.810 ;
        RECT  3.750 0.740 3.820 0.935 ;
        RECT  3.685 0.365 3.755 0.640 ;
        RECT  3.085 0.865 3.750 0.935 ;
        RECT  3.230 0.720 3.670 0.790 ;
        RECT  3.330 0.210 3.450 0.425 ;
        RECT  3.230 0.355 3.330 0.425 ;
        RECT  2.040 0.205 3.260 0.275 ;
        RECT  3.160 0.355 3.230 0.790 ;
        RECT  3.030 0.385 3.160 0.455 ;
        RECT  3.015 0.560 3.085 0.935 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.665 0.350 1.735 0.795 ;
        RECT  1.540 0.350 1.665 0.420 ;
        RECT  1.510 0.725 1.665 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSND4BWP

MACRO SDFSNQD0BWP
    CLASS CORE ;
    FOREIGN SDFSNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0112 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.490 0.500 3.535 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.185 4.445 0.905 ;
        RECT  4.355 0.185 4.375 0.305 ;
        RECT  4.355 0.755 4.375 0.905 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.355 0.810 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 -0.115 4.480 0.115 ;
        RECT  4.175 -0.115 4.245 0.315 ;
        RECT  3.870 -0.115 4.175 0.115 ;
        RECT  3.750 -0.115 3.870 0.280 ;
        RECT  2.380 -0.115 3.750 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.285 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 1.145 4.480 1.375 ;
        RECT  4.175 0.755 4.245 1.375 ;
        RECT  3.870 1.145 4.175 1.375 ;
        RECT  3.750 1.020 3.870 1.375 ;
        RECT  3.460 1.145 3.750 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.545 4.270 0.615 ;
        RECT  4.000 0.350 4.070 0.895 ;
        RECT  3.745 0.350 4.000 0.420 ;
        RECT  3.980 0.755 4.000 0.895 ;
        RECT  3.910 0.520 3.930 0.640 ;
        RECT  3.840 0.520 3.910 0.950 ;
        RECT  3.085 0.880 3.840 0.950 ;
        RECT  3.675 0.350 3.745 0.640 ;
        RECT  3.265 0.740 3.650 0.810 ;
        RECT  3.265 0.355 3.460 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.195 0.355 3.265 0.810 ;
        RECT  3.030 0.385 3.195 0.455 ;
        RECT  3.015 0.560 3.085 0.950 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.740 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.920 0.500 1.000 0.770 ;
        RECT  0.585 0.700 0.920 0.770 ;
        RECT  0.620 0.195 0.740 0.280 ;
        RECT  0.615 0.840 0.685 1.055 ;
        RECT  0.535 0.630 0.585 0.770 ;
        RECT  0.465 0.355 0.535 0.915 ;
        RECT  0.125 0.355 0.465 0.425 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.845 0.125 1.060 ;
    END
END SDFSNQD0BWP

MACRO SDFSNQD1BWP
    CLASS CORE ;
    FOREIGN SDFSNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0404 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.355 0.195 4.445 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 -0.115 4.480 0.115 ;
        RECT  4.175 -0.115 4.245 0.475 ;
        RECT  3.890 -0.115 4.175 0.115 ;
        RECT  3.770 -0.115 3.890 0.285 ;
        RECT  2.380 -0.115 3.770 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 1.145 4.480 1.375 ;
        RECT  4.175 0.735 4.245 1.375 ;
        RECT  3.890 1.145 4.175 1.375 ;
        RECT  3.770 1.020 3.890 1.375 ;
        RECT  3.460 1.145 3.770 1.375 ;
        RECT  3.340 1.020 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.070 0.545 4.270 0.615 ;
        RECT  4.045 0.370 4.070 1.035 ;
        RECT  4.000 0.185 4.045 1.035 ;
        RECT  3.975 0.185 4.000 0.440 ;
        RECT  3.980 0.735 4.000 1.035 ;
        RECT  3.745 0.370 3.975 0.440 ;
        RECT  3.910 0.520 3.930 0.640 ;
        RECT  3.840 0.520 3.910 0.950 ;
        RECT  3.085 0.880 3.840 0.950 ;
        RECT  3.675 0.370 3.745 0.640 ;
        RECT  3.265 0.740 3.650 0.810 ;
        RECT  3.265 0.355 3.460 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.195 0.355 3.265 0.810 ;
        RECT  3.030 0.385 3.195 0.455 ;
        RECT  3.015 0.560 3.085 0.950 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSNQD1BWP

MACRO SDFSNQD2BWP
    CLASS CORE ;
    FOREIGN SDFSNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  3.470 0.510 3.535 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.385 0.355 4.445 0.815 ;
        RECT  4.375 0.185 4.385 1.035 ;
        RECT  4.315 0.185 4.375 0.465 ;
        RECT  4.315 0.745 4.375 1.035 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.300 ;
        RECT  4.195 -0.115 4.490 0.115 ;
        RECT  4.125 -0.115 4.195 0.300 ;
        RECT  3.850 -0.115 4.125 0.115 ;
        RECT  3.730 -0.115 3.850 0.280 ;
        RECT  2.380 -0.115 3.730 0.115 ;
        RECT  2.260 -0.115 2.380 0.130 ;
        RECT  1.440 -0.115 2.260 0.115 ;
        RECT  1.320 -0.115 1.440 0.125 ;
        RECT  1.140 -0.115 1.320 0.115 ;
        RECT  1.020 -0.115 1.140 0.125 ;
        RECT  0.330 -0.115 1.020 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.490 0.905 4.570 1.375 ;
        RECT  4.220 1.145 4.490 1.375 ;
        RECT  4.100 1.005 4.220 1.375 ;
        RECT  3.850 1.145 4.100 1.375 ;
        RECT  3.730 1.005 3.850 1.375 ;
        RECT  3.460 1.145 3.730 1.375 ;
        RECT  3.340 1.015 3.460 1.375 ;
        RECT  2.730 1.145 3.340 1.375 ;
        RECT  2.610 0.990 2.730 1.375 ;
        RECT  2.370 1.145 2.610 1.375 ;
        RECT  2.250 1.005 2.370 1.375 ;
        RECT  1.400 1.145 2.250 1.375 ;
        RECT  1.280 1.130 1.400 1.375 ;
        RECT  1.100 1.145 1.280 1.375 ;
        RECT  0.980 1.130 1.100 1.375 ;
        RECT  0.330 1.145 0.980 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.180 0.520 4.270 0.640 ;
        RECT  4.110 0.370 4.180 0.935 ;
        RECT  4.005 0.370 4.110 0.440 ;
        RECT  3.900 0.865 4.110 0.935 ;
        RECT  3.935 0.185 4.005 0.440 ;
        RECT  3.745 0.370 3.935 0.440 ;
        RECT  3.865 0.520 3.935 0.790 ;
        RECT  3.810 0.720 3.865 0.790 ;
        RECT  3.740 0.720 3.810 0.935 ;
        RECT  3.675 0.370 3.745 0.640 ;
        RECT  3.085 0.865 3.740 0.935 ;
        RECT  3.265 0.720 3.650 0.790 ;
        RECT  3.265 0.355 3.450 0.425 ;
        RECT  2.020 0.205 3.270 0.275 ;
        RECT  3.195 0.355 3.265 0.790 ;
        RECT  3.030 0.385 3.195 0.455 ;
        RECT  3.015 0.560 3.085 0.935 ;
        RECT  2.925 0.560 3.015 0.630 ;
        RECT  2.745 0.710 2.930 0.780 ;
        RECT  2.855 0.360 2.925 0.630 ;
        RECT  2.815 0.850 2.885 1.060 ;
        RECT  2.145 0.850 2.815 0.920 ;
        RECT  2.675 0.360 2.745 0.780 ;
        RECT  2.140 0.710 2.675 0.780 ;
        RECT  2.385 0.375 2.455 0.640 ;
        RECT  1.965 0.375 2.385 0.445 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.195 1.840 0.265 ;
        RECT  1.720 0.740 1.790 1.055 ;
        RECT  1.650 0.575 1.730 0.645 ;
        RECT  0.685 0.985 1.720 1.055 ;
        RECT  1.580 0.350 1.650 0.795 ;
        RECT  1.520 0.350 1.580 0.420 ;
        RECT  1.490 0.725 1.580 0.795 ;
        RECT  1.410 0.520 1.510 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.350 0.935 0.420 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.350 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSNQD2BWP

MACRO SDFSNQD4BWP
    CLASS CORE ;
    FOREIGN SDFSNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0308 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.0432 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.640 ;
        RECT  3.470 0.520 3.535 0.640 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.805 0.465 ;
        RECT  4.795 0.765 4.805 1.065 ;
        RECT  4.735 0.185 4.795 1.065 ;
        RECT  4.585 0.355 4.735 0.905 ;
        RECT  4.445 0.355 4.585 0.465 ;
        RECT  4.445 0.765 4.585 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.765 4.445 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.905 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.465 ;
        RECT  4.650 -0.115 4.910 0.115 ;
        RECT  4.530 -0.115 4.650 0.275 ;
        RECT  4.260 -0.115 4.530 0.115 ;
        RECT  4.140 -0.115 4.260 0.280 ;
        RECT  3.870 -0.115 4.140 0.115 ;
        RECT  3.750 -0.115 3.870 0.280 ;
        RECT  2.400 -0.115 3.750 0.115 ;
        RECT  2.280 -0.115 2.400 0.130 ;
        RECT  1.480 -0.115 2.280 0.115 ;
        RECT  1.360 -0.115 1.480 0.130 ;
        RECT  1.120 -0.115 1.360 0.115 ;
        RECT  1.000 -0.115 1.120 0.130 ;
        RECT  0.330 -0.115 1.000 0.115 ;
        RECT  0.210 -0.115 0.330 0.280 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.685 4.990 1.375 ;
        RECT  4.625 1.145 4.910 1.375 ;
        RECT  4.555 0.975 4.625 1.375 ;
        RECT  4.260 1.145 4.555 1.375 ;
        RECT  4.140 1.005 4.260 1.375 ;
        RECT  3.870 1.145 4.140 1.375 ;
        RECT  3.750 1.005 3.870 1.375 ;
        RECT  3.480 1.145 3.750 1.375 ;
        RECT  3.360 1.015 3.480 1.375 ;
        RECT  2.750 1.145 3.360 1.375 ;
        RECT  2.630 0.990 2.750 1.375 ;
        RECT  2.390 1.145 2.630 1.375 ;
        RECT  2.270 0.990 2.390 1.375 ;
        RECT  1.440 1.145 2.270 1.375 ;
        RECT  1.320 1.125 1.440 1.375 ;
        RECT  1.080 1.145 1.320 1.375 ;
        RECT  0.960 1.125 1.080 1.375 ;
        RECT  0.330 1.145 0.960 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.355 4.515 0.465 ;
        RECT  4.445 0.765 4.515 0.905 ;
        RECT  4.375 0.185 4.445 0.465 ;
        RECT  4.375 0.765 4.445 1.065 ;
        RECT  4.200 0.545 4.410 0.615 ;
        RECT  4.130 0.370 4.200 0.935 ;
        RECT  4.025 0.370 4.130 0.440 ;
        RECT  3.920 0.865 4.130 0.935 ;
        RECT  3.955 0.185 4.025 0.440 ;
        RECT  3.955 0.520 4.025 0.790 ;
        RECT  3.765 0.370 3.955 0.440 ;
        RECT  3.830 0.720 3.955 0.790 ;
        RECT  3.760 0.720 3.830 0.935 ;
        RECT  3.695 0.370 3.765 0.640 ;
        RECT  3.105 0.865 3.760 0.935 ;
        RECT  3.285 0.720 3.670 0.790 ;
        RECT  3.285 0.355 3.465 0.425 ;
        RECT  2.040 0.205 3.290 0.275 ;
        RECT  3.215 0.355 3.285 0.790 ;
        RECT  3.050 0.385 3.215 0.455 ;
        RECT  3.035 0.560 3.105 0.935 ;
        RECT  2.945 0.560 3.035 0.630 ;
        RECT  2.765 0.710 2.950 0.780 ;
        RECT  2.875 0.360 2.945 0.630 ;
        RECT  2.835 0.850 2.905 1.060 ;
        RECT  2.145 0.850 2.835 0.920 ;
        RECT  2.695 0.360 2.765 0.780 ;
        RECT  2.295 0.710 2.695 0.780 ;
        RECT  2.405 0.375 2.475 0.640 ;
        RECT  1.965 0.375 2.405 0.445 ;
        RECT  2.225 0.520 2.295 0.780 ;
        RECT  2.075 0.850 2.145 1.075 ;
        RECT  1.970 1.005 2.075 1.075 ;
        RECT  1.895 0.375 1.965 0.930 ;
        RECT  0.610 0.205 1.860 0.275 ;
        RECT  1.630 0.875 1.810 0.945 ;
        RECT  1.665 0.350 1.735 0.795 ;
        RECT  1.540 0.350 1.665 0.420 ;
        RECT  1.510 0.725 1.665 0.795 ;
        RECT  1.560 0.875 1.630 1.055 ;
        RECT  0.685 0.985 1.560 1.055 ;
        RECT  1.410 0.520 1.535 0.640 ;
        RECT  1.340 0.345 1.410 0.915 ;
        RECT  1.170 0.345 1.340 0.415 ;
        RECT  1.120 0.845 1.340 0.915 ;
        RECT  0.830 0.355 0.935 0.425 ;
        RECT  0.830 0.845 0.900 0.915 ;
        RECT  0.760 0.355 0.830 0.915 ;
        RECT  0.615 0.795 0.685 1.055 ;
        RECT  0.535 0.530 0.585 0.650 ;
        RECT  0.465 0.350 0.535 0.915 ;
        RECT  0.125 0.350 0.465 0.420 ;
        RECT  0.125 0.845 0.465 0.915 ;
        RECT  0.055 0.200 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFSNQD4BWP

MACRO SDFXD0BWP
    CLASS CORE ;
    FOREIGN SDFXD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.355 0.345 5.425 0.905 ;
        RECT  5.335 0.345 5.355 0.465 ;
        RECT  5.335 0.735 5.355 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.210 5.145 0.485 ;
        RECT  5.030 0.370 5.075 0.485 ;
        RECT  4.960 0.370 5.030 0.790 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.365 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 -0.115 5.460 0.115 ;
        RECT  5.120 -0.115 5.240 0.140 ;
        RECT  4.665 -0.115 5.120 0.115 ;
        RECT  4.595 -0.115 4.665 0.310 ;
        RECT  3.940 -0.115 4.595 0.115 ;
        RECT  3.840 -0.115 3.940 0.420 ;
        RECT  3.555 -0.115 3.840 0.115 ;
        RECT  3.485 -0.115 3.555 0.250 ;
        RECT  2.520 -0.115 3.485 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.215 1.145 5.460 1.375 ;
        RECT  5.145 1.010 5.215 1.375 ;
        RECT  4.670 1.145 5.145 1.375 ;
        RECT  4.600 0.950 4.670 1.375 ;
        RECT  3.900 1.145 4.600 1.375 ;
        RECT  3.780 1.040 3.900 1.375 ;
        RECT  3.550 1.145 3.780 1.375 ;
        RECT  3.430 0.980 3.550 1.375 ;
        RECT  2.520 1.145 3.430 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.265 0.515 5.285 0.670 ;
        RECT  5.215 0.515 5.265 0.940 ;
        RECT  5.195 0.600 5.215 0.940 ;
        RECT  4.890 0.870 5.195 0.940 ;
        RECT  4.845 0.385 4.890 0.940 ;
        RECT  4.820 0.190 4.845 1.070 ;
        RECT  4.775 0.190 4.820 0.455 ;
        RECT  4.775 0.870 4.820 1.070 ;
        RECT  4.460 0.385 4.775 0.455 ;
        RECT  4.650 0.530 4.750 0.630 ;
        RECT  4.530 0.560 4.650 0.630 ;
        RECT  4.460 0.560 4.530 1.065 ;
        RECT  4.390 0.560 4.460 0.630 ;
        RECT  4.210 0.995 4.460 1.065 ;
        RECT  4.320 0.315 4.390 0.630 ;
        RECT  4.250 0.790 4.385 0.910 ;
        RECT  4.190 0.315 4.320 0.385 ;
        RECT  4.180 0.490 4.250 0.910 ;
        RECT  3.745 0.490 4.180 0.560 ;
        RECT  3.300 0.840 4.180 0.910 ;
        RECT  3.475 0.630 4.010 0.700 ;
        RECT  3.675 0.320 3.745 0.560 ;
        RECT  3.405 0.345 3.475 0.700 ;
        RECT  3.300 0.345 3.405 0.415 ;
        RECT  3.230 0.195 3.300 0.415 ;
        RECT  3.230 0.500 3.300 0.910 ;
        RECT  3.020 0.195 3.230 0.265 ;
        RECT  3.140 1.005 3.205 1.075 ;
        RECT  3.090 0.350 3.160 0.615 ;
        RECT  3.070 0.850 3.140 1.075 ;
        RECT  3.080 0.545 3.090 0.615 ;
        RECT  2.980 0.545 3.080 0.780 ;
        RECT  2.505 0.850 3.070 0.920 ;
        RECT  2.950 0.195 3.020 0.465 ;
        RECT  2.720 0.545 2.980 0.615 ;
        RECT  2.645 0.395 2.950 0.465 ;
        RECT  2.120 0.990 2.920 1.060 ;
        RECT  2.790 0.200 2.880 0.320 ;
        RECT  0.370 0.200 2.790 0.270 ;
        RECT  2.645 0.710 2.710 0.780 ;
        RECT  2.575 0.395 2.645 0.780 ;
        RECT  2.435 0.350 2.505 0.920 ;
        RECT  2.205 0.350 2.435 0.420 ;
        RECT  2.205 0.850 2.435 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.365 0.700 0.925 ;
        RECT  0.570 0.365 0.630 0.435 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXD0BWP

MACRO SDFXD1BWP
    CLASS CORE ;
    FOREIGN SDFXD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.355 0.185 5.425 1.045 ;
        RECT  5.335 0.185 5.355 0.465 ;
        RECT  5.335 0.735 5.355 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.030 0.210 5.145 0.485 ;
        RECT  4.960 0.210 5.030 0.790 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 -0.115 5.460 0.115 ;
        RECT  5.120 -0.115 5.240 0.140 ;
        RECT  4.665 -0.115 5.120 0.115 ;
        RECT  4.595 -0.115 4.665 0.310 ;
        RECT  3.950 -0.115 4.595 0.115 ;
        RECT  3.830 -0.115 3.950 0.400 ;
        RECT  3.555 -0.115 3.830 0.115 ;
        RECT  3.485 -0.115 3.555 0.250 ;
        RECT  2.520 -0.115 3.485 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 1.145 5.460 1.375 ;
        RECT  5.120 1.010 5.240 1.375 ;
        RECT  4.670 1.145 5.120 1.375 ;
        RECT  4.600 0.950 4.670 1.375 ;
        RECT  3.875 1.145 4.600 1.375 ;
        RECT  3.805 1.010 3.875 1.375 ;
        RECT  3.550 1.145 3.805 1.375 ;
        RECT  3.430 0.980 3.550 1.375 ;
        RECT  2.520 1.145 3.430 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.265 0.515 5.285 0.670 ;
        RECT  5.215 0.515 5.265 0.940 ;
        RECT  5.195 0.600 5.215 0.940 ;
        RECT  4.890 0.870 5.195 0.940 ;
        RECT  4.845 0.385 4.890 0.940 ;
        RECT  4.820 0.190 4.845 1.070 ;
        RECT  4.775 0.190 4.820 0.455 ;
        RECT  4.775 0.870 4.820 1.070 ;
        RECT  4.460 0.385 4.775 0.455 ;
        RECT  4.650 0.530 4.750 0.630 ;
        RECT  4.530 0.560 4.650 0.630 ;
        RECT  4.460 0.560 4.530 1.065 ;
        RECT  4.390 0.560 4.460 0.630 ;
        RECT  4.210 0.995 4.460 1.065 ;
        RECT  4.320 0.315 4.390 0.630 ;
        RECT  4.250 0.790 4.385 0.910 ;
        RECT  4.190 0.315 4.320 0.385 ;
        RECT  4.180 0.490 4.250 0.910 ;
        RECT  3.745 0.490 4.180 0.560 ;
        RECT  3.300 0.840 4.180 0.910 ;
        RECT  3.475 0.630 4.010 0.700 ;
        RECT  3.675 0.290 3.745 0.560 ;
        RECT  3.405 0.345 3.475 0.700 ;
        RECT  3.300 0.345 3.405 0.415 ;
        RECT  3.230 0.195 3.300 0.415 ;
        RECT  3.230 0.500 3.300 0.910 ;
        RECT  3.020 0.195 3.230 0.265 ;
        RECT  3.140 1.005 3.205 1.075 ;
        RECT  3.090 0.350 3.160 0.615 ;
        RECT  3.070 0.850 3.140 1.075 ;
        RECT  3.080 0.545 3.090 0.615 ;
        RECT  2.980 0.545 3.080 0.780 ;
        RECT  2.505 0.850 3.070 0.920 ;
        RECT  2.950 0.195 3.020 0.460 ;
        RECT  2.720 0.545 2.980 0.615 ;
        RECT  2.645 0.390 2.950 0.460 ;
        RECT  2.120 0.990 2.920 1.060 ;
        RECT  2.790 0.200 2.880 0.320 ;
        RECT  0.370 0.200 2.790 0.270 ;
        RECT  2.645 0.710 2.710 0.780 ;
        RECT  2.575 0.390 2.645 0.780 ;
        RECT  2.435 0.350 2.505 0.920 ;
        RECT  2.205 0.350 2.435 0.420 ;
        RECT  2.205 0.850 2.435 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXD1BWP

MACRO SDFXD2BWP
    CLASS CORE ;
    FOREIGN SDFXD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.505 0.355 5.565 0.805 ;
        RECT  5.495 0.185 5.505 1.035 ;
        RECT  5.435 0.185 5.495 0.465 ;
        RECT  5.435 0.735 5.495 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.075 0.215 5.145 0.800 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.360 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.300 ;
        RECT  5.325 -0.115 5.610 0.115 ;
        RECT  5.255 -0.115 5.325 0.465 ;
        RECT  4.965 -0.115 5.255 0.115 ;
        RECT  4.895 -0.115 4.965 0.425 ;
        RECT  4.605 -0.115 4.895 0.115 ;
        RECT  4.535 -0.115 4.605 0.420 ;
        RECT  3.885 -0.115 4.535 0.115 ;
        RECT  3.815 -0.115 3.885 0.420 ;
        RECT  3.540 -0.115 3.815 0.115 ;
        RECT  3.420 -0.115 3.540 0.245 ;
        RECT  2.520 -0.115 3.420 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.905 5.690 1.375 ;
        RECT  5.350 1.145 5.610 1.375 ;
        RECT  5.230 1.010 5.350 1.375 ;
        RECT  4.990 1.145 5.230 1.375 ;
        RECT  4.870 1.010 4.990 1.375 ;
        RECT  4.610 1.145 4.870 1.375 ;
        RECT  4.540 0.950 4.610 1.375 ;
        RECT  3.825 1.145 4.540 1.375 ;
        RECT  3.755 0.980 3.825 1.375 ;
        RECT  3.445 1.145 3.755 1.375 ;
        RECT  3.375 0.980 3.445 1.375 ;
        RECT  2.520 1.145 3.375 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.350 0.545 5.420 0.615 ;
        RECT  5.280 0.545 5.350 0.940 ;
        RECT  4.850 0.870 5.280 0.940 ;
        RECT  4.785 0.490 4.850 0.940 ;
        RECT  4.780 0.300 4.785 1.070 ;
        RECT  4.715 0.300 4.780 0.560 ;
        RECT  4.715 0.870 4.780 1.070 ;
        RECT  4.400 0.490 4.715 0.560 ;
        RECT  4.470 0.635 4.700 0.705 ;
        RECT  4.400 0.635 4.470 1.045 ;
        RECT  4.320 0.635 4.400 0.705 ;
        RECT  4.130 0.975 4.400 1.045 ;
        RECT  4.180 0.785 4.325 0.905 ;
        RECT  4.250 0.315 4.320 0.705 ;
        RECT  4.140 0.315 4.250 0.385 ;
        RECT  4.110 0.490 4.180 0.905 ;
        RECT  3.705 0.490 4.110 0.560 ;
        RECT  3.645 0.835 4.110 0.905 ;
        RECT  3.635 0.185 3.705 0.560 ;
        RECT  3.575 0.835 3.645 1.070 ;
        RECT  3.260 0.835 3.575 0.905 ;
        RECT  3.375 0.315 3.445 0.670 ;
        RECT  3.280 0.315 3.375 0.385 ;
        RECT  3.210 0.195 3.280 0.385 ;
        RECT  3.190 0.500 3.260 0.905 ;
        RECT  2.980 0.195 3.210 0.265 ;
        RECT  3.100 1.005 3.185 1.075 ;
        RECT  3.060 0.350 3.120 0.630 ;
        RECT  3.030 0.850 3.100 1.075 ;
        RECT  3.050 0.350 3.060 0.780 ;
        RECT  2.960 0.560 3.050 0.780 ;
        RECT  2.500 0.850 3.030 0.920 ;
        RECT  2.910 0.195 2.980 0.460 ;
        RECT  2.810 0.560 2.960 0.630 ;
        RECT  2.640 0.390 2.910 0.460 ;
        RECT  2.120 0.990 2.900 1.060 ;
        RECT  2.750 0.200 2.840 0.320 ;
        RECT  2.710 0.530 2.810 0.630 ;
        RECT  0.370 0.200 2.750 0.270 ;
        RECT  2.640 0.710 2.690 0.780 ;
        RECT  2.570 0.390 2.640 0.780 ;
        RECT  2.430 0.345 2.500 0.920 ;
        RECT  2.205 0.345 2.430 0.415 ;
        RECT  2.205 0.850 2.430 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXD2BWP

MACRO SDFXD4BWP
    CLASS CORE ;
    FOREIGN SDFXD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.755 0.185 6.765 0.465 ;
        RECT  6.755 0.765 6.765 1.065 ;
        RECT  6.695 0.185 6.755 1.065 ;
        RECT  6.545 0.355 6.695 0.905 ;
        RECT  6.405 0.355 6.545 0.465 ;
        RECT  6.405 0.765 6.545 0.905 ;
        RECT  6.335 0.185 6.405 0.465 ;
        RECT  6.335 0.765 6.405 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.700 6.070 0.800 ;
        RECT  5.975 0.185 6.060 0.485 ;
        RECT  5.915 0.355 5.975 0.485 ;
        RECT  5.705 0.355 5.915 0.800 ;
        RECT  5.685 0.355 5.705 0.485 ;
        RECT  5.600 0.700 5.705 0.800 ;
        RECT  5.615 0.185 5.685 0.485 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 -0.115 7.000 0.115 ;
        RECT  6.870 -0.115 6.950 0.465 ;
        RECT  6.610 -0.115 6.870 0.115 ;
        RECT  6.490 -0.115 6.610 0.275 ;
        RECT  6.225 -0.115 6.490 0.115 ;
        RECT  6.155 -0.115 6.225 0.465 ;
        RECT  5.890 -0.115 6.155 0.115 ;
        RECT  5.770 -0.115 5.890 0.280 ;
        RECT  5.505 -0.115 5.770 0.115 ;
        RECT  5.435 -0.115 5.505 0.305 ;
        RECT  5.075 -0.115 5.435 0.115 ;
        RECT  5.005 -0.115 5.075 0.305 ;
        RECT  4.340 -0.115 5.005 0.115 ;
        RECT  4.220 -0.115 4.340 0.225 ;
        RECT  3.555 -0.115 4.220 0.115 ;
        RECT  3.485 -0.115 3.555 0.250 ;
        RECT  2.520 -0.115 3.485 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 1.145 7.000 1.375 ;
        RECT  6.870 0.685 6.950 1.375 ;
        RECT  6.585 1.145 6.870 1.375 ;
        RECT  6.515 0.975 6.585 1.375 ;
        RECT  6.250 1.145 6.515 1.375 ;
        RECT  6.130 1.010 6.250 1.375 ;
        RECT  5.890 1.145 6.130 1.375 ;
        RECT  5.770 1.010 5.890 1.375 ;
        RECT  5.530 1.145 5.770 1.375 ;
        RECT  5.410 1.010 5.530 1.375 ;
        RECT  5.085 1.145 5.410 1.375 ;
        RECT  5.015 0.735 5.085 1.375 ;
        RECT  4.320 1.145 5.015 1.375 ;
        RECT  4.200 1.040 4.320 1.375 ;
        RECT  3.525 1.145 4.200 1.375 ;
        RECT  3.455 0.930 3.525 1.375 ;
        RECT  2.520 1.145 3.455 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.405 0.355 6.475 0.465 ;
        RECT  6.405 0.765 6.475 0.905 ;
        RECT  6.335 0.185 6.405 0.465 ;
        RECT  6.335 0.765 6.405 1.065 ;
        RECT  5.985 0.700 6.070 0.800 ;
        RECT  5.985 0.185 6.060 0.485 ;
        RECT  5.615 0.185 5.635 0.485 ;
        RECT  5.600 0.700 5.635 0.800 ;
        RECT  6.220 0.545 6.380 0.615 ;
        RECT  6.150 0.545 6.220 0.940 ;
        RECT  5.530 0.870 6.150 0.940 ;
        RECT  5.460 0.395 5.530 0.940 ;
        RECT  5.265 0.395 5.460 0.465 ;
        RECT  5.265 0.870 5.460 0.940 ;
        RECT  4.930 0.545 5.390 0.615 ;
        RECT  5.195 0.185 5.265 0.465 ;
        RECT  5.195 0.735 5.265 1.035 ;
        RECT  4.860 0.395 5.195 0.465 ;
        RECT  4.860 0.545 4.930 1.065 ;
        RECT  4.790 0.545 4.860 0.615 ;
        RECT  4.475 0.995 4.860 1.065 ;
        RECT  4.720 0.315 4.790 0.615 ;
        RECT  4.710 0.760 4.780 0.920 ;
        RECT  3.850 0.315 4.720 0.385 ;
        RECT  4.650 0.760 4.710 0.830 ;
        RECT  4.580 0.480 4.650 0.830 ;
        RECT  3.745 0.480 4.580 0.550 ;
        RECT  3.705 0.760 4.580 0.830 ;
        RECT  4.405 0.900 4.475 1.065 ;
        RECT  3.475 0.620 4.420 0.690 ;
        RECT  4.100 0.900 4.405 0.970 ;
        RECT  4.030 0.900 4.100 1.045 ;
        RECT  3.810 0.975 4.030 1.045 ;
        RECT  3.675 0.290 3.745 0.550 ;
        RECT  3.635 0.760 3.705 1.050 ;
        RECT  3.300 0.760 3.635 0.830 ;
        RECT  3.405 0.345 3.475 0.690 ;
        RECT  3.300 0.345 3.405 0.415 ;
        RECT  3.230 0.195 3.300 0.415 ;
        RECT  3.230 0.500 3.300 0.830 ;
        RECT  3.020 0.195 3.230 0.265 ;
        RECT  3.140 1.005 3.205 1.075 ;
        RECT  3.090 0.350 3.160 0.615 ;
        RECT  3.070 0.850 3.140 1.075 ;
        RECT  3.080 0.545 3.090 0.615 ;
        RECT  2.980 0.545 3.080 0.780 ;
        RECT  2.505 0.850 3.070 0.920 ;
        RECT  2.950 0.195 3.020 0.460 ;
        RECT  2.720 0.545 2.980 0.615 ;
        RECT  2.645 0.390 2.950 0.460 ;
        RECT  2.120 0.990 2.920 1.060 ;
        RECT  2.790 0.200 2.880 0.320 ;
        RECT  0.370 0.200 2.790 0.270 ;
        RECT  2.645 0.710 2.710 0.780 ;
        RECT  2.575 0.390 2.645 0.780 ;
        RECT  2.435 0.350 2.505 0.920 ;
        RECT  2.205 0.350 2.435 0.420 ;
        RECT  2.205 0.850 2.435 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXD4BWP

MACRO SDFXQD0BWP
    CLASS CORE ;
    FOREIGN SDFXQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.345 0.765 ;
        RECT  2.225 0.495 2.275 0.640 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.185 0.640 1.295 0.765 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0262 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SA
    PIN Q
        ANTENNAGATEAREA 0.0096 ;
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.215 4.725 1.045 ;
        RECT  4.635 0.215 4.655 0.415 ;
        RECT  4.635 0.905 4.655 1.045 ;
        RECT  4.355 0.345 4.635 0.415 ;
        RECT  4.285 0.345 4.355 0.610 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0146 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.640 ;
        RECT  0.685 0.520 0.715 0.640 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0146 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.535 0.520 0.575 0.640 ;
        RECT  0.455 0.355 0.535 0.640 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.495 2.635 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.115 4.760 0.115 ;
        RECT  4.400 -0.115 4.520 0.275 ;
        RECT  3.685 -0.115 4.400 0.115 ;
        RECT  3.615 -0.115 3.685 0.430 ;
        RECT  2.740 -0.115 3.615 0.115 ;
        RECT  2.620 -0.115 2.740 0.125 ;
        RECT  2.240 -0.115 2.620 0.115 ;
        RECT  2.120 -0.115 2.240 0.125 ;
        RECT  1.425 -0.115 2.120 0.115 ;
        RECT  1.355 -0.115 1.425 0.260 ;
        RECT  1.080 -0.115 1.355 0.115 ;
        RECT  0.960 -0.115 1.080 0.145 ;
        RECT  0.340 -0.115 0.960 0.115 ;
        RECT  0.220 -0.115 0.340 0.185 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.145 4.760 1.375 ;
        RECT  4.455 0.915 4.525 1.375 ;
        RECT  3.700 1.145 4.455 1.375 ;
        RECT  3.580 0.880 3.700 1.375 ;
        RECT  2.740 1.145 3.580 1.375 ;
        RECT  2.620 1.130 2.740 1.375 ;
        RECT  2.240 1.145 2.620 1.375 ;
        RECT  2.120 1.135 2.240 1.375 ;
        RECT  1.465 1.145 2.120 1.375 ;
        RECT  1.340 1.135 1.465 1.375 ;
        RECT  1.100 1.145 1.340 1.375 ;
        RECT  0.980 1.135 1.100 1.375 ;
        RECT  0.380 1.145 0.980 1.375 ;
        RECT  0.305 0.985 0.380 1.375 ;
        RECT  0.210 0.985 0.305 1.055 ;
        RECT  0.000 1.145 0.305 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.510 0.510 4.585 0.750 ;
        RECT  4.360 0.680 4.510 0.750 ;
        RECT  4.290 0.680 4.360 1.065 ;
        RECT  4.185 0.680 4.290 0.750 ;
        RECT  3.940 0.995 4.290 1.065 ;
        RECT  4.115 0.215 4.185 0.750 ;
        RECT  4.020 0.830 4.180 0.900 ;
        RECT  3.970 0.215 4.115 0.285 ;
        RECT  3.950 0.420 4.020 0.900 ;
        RECT  3.865 0.220 3.880 0.800 ;
        RECT  3.810 0.220 3.865 1.050 ;
        RECT  3.795 0.730 3.810 1.050 ;
        RECT  3.555 0.730 3.795 0.800 ;
        RECT  3.670 0.510 3.740 0.640 ;
        RECT  3.295 0.510 3.670 0.580 ;
        RECT  3.485 0.680 3.555 0.800 ;
        RECT  3.285 0.300 3.295 0.580 ;
        RECT  3.215 0.300 3.285 0.960 ;
        RECT  1.825 0.195 3.140 0.265 ;
        RECT  3.035 0.840 3.105 1.060 ;
        RECT  1.830 0.990 3.035 1.060 ;
        RECT  2.925 0.340 2.995 0.765 ;
        RECT  2.855 0.340 2.925 0.460 ;
        RECT  2.855 0.695 2.925 0.920 ;
        RECT  2.775 0.520 2.810 0.640 ;
        RECT  2.705 0.355 2.775 0.920 ;
        RECT  2.470 0.355 2.705 0.425 ;
        RECT  2.470 0.850 2.705 0.920 ;
        RECT  2.115 0.355 2.390 0.425 ;
        RECT  2.115 0.850 2.390 0.920 ;
        RECT  2.045 0.355 2.115 0.920 ;
        RECT  1.835 0.510 1.905 0.770 ;
        RECT  1.515 0.510 1.835 0.580 ;
        RECT  1.760 0.850 1.830 1.060 ;
        RECT  1.755 0.195 1.825 0.430 ;
        RECT  1.685 0.670 1.755 0.750 ;
        RECT  1.615 0.670 1.685 1.065 ;
        RECT  1.110 0.995 1.615 1.065 ;
        RECT  1.445 0.340 1.515 0.915 ;
        RECT  1.250 0.340 1.445 0.410 ;
        RECT  1.190 0.845 1.445 0.915 ;
        RECT  1.180 0.220 1.250 0.410 ;
        RECT  1.040 0.215 1.110 1.065 ;
        RECT  0.590 0.215 1.040 0.285 ;
        RECT  0.580 0.865 1.040 0.935 ;
        RECT  0.900 0.370 0.970 0.795 ;
        RECT  0.385 0.725 0.900 0.795 ;
        RECT  0.315 0.265 0.385 0.915 ;
        RECT  0.125 0.265 0.315 0.340 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.055 0.200 0.125 0.340 ;
        RECT  0.055 0.845 0.125 1.030 ;
    END
END SDFXQD0BWP

MACRO SDFXQD1BWP
    CLASS CORE ;
    FOREIGN SDFXQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.195 0.195 5.285 1.070 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.085 -0.115 5.320 0.115 ;
        RECT  5.015 -0.115 5.085 0.475 ;
        RECT  4.695 -0.115 5.015 0.115 ;
        RECT  4.625 -0.115 4.695 0.310 ;
        RECT  3.950 -0.115 4.625 0.115 ;
        RECT  3.830 -0.115 3.950 0.420 ;
        RECT  3.555 -0.115 3.830 0.115 ;
        RECT  3.485 -0.115 3.555 0.250 ;
        RECT  2.520 -0.115 3.485 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.085 1.145 5.320 1.375 ;
        RECT  5.015 0.685 5.085 1.375 ;
        RECT  4.695 1.145 5.015 1.375 ;
        RECT  4.625 0.950 4.695 1.375 ;
        RECT  3.875 1.145 4.625 1.375 ;
        RECT  3.805 1.010 3.875 1.375 ;
        RECT  3.550 1.145 3.805 1.375 ;
        RECT  3.430 0.980 3.550 1.375 ;
        RECT  2.520 1.145 3.430 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.885 0.385 4.930 0.940 ;
        RECT  4.860 0.190 4.885 1.070 ;
        RECT  4.815 0.190 4.860 0.455 ;
        RECT  4.815 0.870 4.860 1.070 ;
        RECT  4.480 0.385 4.815 0.455 ;
        RECT  4.690 0.530 4.790 0.630 ;
        RECT  4.550 0.560 4.690 0.630 ;
        RECT  4.480 0.560 4.550 1.065 ;
        RECT  4.390 0.560 4.480 0.630 ;
        RECT  4.210 0.995 4.480 1.065 ;
        RECT  4.320 0.315 4.390 0.630 ;
        RECT  4.250 0.790 4.385 0.910 ;
        RECT  4.190 0.315 4.320 0.385 ;
        RECT  4.180 0.490 4.250 0.910 ;
        RECT  3.745 0.490 4.180 0.560 ;
        RECT  3.300 0.840 4.180 0.910 ;
        RECT  3.475 0.630 4.010 0.700 ;
        RECT  3.675 0.290 3.745 0.560 ;
        RECT  3.405 0.345 3.475 0.700 ;
        RECT  3.300 0.345 3.405 0.415 ;
        RECT  3.230 0.195 3.300 0.415 ;
        RECT  3.230 0.500 3.300 0.910 ;
        RECT  3.020 0.195 3.230 0.265 ;
        RECT  3.140 1.005 3.205 1.075 ;
        RECT  3.090 0.350 3.160 0.615 ;
        RECT  3.070 0.850 3.140 1.075 ;
        RECT  3.080 0.545 3.090 0.615 ;
        RECT  2.980 0.545 3.080 0.780 ;
        RECT  2.505 0.850 3.070 0.920 ;
        RECT  2.950 0.195 3.020 0.460 ;
        RECT  2.720 0.545 2.980 0.615 ;
        RECT  2.645 0.390 2.950 0.460 ;
        RECT  2.120 0.990 2.920 1.060 ;
        RECT  2.790 0.200 2.880 0.320 ;
        RECT  0.370 0.200 2.790 0.270 ;
        RECT  2.645 0.710 2.710 0.780 ;
        RECT  2.575 0.390 2.645 0.780 ;
        RECT  2.435 0.350 2.505 0.920 ;
        RECT  2.205 0.350 2.435 0.420 ;
        RECT  2.205 0.850 2.435 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXQD1BWP

MACRO SDFXQD2BWP
    CLASS CORE ;
    FOREIGN SDFXQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.225 0.355 5.285 0.805 ;
        RECT  5.215 0.185 5.225 1.035 ;
        RECT  5.155 0.185 5.215 0.465 ;
        RECT  5.155 0.735 5.215 1.035 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0142 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.360 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.410 -0.115 5.460 0.115 ;
        RECT  5.330 -0.115 5.410 0.300 ;
        RECT  5.045 -0.115 5.330 0.115 ;
        RECT  4.975 -0.115 5.045 0.465 ;
        RECT  4.665 -0.115 4.975 0.115 ;
        RECT  4.595 -0.115 4.665 0.420 ;
        RECT  3.905 -0.115 4.595 0.115 ;
        RECT  3.835 -0.115 3.905 0.420 ;
        RECT  3.560 -0.115 3.835 0.115 ;
        RECT  3.440 -0.115 3.560 0.245 ;
        RECT  2.520 -0.115 3.440 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.410 1.145 5.460 1.375 ;
        RECT  5.330 0.905 5.410 1.375 ;
        RECT  5.045 1.145 5.330 1.375 ;
        RECT  4.975 0.685 5.045 1.375 ;
        RECT  4.655 1.145 4.975 1.375 ;
        RECT  4.585 0.940 4.655 1.375 ;
        RECT  3.845 1.145 4.585 1.375 ;
        RECT  3.775 0.980 3.845 1.375 ;
        RECT  3.465 1.145 3.775 1.375 ;
        RECT  3.395 0.980 3.465 1.375 ;
        RECT  2.520 1.145 3.395 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.845 0.490 4.905 1.045 ;
        RECT  4.835 0.300 4.845 1.045 ;
        RECT  4.775 0.300 4.835 0.560 ;
        RECT  4.740 0.975 4.835 1.045 ;
        RECT  4.460 0.490 4.775 0.560 ;
        RECT  4.510 0.645 4.760 0.715 ;
        RECT  4.440 0.645 4.510 1.045 ;
        RECT  4.360 0.645 4.440 0.715 ;
        RECT  4.170 0.975 4.440 1.045 ;
        RECT  4.220 0.785 4.365 0.905 ;
        RECT  4.290 0.315 4.360 0.715 ;
        RECT  4.180 0.315 4.290 0.385 ;
        RECT  4.150 0.490 4.220 0.905 ;
        RECT  3.725 0.490 4.150 0.560 ;
        RECT  3.665 0.835 4.150 0.905 ;
        RECT  3.655 0.185 3.725 0.560 ;
        RECT  3.595 0.835 3.665 1.070 ;
        RECT  3.260 0.835 3.595 0.905 ;
        RECT  3.395 0.315 3.465 0.670 ;
        RECT  3.280 0.315 3.395 0.385 ;
        RECT  3.210 0.195 3.280 0.385 ;
        RECT  3.190 0.500 3.260 0.905 ;
        RECT  2.980 0.195 3.210 0.265 ;
        RECT  3.100 1.005 3.185 1.075 ;
        RECT  3.060 0.350 3.120 0.630 ;
        RECT  3.030 0.850 3.100 1.075 ;
        RECT  3.050 0.350 3.060 0.780 ;
        RECT  2.960 0.560 3.050 0.780 ;
        RECT  2.500 0.850 3.030 0.920 ;
        RECT  2.910 0.195 2.980 0.460 ;
        RECT  2.810 0.560 2.960 0.630 ;
        RECT  2.640 0.390 2.910 0.460 ;
        RECT  2.120 0.990 2.900 1.060 ;
        RECT  2.750 0.200 2.840 0.320 ;
        RECT  2.710 0.530 2.810 0.630 ;
        RECT  0.370 0.200 2.750 0.270 ;
        RECT  2.640 0.710 2.690 0.780 ;
        RECT  2.570 0.390 2.640 0.780 ;
        RECT  2.430 0.345 2.500 0.920 ;
        RECT  2.205 0.345 2.430 0.415 ;
        RECT  2.205 0.850 2.430 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXQD2BWP

MACRO SDFXQD4BWP
    CLASS CORE ;
    FOREIGN SDFXQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.495 2.205 0.765 ;
        RECT  2.015 0.495 2.115 0.640 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.185 6.065 0.465 ;
        RECT  6.055 0.765 6.065 1.065 ;
        RECT  5.995 0.185 6.055 1.065 ;
        RECT  5.845 0.355 5.995 0.905 ;
        RECT  5.705 0.355 5.845 0.465 ;
        RECT  5.705 0.765 5.845 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.765 5.705 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.630 1.785 0.770 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.0168 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.285 0.625 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.465 ;
        RECT  5.910 -0.115 6.170 0.115 ;
        RECT  5.790 -0.115 5.910 0.275 ;
        RECT  5.525 -0.115 5.790 0.115 ;
        RECT  5.455 -0.115 5.525 0.305 ;
        RECT  5.115 -0.115 5.455 0.115 ;
        RECT  5.045 -0.115 5.115 0.305 ;
        RECT  4.360 -0.115 5.045 0.115 ;
        RECT  4.240 -0.115 4.360 0.225 ;
        RECT  3.555 -0.115 4.240 0.115 ;
        RECT  3.485 -0.115 3.555 0.250 ;
        RECT  2.520 -0.115 3.485 0.115 ;
        RECT  2.400 -0.115 2.520 0.130 ;
        RECT  2.130 -0.115 2.400 0.115 ;
        RECT  2.010 -0.115 2.130 0.125 ;
        RECT  0.840 -0.115 2.010 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.685 6.250 1.375 ;
        RECT  5.885 1.145 6.170 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  5.525 1.145 5.815 1.375 ;
        RECT  5.455 0.905 5.525 1.375 ;
        RECT  5.125 1.145 5.455 1.375 ;
        RECT  5.055 0.735 5.125 1.375 ;
        RECT  4.340 1.145 5.055 1.375 ;
        RECT  4.220 1.040 4.340 1.375 ;
        RECT  3.525 1.145 4.220 1.375 ;
        RECT  3.455 0.930 3.525 1.375 ;
        RECT  2.520 1.145 3.455 1.375 ;
        RECT  2.400 1.130 2.520 1.375 ;
        RECT  2.130 1.145 2.400 1.375 ;
        RECT  2.010 1.135 2.130 1.375 ;
        RECT  0.125 1.145 2.010 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.355 5.775 0.465 ;
        RECT  5.705 0.765 5.775 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.765 5.705 1.065 ;
        RECT  5.480 0.395 5.550 0.805 ;
        RECT  5.305 0.395 5.480 0.465 ;
        RECT  5.305 0.735 5.480 0.805 ;
        RECT  4.970 0.545 5.410 0.615 ;
        RECT  5.235 0.185 5.305 0.465 ;
        RECT  5.235 0.735 5.305 1.035 ;
        RECT  4.900 0.395 5.235 0.465 ;
        RECT  4.900 0.545 4.970 1.065 ;
        RECT  4.830 0.545 4.900 0.615 ;
        RECT  4.515 0.995 4.900 1.065 ;
        RECT  4.760 0.315 4.830 0.615 ;
        RECT  4.750 0.760 4.820 0.920 ;
        RECT  3.850 0.315 4.760 0.385 ;
        RECT  4.690 0.760 4.750 0.830 ;
        RECT  4.620 0.480 4.690 0.830 ;
        RECT  3.745 0.480 4.620 0.550 ;
        RECT  3.705 0.760 4.620 0.830 ;
        RECT  4.445 0.900 4.515 1.065 ;
        RECT  4.100 0.900 4.445 0.970 ;
        RECT  3.475 0.620 4.440 0.690 ;
        RECT  4.030 0.900 4.100 1.045 ;
        RECT  3.810 0.975 4.030 1.045 ;
        RECT  3.675 0.290 3.745 0.550 ;
        RECT  3.635 0.760 3.705 1.050 ;
        RECT  3.300 0.760 3.635 0.830 ;
        RECT  3.405 0.345 3.475 0.690 ;
        RECT  3.300 0.345 3.405 0.415 ;
        RECT  3.230 0.195 3.300 0.415 ;
        RECT  3.230 0.500 3.300 0.830 ;
        RECT  3.020 0.195 3.230 0.265 ;
        RECT  3.140 1.005 3.205 1.075 ;
        RECT  3.090 0.350 3.160 0.615 ;
        RECT  3.070 0.850 3.140 1.075 ;
        RECT  3.080 0.545 3.090 0.615 ;
        RECT  2.980 0.545 3.080 0.780 ;
        RECT  2.505 0.850 3.070 0.920 ;
        RECT  2.950 0.195 3.020 0.460 ;
        RECT  2.720 0.545 2.980 0.615 ;
        RECT  2.645 0.390 2.950 0.460 ;
        RECT  2.120 0.990 2.920 1.060 ;
        RECT  2.790 0.200 2.880 0.320 ;
        RECT  0.370 0.200 2.790 0.270 ;
        RECT  2.645 0.710 2.710 0.780 ;
        RECT  2.575 0.390 2.645 0.780 ;
        RECT  2.435 0.350 2.505 0.920 ;
        RECT  2.205 0.350 2.435 0.420 ;
        RECT  2.205 0.850 2.435 0.920 ;
        RECT  2.050 0.990 2.120 1.065 ;
        RECT  1.530 0.995 2.050 1.065 ;
        RECT  1.875 0.350 1.945 0.925 ;
        RECT  1.485 0.480 1.875 0.550 ;
        RECT  0.930 0.340 1.790 0.410 ;
        RECT  1.170 0.840 1.790 0.910 ;
        RECT  1.460 0.990 1.530 1.065 ;
        RECT  1.415 0.480 1.485 0.765 ;
        RECT  1.285 0.990 1.460 1.060 ;
        RECT  1.030 0.695 1.415 0.765 ;
        RECT  1.225 0.990 1.285 1.065 ;
        RECT  0.485 0.995 1.225 1.065 ;
        RECT  1.110 0.840 1.170 0.925 ;
        RECT  0.930 0.855 1.110 0.925 ;
        RECT  0.700 0.515 0.940 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SDFXQD4BWP

MACRO SEDFCND0BWP
    CLASS CORE ;
    FOREIGN SEDFCND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.330 5.705 0.905 ;
        RECT  5.615 0.330 5.635 0.450 ;
        RECT  5.615 0.765 5.635 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.405 0.215 5.425 0.485 ;
        RECT  5.335 0.215 5.405 0.905 ;
        RECT  5.215 0.215 5.335 0.345 ;
        RECT  5.235 0.775 5.335 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0348 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0176 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.295 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.495 4.865 0.765 ;
        RECT  4.745 0.495 4.795 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 -0.115 5.740 0.115 ;
        RECT  5.400 -0.115 5.520 0.140 ;
        RECT  4.740 -0.115 5.400 0.115 ;
        RECT  4.620 -0.115 4.740 0.200 ;
        RECT  3.690 -0.115 4.620 0.115 ;
        RECT  3.620 -0.115 3.690 0.265 ;
        RECT  2.580 -0.115 3.620 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.145 5.740 1.375 ;
        RECT  5.400 1.120 5.520 1.375 ;
        RECT  5.150 1.145 5.400 1.375 ;
        RECT  5.030 1.120 5.150 1.375 ;
        RECT  4.740 1.145 5.030 1.375 ;
        RECT  4.620 1.120 4.740 1.375 ;
        RECT  3.785 1.145 4.620 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.545 0.515 5.565 0.710 ;
        RECT  5.495 0.515 5.545 1.050 ;
        RECT  5.475 0.640 5.495 1.050 ;
        RECT  4.500 0.980 5.475 1.050 ;
        RECT  5.145 0.545 5.250 0.615 ;
        RECT  5.075 0.185 5.145 0.910 ;
        RECT  5.040 0.185 5.075 0.285 ;
        RECT  4.640 0.840 5.075 0.910 ;
        RECT  4.935 0.355 5.005 0.640 ;
        RECT  4.850 0.355 4.935 0.425 ;
        RECT  4.780 0.270 4.850 0.425 ;
        RECT  4.200 0.270 4.780 0.340 ;
        RECT  4.570 0.640 4.640 0.910 ;
        RECT  4.500 0.410 4.570 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.935 0.980 4.430 1.050 ;
        RECT  4.225 0.630 4.295 0.910 ;
        RECT  4.200 0.630 4.225 0.700 ;
        RECT  4.130 0.270 4.200 0.700 ;
        RECT  4.080 0.375 4.130 0.445 ;
        RECT  3.990 0.780 4.110 0.850 ;
        RECT  3.830 0.200 4.060 0.270 ;
        RECT  3.920 0.350 3.990 0.850 ;
        RECT  3.865 0.920 3.935 1.050 ;
        RECT  3.915 0.350 3.920 0.560 ;
        RECT  3.320 0.490 3.915 0.560 ;
        RECT  3.550 0.920 3.865 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.760 0.200 3.830 0.420 ;
        RECT  3.380 0.350 3.760 0.420 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.310 0.195 3.380 0.420 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.880 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  2.030 0.685 2.060 0.785 ;
        RECT  1.965 0.480 2.030 0.785 ;
        RECT  1.960 0.340 1.965 0.785 ;
        RECT  1.895 0.340 1.960 0.550 ;
        RECT  1.495 0.480 1.895 0.550 ;
        RECT  1.810 0.635 1.880 0.925 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.570 0.635 1.810 0.705 ;
        RECT  1.670 0.790 1.740 0.925 ;
        RECT  0.930 0.855 1.670 0.925 ;
        RECT  1.425 0.480 1.495 0.765 ;
        RECT  1.030 0.695 1.425 0.765 ;
        RECT  0.700 0.515 0.940 0.615 ;
        RECT  0.630 0.365 0.700 0.925 ;
        RECT  0.570 0.365 0.630 0.435 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCND0BWP

MACRO SEDFCND1BWP
    CLASS CORE ;
    FOREIGN SEDFCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.185 5.705 1.065 ;
        RECT  5.615 0.185 5.635 0.465 ;
        RECT  5.615 0.765 5.635 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.405 0.215 5.425 0.485 ;
        RECT  5.335 0.215 5.405 0.905 ;
        RECT  5.235 0.215 5.335 0.475 ;
        RECT  5.235 0.775 5.335 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.495 4.865 0.770 ;
        RECT  4.745 0.495 4.795 0.640 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 -0.115 5.740 0.115 ;
        RECT  5.400 -0.115 5.520 0.140 ;
        RECT  4.740 -0.115 5.400 0.115 ;
        RECT  4.620 -0.115 4.740 0.200 ;
        RECT  3.690 -0.115 4.620 0.115 ;
        RECT  3.620 -0.115 3.690 0.265 ;
        RECT  2.580 -0.115 3.620 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.145 5.740 1.375 ;
        RECT  5.400 1.120 5.520 1.375 ;
        RECT  5.150 1.145 5.400 1.375 ;
        RECT  5.030 1.120 5.150 1.375 ;
        RECT  4.740 1.145 5.030 1.375 ;
        RECT  4.620 1.120 4.740 1.375 ;
        RECT  3.785 1.145 4.620 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.545 0.515 5.565 0.710 ;
        RECT  5.495 0.515 5.545 1.050 ;
        RECT  5.475 0.640 5.495 1.050 ;
        RECT  4.500 0.980 5.475 1.050 ;
        RECT  5.145 0.545 5.230 0.615 ;
        RECT  5.075 0.185 5.145 0.910 ;
        RECT  5.040 0.185 5.075 0.285 ;
        RECT  4.640 0.840 5.075 0.910 ;
        RECT  4.935 0.355 5.005 0.640 ;
        RECT  4.850 0.355 4.935 0.425 ;
        RECT  4.780 0.270 4.850 0.425 ;
        RECT  4.200 0.270 4.780 0.340 ;
        RECT  4.570 0.640 4.640 0.910 ;
        RECT  4.500 0.410 4.570 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.935 0.980 4.430 1.050 ;
        RECT  4.225 0.630 4.295 0.910 ;
        RECT  4.200 0.630 4.225 0.700 ;
        RECT  4.130 0.270 4.200 0.700 ;
        RECT  4.080 0.375 4.130 0.445 ;
        RECT  3.990 0.780 4.110 0.850 ;
        RECT  3.830 0.200 4.060 0.270 ;
        RECT  3.920 0.350 3.990 0.850 ;
        RECT  3.865 0.920 3.935 1.050 ;
        RECT  3.915 0.350 3.920 0.560 ;
        RECT  3.320 0.490 3.915 0.560 ;
        RECT  3.550 0.920 3.865 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.760 0.200 3.830 0.420 ;
        RECT  3.380 0.350 3.760 0.420 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.310 0.195 3.380 0.420 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.905 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCND1BWP

MACRO SEDFCND2BWP
    CLASS CORE ;
    FOREIGN SEDFCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.785 0.355 5.845 0.805 ;
        RECT  5.775 0.185 5.785 1.035 ;
        RECT  5.715 0.185 5.775 0.465 ;
        RECT  5.715 0.735 5.775 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.355 0.215 5.425 0.780 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.495 4.865 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 -0.115 6.020 0.115 ;
        RECT  5.890 -0.115 5.970 0.300 ;
        RECT  5.605 -0.115 5.890 0.115 ;
        RECT  5.535 -0.115 5.605 0.465 ;
        RECT  5.250 -0.115 5.535 0.115 ;
        RECT  5.130 -0.115 5.250 0.145 ;
        RECT  4.680 -0.115 5.130 0.115 ;
        RECT  4.560 -0.115 4.680 0.200 ;
        RECT  3.720 -0.115 4.560 0.115 ;
        RECT  3.600 -0.115 3.720 0.220 ;
        RECT  2.580 -0.115 3.600 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 1.145 6.020 1.375 ;
        RECT  5.890 0.905 5.970 1.375 ;
        RECT  5.630 1.145 5.890 1.375 ;
        RECT  5.510 1.005 5.630 1.375 ;
        RECT  5.090 1.145 5.510 1.375 ;
        RECT  4.970 1.005 5.090 1.375 ;
        RECT  4.730 1.145 4.970 1.375 ;
        RECT  4.610 1.005 4.730 1.375 ;
        RECT  3.785 1.145 4.610 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.615 0.545 5.700 0.615 ;
        RECT  5.545 0.545 5.615 0.935 ;
        RECT  4.440 0.865 5.545 0.935 ;
        RECT  5.205 0.215 5.275 0.795 ;
        RECT  4.950 0.215 5.205 0.285 ;
        RECT  4.600 0.725 5.205 0.795 ;
        RECT  4.935 0.355 5.005 0.640 ;
        RECT  4.865 0.355 4.935 0.425 ;
        RECT  4.795 0.270 4.865 0.425 ;
        RECT  4.145 0.270 4.795 0.340 ;
        RECT  4.530 0.670 4.600 0.795 ;
        RECT  4.440 0.410 4.530 0.480 ;
        RECT  4.370 0.410 4.440 1.050 ;
        RECT  4.240 0.460 4.370 0.560 ;
        RECT  3.955 0.980 4.370 1.050 ;
        RECT  4.190 0.630 4.290 0.910 ;
        RECT  4.145 0.630 4.190 0.700 ;
        RECT  4.075 0.270 4.145 0.700 ;
        RECT  3.980 0.780 4.110 0.850 ;
        RECT  3.900 0.205 4.005 0.275 ;
        RECT  3.910 0.435 3.980 0.850 ;
        RECT  3.885 0.920 3.955 1.050 ;
        RECT  3.440 0.435 3.910 0.505 ;
        RECT  3.830 0.205 3.900 0.365 ;
        RECT  3.550 0.920 3.885 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.380 0.295 3.830 0.365 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.320 0.435 3.440 0.560 ;
        RECT  3.310 0.195 3.380 0.365 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.905 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCND2BWP

MACRO SEDFCND4BWP
    CLASS CORE ;
    FOREIGN SEDFCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.755 0.185 6.765 0.465 ;
        RECT  6.755 0.765 6.765 1.065 ;
        RECT  6.695 0.185 6.755 1.065 ;
        RECT  6.545 0.355 6.695 0.905 ;
        RECT  6.405 0.355 6.545 0.465 ;
        RECT  6.405 0.765 6.545 0.905 ;
        RECT  6.335 0.185 6.405 0.465 ;
        RECT  6.335 0.765 6.405 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.705 6.060 0.805 ;
        RECT  5.975 0.185 6.045 0.465 ;
        RECT  5.915 0.355 5.975 0.465 ;
        RECT  5.705 0.355 5.915 0.805 ;
        RECT  5.685 0.355 5.705 0.465 ;
        RECT  5.600 0.705 5.705 0.805 ;
        RECT  5.615 0.185 5.685 0.465 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.515 0.630 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.495 5.375 0.640 ;
        RECT  5.215 0.495 5.285 0.770 ;
        RECT  4.865 0.700 5.215 0.770 ;
        RECT  4.785 0.495 4.865 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 -0.115 7.000 0.115 ;
        RECT  6.870 -0.115 6.950 0.465 ;
        RECT  6.610 -0.115 6.870 0.115 ;
        RECT  6.490 -0.115 6.610 0.275 ;
        RECT  6.225 -0.115 6.490 0.115 ;
        RECT  6.155 -0.115 6.225 0.465 ;
        RECT  5.890 -0.115 6.155 0.115 ;
        RECT  5.770 -0.115 5.890 0.275 ;
        RECT  5.520 -0.115 5.770 0.115 ;
        RECT  5.400 -0.115 5.520 0.145 ;
        RECT  4.560 -0.115 5.400 0.115 ;
        RECT  4.440 -0.115 4.560 0.200 ;
        RECT  3.760 -0.115 4.440 0.115 ;
        RECT  3.640 -0.115 3.760 0.220 ;
        RECT  2.600 -0.115 3.640 0.115 ;
        RECT  2.480 -0.115 2.600 0.125 ;
        RECT  2.200 -0.115 2.480 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 1.145 7.000 1.375 ;
        RECT  6.870 0.675 6.950 1.375 ;
        RECT  6.585 1.145 6.870 1.375 ;
        RECT  6.515 0.975 6.585 1.375 ;
        RECT  6.250 1.145 6.515 1.375 ;
        RECT  6.130 1.025 6.250 1.375 ;
        RECT  5.890 1.145 6.130 1.375 ;
        RECT  5.770 1.025 5.890 1.375 ;
        RECT  5.520 1.145 5.770 1.375 ;
        RECT  5.400 1.120 5.520 1.375 ;
        RECT  5.140 1.145 5.400 1.375 ;
        RECT  5.020 1.120 5.140 1.375 ;
        RECT  4.760 1.145 5.020 1.375 ;
        RECT  4.640 1.120 4.760 1.375 ;
        RECT  3.825 1.145 4.640 1.375 ;
        RECT  3.705 1.060 3.825 1.375 ;
        RECT  2.640 1.145 3.705 1.375 ;
        RECT  2.520 1.135 2.640 1.375 ;
        RECT  2.230 1.145 2.520 1.375 ;
        RECT  2.110 1.135 2.230 1.375 ;
        RECT  0.125 1.145 2.110 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.405 0.355 6.475 0.465 ;
        RECT  6.405 0.765 6.475 0.905 ;
        RECT  6.335 0.185 6.405 0.465 ;
        RECT  6.335 0.765 6.405 1.065 ;
        RECT  5.985 0.705 6.060 0.805 ;
        RECT  5.985 0.185 6.045 0.465 ;
        RECT  5.615 0.185 5.635 0.465 ;
        RECT  5.600 0.705 5.635 0.805 ;
        RECT  6.220 0.545 6.370 0.615 ;
        RECT  6.150 0.545 6.220 0.955 ;
        RECT  5.660 0.885 6.150 0.955 ;
        RECT  5.590 0.885 5.660 1.050 ;
        RECT  5.515 0.545 5.595 0.615 ;
        RECT  4.500 0.980 5.590 1.050 ;
        RECT  5.445 0.215 5.515 0.910 ;
        RECT  5.020 0.215 5.445 0.285 ;
        RECT  4.640 0.840 5.445 0.910 ;
        RECT  5.030 0.355 5.130 0.630 ;
        RECT  4.935 0.355 5.030 0.425 ;
        RECT  4.865 0.270 4.935 0.425 ;
        RECT  4.185 0.270 4.865 0.340 ;
        RECT  4.570 0.660 4.640 0.910 ;
        RECT  4.500 0.410 4.590 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.995 0.980 4.430 1.050 ;
        RECT  4.250 0.630 4.350 0.910 ;
        RECT  4.185 0.630 4.250 0.700 ;
        RECT  4.115 0.270 4.185 0.700 ;
        RECT  4.020 0.780 4.150 0.850 ;
        RECT  3.940 0.205 4.045 0.275 ;
        RECT  3.950 0.435 4.020 0.850 ;
        RECT  3.925 0.920 3.995 1.050 ;
        RECT  3.500 0.435 3.950 0.505 ;
        RECT  3.870 0.205 3.940 0.365 ;
        RECT  3.590 0.920 3.925 0.990 ;
        RECT  3.755 0.615 3.880 0.685 ;
        RECT  3.420 0.295 3.870 0.365 ;
        RECT  3.405 0.780 3.790 0.850 ;
        RECT  3.700 0.615 3.755 0.700 ;
        RECT  3.240 0.630 3.700 0.700 ;
        RECT  3.520 0.920 3.590 1.065 ;
        RECT  3.220 0.995 3.520 1.065 ;
        RECT  3.380 0.435 3.500 0.560 ;
        RECT  3.350 0.195 3.420 0.365 ;
        RECT  3.335 0.780 3.405 0.925 ;
        RECT  3.320 0.195 3.350 0.265 ;
        RECT  3.200 0.185 3.320 0.265 ;
        RECT  3.170 0.345 3.240 0.780 ;
        RECT  3.150 0.855 3.220 1.065 ;
        RECT  3.090 0.345 3.170 0.415 ;
        RECT  3.120 0.710 3.170 0.780 ;
        RECT  1.905 0.855 3.150 0.925 ;
        RECT  2.910 0.995 3.030 1.075 ;
        RECT  0.370 0.195 3.020 0.265 ;
        RECT  2.935 0.395 3.005 0.785 ;
        RECT  2.785 0.395 2.935 0.465 ;
        RECT  2.740 0.685 2.935 0.785 ;
        RECT  0.485 0.995 2.910 1.065 ;
        RECT  2.715 0.345 2.785 0.465 ;
        RECT  2.655 0.545 2.750 0.615 ;
        RECT  2.585 0.545 2.655 0.785 ;
        RECT  2.345 0.715 2.585 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCND4BWP

MACRO SEDFCNQD0BWP
    CLASS CORE ;
    FOREIGN SEDFCNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.330 5.565 0.905 ;
        RECT  5.475 0.330 5.495 0.450 ;
        RECT  5.475 0.765 5.495 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0348 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0176 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.295 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.495 4.865 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 -0.115 5.600 0.115 ;
        RECT  5.295 -0.115 5.365 0.450 ;
        RECT  4.780 -0.115 5.295 0.115 ;
        RECT  4.660 -0.115 4.780 0.200 ;
        RECT  3.690 -0.115 4.660 0.115 ;
        RECT  3.620 -0.115 3.690 0.265 ;
        RECT  2.580 -0.115 3.620 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 1.145 5.600 1.375 ;
        RECT  5.285 0.765 5.355 1.375 ;
        RECT  5.115 1.145 5.285 1.375 ;
        RECT  5.045 0.980 5.115 1.375 ;
        RECT  4.745 1.145 5.045 1.375 ;
        RECT  4.675 0.980 4.745 1.375 ;
        RECT  3.785 1.145 4.675 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.215 0.545 5.425 0.615 ;
        RECT  5.145 0.210 5.215 0.910 ;
        RECT  5.060 0.210 5.145 0.280 ;
        RECT  4.925 0.840 5.145 0.910 ;
        RECT  4.975 0.355 5.045 0.640 ;
        RECT  4.865 0.355 4.975 0.425 ;
        RECT  4.855 0.840 4.925 1.075 ;
        RECT  4.795 0.270 4.865 0.425 ;
        RECT  4.640 0.840 4.855 0.910 ;
        RECT  4.200 0.270 4.795 0.340 ;
        RECT  4.570 0.640 4.640 0.910 ;
        RECT  4.500 0.410 4.570 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.935 0.980 4.430 1.050 ;
        RECT  4.225 0.630 4.295 0.910 ;
        RECT  4.200 0.630 4.225 0.700 ;
        RECT  4.130 0.270 4.200 0.700 ;
        RECT  4.080 0.375 4.130 0.445 ;
        RECT  3.990 0.780 4.110 0.850 ;
        RECT  3.830 0.200 4.060 0.270 ;
        RECT  3.920 0.350 3.990 0.850 ;
        RECT  3.865 0.920 3.935 1.050 ;
        RECT  3.915 0.350 3.920 0.560 ;
        RECT  3.320 0.490 3.915 0.560 ;
        RECT  3.550 0.920 3.865 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.760 0.200 3.830 0.420 ;
        RECT  3.380 0.350 3.760 0.420 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.310 0.195 3.380 0.420 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.880 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  2.030 0.685 2.060 0.785 ;
        RECT  1.965 0.480 2.030 0.785 ;
        RECT  1.960 0.340 1.965 0.785 ;
        RECT  1.895 0.340 1.960 0.550 ;
        RECT  1.495 0.480 1.895 0.550 ;
        RECT  1.810 0.635 1.880 0.925 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.570 0.635 1.810 0.705 ;
        RECT  1.670 0.790 1.740 0.925 ;
        RECT  0.930 0.855 1.670 0.925 ;
        RECT  1.425 0.480 1.495 0.765 ;
        RECT  1.030 0.695 1.425 0.765 ;
        RECT  0.700 0.515 0.940 0.615 ;
        RECT  0.630 0.365 0.700 0.925 ;
        RECT  0.570 0.365 0.630 0.435 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCNQD0BWP

MACRO SEDFCNQD1BWP
    CLASS CORE ;
    FOREIGN SEDFCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.185 5.565 1.045 ;
        RECT  5.475 0.185 5.495 0.465 ;
        RECT  5.475 0.735 5.495 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.495 4.865 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 -0.115 5.600 0.115 ;
        RECT  5.295 -0.115 5.365 0.465 ;
        RECT  4.780 -0.115 5.295 0.115 ;
        RECT  4.660 -0.115 4.780 0.200 ;
        RECT  3.690 -0.115 4.660 0.115 ;
        RECT  3.620 -0.115 3.690 0.265 ;
        RECT  2.580 -0.115 3.620 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 1.145 5.600 1.375 ;
        RECT  5.285 0.735 5.355 1.375 ;
        RECT  4.745 1.145 5.285 1.375 ;
        RECT  4.675 0.980 4.745 1.375 ;
        RECT  3.785 1.145 4.675 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.215 0.545 5.425 0.615 ;
        RECT  5.145 0.205 5.215 0.910 ;
        RECT  5.070 0.205 5.145 0.275 ;
        RECT  4.925 0.840 5.145 0.910 ;
        RECT  4.975 0.355 5.045 0.640 ;
        RECT  4.865 0.355 4.975 0.425 ;
        RECT  4.855 0.840 4.925 1.075 ;
        RECT  4.795 0.270 4.865 0.425 ;
        RECT  4.640 0.840 4.855 0.910 ;
        RECT  4.200 0.270 4.795 0.340 ;
        RECT  4.570 0.640 4.640 0.910 ;
        RECT  4.500 0.410 4.570 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.935 0.980 4.430 1.050 ;
        RECT  4.225 0.630 4.295 0.910 ;
        RECT  4.200 0.630 4.225 0.700 ;
        RECT  4.130 0.270 4.200 0.700 ;
        RECT  4.080 0.375 4.130 0.445 ;
        RECT  3.990 0.780 4.110 0.850 ;
        RECT  3.830 0.200 4.060 0.270 ;
        RECT  3.920 0.350 3.990 0.850 ;
        RECT  3.865 0.920 3.935 1.050 ;
        RECT  3.915 0.350 3.920 0.560 ;
        RECT  3.320 0.490 3.915 0.560 ;
        RECT  3.550 0.920 3.865 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.760 0.200 3.830 0.420 ;
        RECT  3.380 0.350 3.760 0.420 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.310 0.195 3.380 0.420 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.905 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCNQD1BWP

MACRO SEDFCNQD2BWP
    CLASS CORE ;
    FOREIGN SEDFCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.505 0.355 5.565 0.805 ;
        RECT  5.495 0.185 5.505 1.035 ;
        RECT  5.435 0.185 5.495 0.465 ;
        RECT  5.435 0.735 5.495 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.345 2.505 0.475 ;
        RECT  2.415 0.345 2.490 0.635 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0384 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.495 4.865 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.300 ;
        RECT  5.325 -0.115 5.610 0.115 ;
        RECT  5.255 -0.115 5.325 0.465 ;
        RECT  4.740 -0.115 5.255 0.115 ;
        RECT  4.620 -0.115 4.740 0.200 ;
        RECT  3.690 -0.115 4.620 0.115 ;
        RECT  3.620 -0.115 3.690 0.265 ;
        RECT  2.580 -0.115 3.620 0.115 ;
        RECT  2.460 -0.115 2.580 0.125 ;
        RECT  2.200 -0.115 2.460 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.895 5.690 1.375 ;
        RECT  5.325 1.145 5.610 1.375 ;
        RECT  5.255 0.745 5.325 1.375 ;
        RECT  5.105 1.145 5.255 1.375 ;
        RECT  5.035 0.980 5.105 1.375 ;
        RECT  4.745 1.145 5.035 1.375 ;
        RECT  4.675 0.980 4.745 1.375 ;
        RECT  3.785 1.145 4.675 1.375 ;
        RECT  3.665 1.060 3.785 1.375 ;
        RECT  2.600 1.145 3.665 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.280 1.145 2.480 1.375 ;
        RECT  2.160 1.135 2.280 1.375 ;
        RECT  0.125 1.145 2.160 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.185 0.545 5.420 0.615 ;
        RECT  5.115 0.205 5.185 0.910 ;
        RECT  5.030 0.205 5.115 0.275 ;
        RECT  4.925 0.840 5.115 0.910 ;
        RECT  4.965 0.355 5.035 0.640 ;
        RECT  4.865 0.355 4.965 0.425 ;
        RECT  4.855 0.840 4.925 1.075 ;
        RECT  4.795 0.270 4.865 0.425 ;
        RECT  4.640 0.840 4.855 0.910 ;
        RECT  4.200 0.270 4.795 0.340 ;
        RECT  4.570 0.640 4.640 0.910 ;
        RECT  4.500 0.410 4.570 0.480 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.935 0.980 4.430 1.050 ;
        RECT  4.225 0.630 4.295 0.910 ;
        RECT  4.200 0.630 4.225 0.700 ;
        RECT  4.130 0.270 4.200 0.700 ;
        RECT  4.080 0.375 4.130 0.445 ;
        RECT  3.990 0.780 4.110 0.850 ;
        RECT  3.830 0.205 4.060 0.275 ;
        RECT  3.920 0.350 3.990 0.850 ;
        RECT  3.865 0.920 3.935 1.050 ;
        RECT  3.915 0.350 3.920 0.560 ;
        RECT  3.320 0.490 3.915 0.560 ;
        RECT  3.550 0.920 3.865 0.990 ;
        RECT  3.200 0.630 3.840 0.700 ;
        RECT  3.760 0.205 3.830 0.420 ;
        RECT  3.380 0.350 3.760 0.420 ;
        RECT  3.345 0.780 3.730 0.850 ;
        RECT  3.480 0.920 3.550 1.065 ;
        RECT  3.160 0.995 3.480 1.065 ;
        RECT  3.310 0.195 3.380 0.420 ;
        RECT  3.275 0.780 3.345 0.925 ;
        RECT  3.280 0.195 3.310 0.265 ;
        RECT  3.160 0.185 3.280 0.265 ;
        RECT  3.130 0.345 3.200 0.780 ;
        RECT  3.090 0.855 3.160 1.065 ;
        RECT  3.050 0.345 3.130 0.415 ;
        RECT  3.060 0.710 3.130 0.780 ;
        RECT  1.905 0.855 3.090 0.925 ;
        RECT  0.370 0.195 2.980 0.265 ;
        RECT  2.860 0.995 2.980 1.075 ;
        RECT  2.895 0.360 2.965 0.785 ;
        RECT  2.650 0.360 2.895 0.440 ;
        RECT  2.700 0.685 2.895 0.785 ;
        RECT  0.485 0.995 2.860 1.065 ;
        RECT  2.630 0.545 2.700 0.615 ;
        RECT  2.560 0.545 2.630 0.785 ;
        RECT  2.345 0.715 2.560 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCNQD2BWP

MACRO SEDFCNQD4BWP
    CLASS CORE ;
    FOREIGN SEDFCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0300 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.425 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.185 6.065 0.465 ;
        RECT  6.055 0.765 6.065 1.065 ;
        RECT  5.995 0.185 6.055 1.065 ;
        RECT  5.845 0.355 5.995 0.905 ;
        RECT  5.685 0.355 5.845 0.465 ;
        RECT  5.685 0.765 5.845 0.905 ;
        RECT  5.615 0.185 5.685 0.465 ;
        RECT  5.615 0.765 5.685 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0368 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.470 2.205 0.770 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0240 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.515 0.630 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.0672 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.495 5.375 0.640 ;
        RECT  5.215 0.495 5.285 0.770 ;
        RECT  4.865 0.700 5.215 0.770 ;
        RECT  4.785 0.495 4.865 0.770 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.465 ;
        RECT  5.900 -0.115 6.170 0.115 ;
        RECT  5.780 -0.115 5.900 0.275 ;
        RECT  5.520 -0.115 5.780 0.115 ;
        RECT  5.400 -0.115 5.520 0.145 ;
        RECT  4.560 -0.115 5.400 0.115 ;
        RECT  4.440 -0.115 4.560 0.200 ;
        RECT  3.760 -0.115 4.440 0.115 ;
        RECT  3.640 -0.115 3.760 0.220 ;
        RECT  2.600 -0.115 3.640 0.115 ;
        RECT  2.480 -0.115 2.600 0.125 ;
        RECT  2.200 -0.115 2.480 0.115 ;
        RECT  2.080 -0.115 2.200 0.125 ;
        RECT  0.840 -0.115 2.080 0.115 ;
        RECT  0.720 -0.115 0.840 0.125 ;
        RECT  0.140 -0.115 0.720 0.115 ;
        RECT  0.040 -0.115 0.140 0.285 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.675 6.250 1.375 ;
        RECT  5.875 1.145 6.170 1.375 ;
        RECT  5.805 0.975 5.875 1.375 ;
        RECT  5.495 1.145 5.805 1.375 ;
        RECT  5.425 0.980 5.495 1.375 ;
        RECT  5.115 1.145 5.425 1.375 ;
        RECT  5.045 0.980 5.115 1.375 ;
        RECT  4.735 1.145 5.045 1.375 ;
        RECT  4.665 0.980 4.735 1.375 ;
        RECT  3.825 1.145 4.665 1.375 ;
        RECT  3.705 1.060 3.825 1.375 ;
        RECT  2.640 1.145 3.705 1.375 ;
        RECT  2.520 1.135 2.640 1.375 ;
        RECT  2.230 1.145 2.520 1.375 ;
        RECT  2.110 1.135 2.230 1.375 ;
        RECT  0.125 1.145 2.110 1.375 ;
        RECT  0.055 0.900 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.685 0.355 5.775 0.465 ;
        RECT  5.685 0.765 5.775 0.905 ;
        RECT  5.615 0.185 5.685 0.465 ;
        RECT  5.615 0.765 5.685 1.065 ;
        RECT  5.515 0.545 5.710 0.615 ;
        RECT  5.445 0.215 5.515 0.910 ;
        RECT  5.020 0.215 5.445 0.285 ;
        RECT  5.305 0.840 5.445 0.910 ;
        RECT  5.235 0.840 5.305 1.075 ;
        RECT  4.925 0.840 5.235 0.910 ;
        RECT  5.030 0.355 5.130 0.630 ;
        RECT  4.935 0.355 5.030 0.425 ;
        RECT  4.865 0.270 4.935 0.425 ;
        RECT  4.855 0.840 4.925 1.075 ;
        RECT  4.185 0.270 4.865 0.340 ;
        RECT  4.640 0.840 4.855 0.910 ;
        RECT  4.570 0.660 4.640 0.910 ;
        RECT  4.500 0.410 4.590 0.480 ;
        RECT  4.500 0.980 4.570 1.050 ;
        RECT  4.430 0.410 4.500 1.050 ;
        RECT  4.270 0.475 4.430 0.545 ;
        RECT  3.995 0.980 4.430 1.050 ;
        RECT  4.250 0.630 4.350 0.910 ;
        RECT  4.185 0.630 4.250 0.700 ;
        RECT  4.115 0.270 4.185 0.700 ;
        RECT  4.020 0.780 4.150 0.850 ;
        RECT  3.940 0.205 4.045 0.275 ;
        RECT  3.950 0.435 4.020 0.850 ;
        RECT  3.925 0.920 3.995 1.050 ;
        RECT  3.500 0.435 3.950 0.505 ;
        RECT  3.870 0.205 3.940 0.365 ;
        RECT  3.590 0.920 3.925 0.990 ;
        RECT  3.755 0.615 3.880 0.685 ;
        RECT  3.420 0.295 3.870 0.365 ;
        RECT  3.405 0.780 3.790 0.850 ;
        RECT  3.700 0.615 3.755 0.700 ;
        RECT  3.240 0.630 3.700 0.700 ;
        RECT  3.520 0.920 3.590 1.065 ;
        RECT  3.220 0.995 3.520 1.065 ;
        RECT  3.380 0.435 3.500 0.560 ;
        RECT  3.350 0.195 3.420 0.365 ;
        RECT  3.335 0.780 3.405 0.925 ;
        RECT  3.320 0.195 3.350 0.265 ;
        RECT  3.200 0.185 3.320 0.265 ;
        RECT  3.170 0.345 3.240 0.780 ;
        RECT  3.150 0.855 3.220 1.065 ;
        RECT  3.090 0.345 3.170 0.415 ;
        RECT  3.120 0.710 3.170 0.780 ;
        RECT  1.905 0.855 3.150 0.925 ;
        RECT  2.910 0.995 3.030 1.075 ;
        RECT  0.370 0.195 3.020 0.265 ;
        RECT  2.935 0.395 3.005 0.785 ;
        RECT  2.785 0.395 2.935 0.465 ;
        RECT  2.740 0.685 2.935 0.785 ;
        RECT  0.485 0.995 2.910 1.065 ;
        RECT  2.715 0.345 2.785 0.465 ;
        RECT  2.655 0.545 2.750 0.615 ;
        RECT  2.585 0.545 2.655 0.785 ;
        RECT  2.345 0.715 2.585 0.785 ;
        RECT  2.275 0.345 2.345 0.785 ;
        RECT  1.975 0.480 2.045 0.775 ;
        RECT  1.965 0.480 1.975 0.550 ;
        RECT  1.895 0.340 1.965 0.550 ;
        RECT  1.835 0.635 1.905 0.925 ;
        RECT  1.515 0.480 1.895 0.550 ;
        RECT  1.590 0.635 1.835 0.705 ;
        RECT  0.930 0.340 1.810 0.410 ;
        RECT  1.695 0.790 1.765 0.925 ;
        RECT  0.930 0.855 1.695 0.925 ;
        RECT  1.445 0.480 1.515 0.780 ;
        RECT  1.090 0.710 1.445 0.780 ;
        RECT  1.020 0.660 1.090 0.780 ;
        RECT  0.700 0.515 0.950 0.585 ;
        RECT  0.630 0.345 0.700 0.925 ;
        RECT  0.570 0.345 0.630 0.415 ;
        RECT  0.375 0.705 0.630 0.775 ;
        RECT  0.570 0.855 0.630 0.925 ;
        RECT  0.415 0.895 0.485 1.065 ;
    END
END SEDFCNQD4BWP

MACRO SEDFD0BWP
    CLASS CORE ;
    FOREIGN SEDFD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0268 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.225 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.350 5.285 0.905 ;
        RECT  5.195 0.350 5.215 0.470 ;
        RECT  5.200 0.760 5.215 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.215 5.005 0.485 ;
        RECT  4.885 0.350 4.935 0.485 ;
        RECT  4.815 0.350 4.885 0.895 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.100 -0.115 5.320 0.115 ;
        RECT  4.980 -0.115 5.100 0.145 ;
        RECT  4.495 -0.115 4.980 0.115 ;
        RECT  4.425 -0.115 4.495 0.280 ;
        RECT  3.660 -0.115 4.425 0.115 ;
        RECT  3.540 -0.115 3.660 0.125 ;
        RECT  2.720 -0.115 3.540 0.115 ;
        RECT  2.600 -0.115 2.720 0.125 ;
        RECT  2.210 -0.115 2.600 0.115 ;
        RECT  2.090 -0.115 2.210 0.125 ;
        RECT  1.420 -0.115 2.090 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  1.060 -0.115 1.300 0.115 ;
        RECT  0.940 -0.115 1.060 0.150 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.080 1.145 5.320 1.375 ;
        RECT  4.960 1.135 5.080 1.375 ;
        RECT  4.560 1.145 4.960 1.375 ;
        RECT  4.440 1.135 4.560 1.375 ;
        RECT  3.700 1.145 4.440 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  2.740 1.145 3.580 1.375 ;
        RECT  2.620 1.135 2.740 1.375 ;
        RECT  2.180 1.145 2.620 1.375 ;
        RECT  2.060 1.135 2.180 1.375 ;
        RECT  0.330 1.145 2.060 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.130 0.520 5.145 0.710 ;
        RECT  5.075 0.520 5.130 1.065 ;
        RECT  5.060 0.640 5.075 1.065 ;
        RECT  4.745 0.995 5.060 1.065 ;
        RECT  4.675 0.365 4.745 1.065 ;
        RECT  4.395 0.365 4.675 0.435 ;
        RECT  4.635 0.840 4.675 1.065 ;
        RECT  3.880 0.995 4.635 1.065 ;
        RECT  4.550 0.520 4.595 0.640 ;
        RECT  4.480 0.520 4.550 0.925 ;
        RECT  4.030 0.855 4.480 0.925 ;
        RECT  4.325 0.365 4.395 0.640 ;
        RECT  4.180 0.715 4.270 0.785 ;
        RECT  4.110 0.195 4.180 0.785 ;
        RECT  3.995 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.925 ;
        RECT  3.855 0.185 3.995 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.065 ;
        RECT  3.295 0.195 3.855 0.265 ;
        RECT  3.780 0.335 3.820 0.455 ;
        RECT  3.555 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.695 0.520 3.750 0.640 ;
        RECT  3.625 0.340 3.695 0.640 ;
        RECT  3.285 0.340 3.625 0.410 ;
        RECT  3.485 0.520 3.555 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.545 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.545 1.765 0.615 ;
        RECT  1.530 0.685 1.680 0.755 ;
        RECT  1.460 0.685 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.640 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.570 0.675 0.640 ;
        RECT  0.345 0.570 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFD0BWP

MACRO SEDFD1BWP
    CLASS CORE ;
    FOREIGN SEDFD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.210 5.285 1.065 ;
        RECT  5.195 0.210 5.215 0.470 ;
        RECT  5.195 0.760 5.215 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.885 0.215 5.005 0.485 ;
        RECT  4.815 0.215 4.885 0.895 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.100 -0.115 5.320 0.115 ;
        RECT  4.980 -0.115 5.100 0.145 ;
        RECT  4.495 -0.115 4.980 0.115 ;
        RECT  4.425 -0.115 4.495 0.280 ;
        RECT  3.660 -0.115 4.425 0.115 ;
        RECT  3.540 -0.115 3.660 0.125 ;
        RECT  2.720 -0.115 3.540 0.115 ;
        RECT  2.600 -0.115 2.720 0.125 ;
        RECT  2.210 -0.115 2.600 0.115 ;
        RECT  2.090 -0.115 2.210 0.125 ;
        RECT  1.420 -0.115 2.090 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  1.060 -0.115 1.300 0.115 ;
        RECT  0.940 -0.115 1.060 0.150 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.100 1.145 5.320 1.375 ;
        RECT  4.980 1.140 5.100 1.375 ;
        RECT  4.560 1.145 4.980 1.375 ;
        RECT  4.440 1.135 4.560 1.375 ;
        RECT  3.700 1.145 4.440 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  2.740 1.145 3.580 1.375 ;
        RECT  2.620 1.135 2.740 1.375 ;
        RECT  2.180 1.145 2.620 1.375 ;
        RECT  2.060 1.135 2.180 1.375 ;
        RECT  0.330 1.145 2.060 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.125 0.520 5.145 0.710 ;
        RECT  5.075 0.520 5.125 1.065 ;
        RECT  5.055 0.640 5.075 1.065 ;
        RECT  4.745 0.995 5.055 1.065 ;
        RECT  4.675 0.365 4.745 1.065 ;
        RECT  4.395 0.365 4.675 0.435 ;
        RECT  4.635 0.840 4.675 1.065 ;
        RECT  3.880 0.995 4.635 1.065 ;
        RECT  4.550 0.520 4.595 0.640 ;
        RECT  4.480 0.520 4.550 0.925 ;
        RECT  4.030 0.855 4.480 0.925 ;
        RECT  4.325 0.365 4.395 0.640 ;
        RECT  4.180 0.715 4.270 0.785 ;
        RECT  4.110 0.195 4.180 0.785 ;
        RECT  3.995 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.925 ;
        RECT  3.855 0.185 3.995 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.065 ;
        RECT  3.295 0.195 3.855 0.265 ;
        RECT  3.780 0.335 3.820 0.455 ;
        RECT  3.555 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.695 0.520 3.750 0.640 ;
        RECT  3.625 0.340 3.695 0.640 ;
        RECT  3.285 0.340 3.625 0.410 ;
        RECT  3.485 0.520 3.555 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.685 1.680 0.755 ;
        RECT  1.460 0.685 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFD1BWP

MACRO SEDFD2BWP
    CLASS CORE ;
    FOREIGN SEDFD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.365 0.355 5.425 0.820 ;
        RECT  5.355 0.185 5.365 1.035 ;
        RECT  5.295 0.185 5.355 0.465 ;
        RECT  5.295 0.735 5.355 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.215 5.005 0.790 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.550 0.300 ;
        RECT  5.185 -0.115 5.470 0.115 ;
        RECT  5.115 -0.115 5.185 0.465 ;
        RECT  4.850 -0.115 5.115 0.115 ;
        RECT  4.730 -0.115 4.850 0.280 ;
        RECT  4.455 -0.115 4.730 0.115 ;
        RECT  4.385 -0.115 4.455 0.280 ;
        RECT  3.640 -0.115 4.385 0.115 ;
        RECT  3.520 -0.115 3.640 0.125 ;
        RECT  2.720 -0.115 3.520 0.115 ;
        RECT  2.600 -0.115 2.720 0.125 ;
        RECT  2.210 -0.115 2.600 0.115 ;
        RECT  2.090 -0.115 2.210 0.125 ;
        RECT  1.420 -0.115 2.090 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  1.060 -0.115 1.300 0.115 ;
        RECT  0.940 -0.115 1.060 0.150 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 1.145 5.600 1.375 ;
        RECT  5.470 0.905 5.550 1.375 ;
        RECT  5.210 1.145 5.470 1.375 ;
        RECT  5.090 1.010 5.210 1.375 ;
        RECT  4.850 1.145 5.090 1.375 ;
        RECT  4.730 1.010 4.850 1.375 ;
        RECT  4.520 1.145 4.730 1.375 ;
        RECT  4.400 1.135 4.520 1.375 ;
        RECT  3.700 1.145 4.400 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  2.740 1.145 3.580 1.375 ;
        RECT  2.620 1.135 2.740 1.375 ;
        RECT  2.180 1.145 2.620 1.375 ;
        RECT  2.060 1.135 2.180 1.375 ;
        RECT  0.330 1.145 2.060 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.170 0.545 5.280 0.615 ;
        RECT  5.100 0.545 5.170 0.940 ;
        RECT  4.865 0.870 5.100 0.940 ;
        RECT  4.795 0.365 4.865 0.940 ;
        RECT  4.355 0.365 4.795 0.435 ;
        RECT  4.645 0.840 4.795 0.940 ;
        RECT  4.505 0.545 4.725 0.615 ;
        RECT  4.575 0.840 4.645 1.065 ;
        RECT  3.880 0.995 4.575 1.065 ;
        RECT  4.435 0.545 4.505 0.925 ;
        RECT  4.030 0.855 4.435 0.925 ;
        RECT  4.285 0.365 4.355 0.620 ;
        RECT  4.180 0.700 4.240 0.770 ;
        RECT  4.110 0.195 4.180 0.770 ;
        RECT  3.975 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.925 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.065 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.820 0.455 ;
        RECT  3.550 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.690 0.520 3.730 0.640 ;
        RECT  3.620 0.340 3.690 0.640 ;
        RECT  3.285 0.340 3.620 0.410 ;
        RECT  3.480 0.520 3.550 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.685 1.680 0.755 ;
        RECT  1.460 0.685 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFD2BWP

MACRO SEDFD4BWP
    CLASS CORE ;
    FOREIGN SEDFD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.415 0.185 6.485 0.465 ;
        RECT  6.415 0.765 6.485 1.065 ;
        RECT  6.335 0.355 6.415 0.465 ;
        RECT  6.335 0.765 6.415 0.905 ;
        RECT  6.125 0.355 6.335 0.905 ;
        RECT  6.055 0.185 6.125 0.465 ;
        RECT  6.055 0.765 6.125 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.695 5.780 0.795 ;
        RECT  5.695 0.185 5.765 0.485 ;
        RECT  5.635 0.355 5.695 0.485 ;
        RECT  5.425 0.355 5.635 0.795 ;
        RECT  5.385 0.355 5.425 0.485 ;
        RECT  5.300 0.695 5.425 0.795 ;
        RECT  5.315 0.185 5.385 0.485 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.670 -0.115 6.720 0.115 ;
        RECT  6.590 -0.115 6.670 0.465 ;
        RECT  6.330 -0.115 6.590 0.115 ;
        RECT  6.210 -0.115 6.330 0.275 ;
        RECT  5.945 -0.115 6.210 0.115 ;
        RECT  5.875 -0.115 5.945 0.465 ;
        RECT  5.600 -0.115 5.875 0.115 ;
        RECT  5.480 -0.115 5.600 0.275 ;
        RECT  5.205 -0.115 5.480 0.115 ;
        RECT  5.135 -0.115 5.205 0.305 ;
        RECT  4.870 -0.115 5.135 0.115 ;
        RECT  4.750 -0.115 4.870 0.280 ;
        RECT  4.040 -0.115 4.750 0.115 ;
        RECT  3.920 -0.115 4.040 0.130 ;
        RECT  3.640 -0.115 3.920 0.115 ;
        RECT  3.520 -0.115 3.640 0.125 ;
        RECT  2.740 -0.115 3.520 0.115 ;
        RECT  2.620 -0.115 2.740 0.130 ;
        RECT  2.210 -0.115 2.620 0.115 ;
        RECT  2.090 -0.115 2.210 0.125 ;
        RECT  1.420 -0.115 2.090 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  1.060 -0.115 1.300 0.115 ;
        RECT  0.940 -0.115 1.060 0.150 ;
        RECT  0.330 -0.115 0.940 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.145 6.720 1.375 ;
        RECT  6.590 0.685 6.670 1.375 ;
        RECT  6.305 1.145 6.590 1.375 ;
        RECT  6.235 0.975 6.305 1.375 ;
        RECT  5.970 1.145 6.235 1.375 ;
        RECT  5.850 1.005 5.970 1.375 ;
        RECT  5.600 1.145 5.850 1.375 ;
        RECT  5.480 1.005 5.600 1.375 ;
        RECT  5.230 1.145 5.480 1.375 ;
        RECT  5.110 1.005 5.230 1.375 ;
        RECT  4.860 1.145 5.110 1.375 ;
        RECT  4.740 1.120 4.860 1.375 ;
        RECT  4.070 1.145 4.740 1.375 ;
        RECT  3.950 1.040 4.070 1.375 ;
        RECT  3.680 1.145 3.950 1.375 ;
        RECT  3.560 1.040 3.680 1.375 ;
        RECT  2.740 1.145 3.560 1.375 ;
        RECT  2.620 1.135 2.740 1.375 ;
        RECT  2.180 1.145 2.620 1.375 ;
        RECT  2.060 1.135 2.180 1.375 ;
        RECT  0.330 1.145 2.060 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.415 0.185 6.485 0.465 ;
        RECT  6.415 0.765 6.485 1.065 ;
        RECT  6.405 0.355 6.415 0.465 ;
        RECT  6.405 0.765 6.415 0.905 ;
        RECT  5.705 0.695 5.780 0.795 ;
        RECT  5.705 0.185 5.765 0.485 ;
        RECT  5.315 0.185 5.355 0.485 ;
        RECT  5.300 0.695 5.355 0.795 ;
        RECT  5.930 0.545 6.040 0.615 ;
        RECT  5.860 0.545 5.930 0.935 ;
        RECT  5.180 0.865 5.860 0.935 ;
        RECT  5.110 0.375 5.180 0.935 ;
        RECT  5.025 0.375 5.110 0.445 ;
        RECT  5.025 0.865 5.110 0.935 ;
        RECT  4.955 0.185 5.025 0.445 ;
        RECT  4.955 0.520 5.025 0.790 ;
        RECT  4.955 0.865 5.025 1.050 ;
        RECT  4.755 0.375 4.955 0.445 ;
        RECT  4.790 0.720 4.955 0.790 ;
        RECT  4.235 0.980 4.955 1.050 ;
        RECT  4.720 0.720 4.790 0.910 ;
        RECT  4.685 0.375 4.755 0.640 ;
        RECT  4.390 0.840 4.720 0.910 ;
        RECT  4.530 0.700 4.600 0.770 ;
        RECT  4.460 0.200 4.530 0.770 ;
        RECT  4.330 0.200 4.460 0.270 ;
        RECT  4.320 0.340 4.390 0.910 ;
        RECT  4.190 0.185 4.330 0.270 ;
        RECT  4.290 0.340 4.320 0.460 ;
        RECT  4.210 0.750 4.250 0.820 ;
        RECT  4.165 0.900 4.235 1.050 ;
        RECT  4.140 0.345 4.210 0.820 ;
        RECT  3.295 0.200 4.190 0.270 ;
        RECT  3.435 0.900 4.165 0.970 ;
        RECT  3.730 0.345 4.140 0.415 ;
        RECT  3.560 0.750 4.140 0.820 ;
        RECT  3.285 0.515 3.930 0.585 ;
        RECT  3.440 0.665 3.560 0.820 ;
        RECT  3.365 0.900 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.200 3.110 0.270 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.200 1.775 0.460 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.685 1.680 0.755 ;
        RECT  1.460 0.685 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFD4BWP

MACRO SEDFKCND0BWP
    CLASS CORE ;
    FOREIGN SEDFKCND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.355 2.205 0.625 ;
        RECT  2.100 0.555 2.135 0.625 ;
        RECT  1.980 0.555 2.100 0.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.635 2.765 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.330 5.705 0.905 ;
        RECT  5.615 0.330 5.635 0.450 ;
        RECT  5.615 0.775 5.635 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.330 0.355 5.400 0.905 ;
        RECT  5.215 0.355 5.330 0.485 ;
        RECT  5.215 0.775 5.330 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0256 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 3.045 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 -0.115 5.740 0.115 ;
        RECT  5.400 -0.115 5.520 0.140 ;
        RECT  4.940 -0.115 5.400 0.115 ;
        RECT  4.820 -0.115 4.940 0.140 ;
        RECT  4.085 -0.115 4.820 0.115 ;
        RECT  4.015 -0.115 4.085 0.420 ;
        RECT  3.175 -0.115 4.015 0.115 ;
        RECT  3.055 -0.115 3.175 0.125 ;
        RECT  2.840 -0.115 3.055 0.115 ;
        RECT  2.720 -0.115 2.840 0.125 ;
        RECT  2.010 -0.115 2.720 0.115 ;
        RECT  1.930 -0.115 2.010 0.455 ;
        RECT  1.470 -0.115 1.930 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.145 5.740 1.375 ;
        RECT  5.400 1.120 5.520 1.375 ;
        RECT  4.940 1.145 5.400 1.375 ;
        RECT  4.820 1.120 4.940 1.375 ;
        RECT  4.100 1.145 4.820 1.375 ;
        RECT  3.975 1.030 4.100 1.375 ;
        RECT  3.175 1.145 3.975 1.375 ;
        RECT  3.055 1.135 3.175 1.375 ;
        RECT  2.840 1.145 3.055 1.375 ;
        RECT  2.720 1.135 2.840 1.375 ;
        RECT  2.040 1.145 2.720 1.375 ;
        RECT  1.920 1.060 2.040 1.375 ;
        RECT  1.420 1.145 1.920 1.375 ;
        RECT  1.300 1.135 1.420 1.375 ;
        RECT  1.120 1.145 1.300 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.545 0.520 5.565 0.640 ;
        RECT  5.475 0.210 5.545 1.050 ;
        RECT  5.110 0.210 5.475 0.280 ;
        RECT  4.270 0.980 5.475 1.050 ;
        RECT  5.110 0.555 5.220 0.625 ;
        RECT  5.040 0.210 5.110 0.305 ;
        RECT  5.040 0.375 5.110 0.895 ;
        RECT  4.740 0.235 5.040 0.305 ;
        RECT  4.820 0.375 5.040 0.445 ;
        RECT  4.900 0.520 4.970 0.910 ;
        RECT  4.880 0.520 4.900 0.630 ;
        RECT  4.380 0.840 4.900 0.910 ;
        RECT  4.580 0.560 4.880 0.630 ;
        RECT  4.700 0.375 4.820 0.465 ;
        RECT  4.650 0.185 4.740 0.305 ;
        RECT  4.440 0.700 4.640 0.770 ;
        RECT  4.510 0.210 4.580 0.630 ;
        RECT  4.420 0.210 4.510 0.280 ;
        RECT  4.370 0.360 4.440 0.770 ;
        RECT  4.230 0.185 4.300 0.820 ;
        RECT  4.200 0.890 4.270 1.050 ;
        RECT  4.000 0.750 4.230 0.820 ;
        RECT  3.880 0.890 4.200 0.960 ;
        RECT  4.090 0.520 4.160 0.640 ;
        RECT  3.725 0.520 4.090 0.590 ;
        RECT  3.880 0.680 4.000 0.820 ;
        RECT  3.810 0.890 3.880 1.065 ;
        RECT  2.250 0.995 3.810 1.065 ;
        RECT  3.705 0.300 3.725 0.590 ;
        RECT  3.655 0.300 3.705 0.920 ;
        RECT  3.635 0.520 3.655 0.920 ;
        RECT  2.750 0.195 3.550 0.265 ;
        RECT  2.330 0.855 3.550 0.925 ;
        RECT  3.435 0.335 3.505 0.785 ;
        RECT  3.260 0.335 3.435 0.435 ;
        RECT  3.260 0.685 3.435 0.785 ;
        RECT  3.185 0.545 3.250 0.615 ;
        RECT  3.115 0.355 3.185 0.785 ;
        RECT  2.870 0.355 3.115 0.425 ;
        RECT  2.870 0.715 3.115 0.785 ;
        RECT  2.680 0.195 2.750 0.405 ;
        RECT  2.345 0.475 2.740 0.545 ;
        RECT  2.320 0.335 2.680 0.405 ;
        RECT  2.275 0.475 2.345 0.775 ;
        RECT  2.250 0.705 2.275 0.775 ;
        RECT  2.180 0.705 2.250 0.850 ;
        RECT  2.180 0.920 2.250 1.065 ;
        RECT  1.780 0.780 2.180 0.850 ;
        RECT  1.805 0.920 2.180 0.990 ;
        RECT  1.780 0.335 1.825 0.545 ;
        RECT  1.735 0.920 1.805 1.065 ;
        RECT  1.755 0.335 1.780 0.850 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.710 0.475 1.755 0.850 ;
        RECT  0.970 0.995 1.735 1.065 ;
        RECT  1.570 0.185 1.640 0.915 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.535 0.795 1.570 0.915 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.870 0.505 0.990 0.775 ;
        RECT  0.850 0.995 0.970 1.070 ;
        RECT  0.385 0.705 0.870 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCND0BWP

MACRO SEDFKCND1BWP
    CLASS CORE ;
    FOREIGN SEDFKCND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.185 5.845 1.045 ;
        RECT  5.755 0.185 5.775 0.465 ;
        RECT  5.755 0.740 5.775 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.470 0.355 5.540 0.905 ;
        RECT  5.355 0.355 5.470 0.485 ;
        RECT  5.355 0.775 5.470 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.115 5.880 0.115 ;
        RECT  5.540 -0.115 5.660 0.140 ;
        RECT  5.080 -0.115 5.540 0.115 ;
        RECT  4.960 -0.115 5.080 0.140 ;
        RECT  4.225 -0.115 4.960 0.115 ;
        RECT  4.155 -0.115 4.225 0.420 ;
        RECT  3.315 -0.115 4.155 0.115 ;
        RECT  3.195 -0.115 3.315 0.125 ;
        RECT  2.980 -0.115 3.195 0.115 ;
        RECT  2.860 -0.115 2.980 0.125 ;
        RECT  2.010 -0.115 2.860 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.145 5.880 1.375 ;
        RECT  5.540 1.120 5.660 1.375 ;
        RECT  5.080 1.145 5.540 1.375 ;
        RECT  4.960 1.120 5.080 1.375 ;
        RECT  4.240 1.145 4.960 1.375 ;
        RECT  4.115 1.030 4.240 1.375 ;
        RECT  3.315 1.145 4.115 1.375 ;
        RECT  3.195 1.135 3.315 1.375 ;
        RECT  2.940 1.145 3.195 1.375 ;
        RECT  2.820 1.135 2.940 1.375 ;
        RECT  2.100 1.145 2.820 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.685 0.520 5.705 0.640 ;
        RECT  5.615 0.210 5.685 1.050 ;
        RECT  5.250 0.210 5.615 0.280 ;
        RECT  4.410 0.980 5.615 1.050 ;
        RECT  5.250 0.555 5.350 0.625 ;
        RECT  5.180 0.210 5.250 0.305 ;
        RECT  5.180 0.375 5.250 0.895 ;
        RECT  4.880 0.235 5.180 0.305 ;
        RECT  4.960 0.375 5.180 0.445 ;
        RECT  5.040 0.520 5.110 0.910 ;
        RECT  5.020 0.520 5.040 0.630 ;
        RECT  4.520 0.840 5.040 0.910 ;
        RECT  4.720 0.560 5.020 0.630 ;
        RECT  4.840 0.375 4.960 0.465 ;
        RECT  4.790 0.185 4.880 0.305 ;
        RECT  4.580 0.700 4.780 0.770 ;
        RECT  4.650 0.210 4.720 0.630 ;
        RECT  4.560 0.210 4.650 0.280 ;
        RECT  4.510 0.360 4.580 0.770 ;
        RECT  4.370 0.185 4.440 0.820 ;
        RECT  4.340 0.890 4.410 1.050 ;
        RECT  4.140 0.750 4.370 0.820 ;
        RECT  4.020 0.890 4.340 0.960 ;
        RECT  4.230 0.520 4.300 0.640 ;
        RECT  3.865 0.520 4.230 0.590 ;
        RECT  4.020 0.680 4.140 0.820 ;
        RECT  3.950 0.890 4.020 1.065 ;
        RECT  2.290 0.995 3.950 1.065 ;
        RECT  3.845 0.300 3.865 0.590 ;
        RECT  3.795 0.300 3.845 0.920 ;
        RECT  3.775 0.520 3.795 0.920 ;
        RECT  2.385 0.195 3.690 0.265 ;
        RECT  2.390 0.855 3.690 0.925 ;
        RECT  3.575 0.335 3.645 0.785 ;
        RECT  3.400 0.335 3.575 0.435 ;
        RECT  3.400 0.685 3.575 0.785 ;
        RECT  3.325 0.545 3.390 0.615 ;
        RECT  3.255 0.355 3.325 0.785 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.715 3.255 0.785 ;
        RECT  2.835 0.335 2.905 0.785 ;
        RECT  2.470 0.335 2.835 0.405 ;
        RECT  2.610 0.715 2.835 0.785 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.195 2.385 0.410 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.065 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCND1BWP

MACRO SEDFKCND2BWP
    CLASS CORE ;
    FOREIGN SEDFKCND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.065 0.355 6.125 0.815 ;
        RECT  6.055 0.185 6.065 1.035 ;
        RECT  5.995 0.185 6.055 0.465 ;
        RECT  5.995 0.745 6.055 1.035 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.615 0.355 5.705 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.300 ;
        RECT  5.900 -0.115 6.170 0.115 ;
        RECT  5.780 -0.115 5.900 0.140 ;
        RECT  5.470 -0.115 5.780 0.115 ;
        RECT  5.350 -0.115 5.470 0.140 ;
        RECT  5.100 -0.115 5.350 0.115 ;
        RECT  4.980 -0.115 5.100 0.140 ;
        RECT  4.245 -0.115 4.980 0.115 ;
        RECT  4.175 -0.115 4.245 0.420 ;
        RECT  3.315 -0.115 4.175 0.115 ;
        RECT  3.195 -0.115 3.315 0.125 ;
        RECT  2.980 -0.115 3.195 0.115 ;
        RECT  2.860 -0.115 2.980 0.125 ;
        RECT  2.010 -0.115 2.860 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.905 6.250 1.375 ;
        RECT  5.900 1.145 6.170 1.375 ;
        RECT  5.780 1.120 5.900 1.375 ;
        RECT  5.470 1.145 5.780 1.375 ;
        RECT  5.350 1.120 5.470 1.375 ;
        RECT  5.100 1.145 5.350 1.375 ;
        RECT  4.980 1.120 5.100 1.375 ;
        RECT  4.260 1.145 4.980 1.375 ;
        RECT  4.135 1.030 4.260 1.375 ;
        RECT  3.315 1.145 4.135 1.375 ;
        RECT  3.195 1.135 3.315 1.375 ;
        RECT  2.940 1.145 3.195 1.375 ;
        RECT  2.820 1.135 2.940 1.375 ;
        RECT  2.100 1.145 2.820 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.890 0.545 5.980 0.615 ;
        RECT  5.820 0.210 5.890 1.050 ;
        RECT  5.270 0.210 5.820 0.280 ;
        RECT  4.430 0.980 5.820 1.050 ;
        RECT  5.440 0.385 5.510 0.875 ;
        RECT  4.860 0.385 5.440 0.455 ;
        RECT  5.160 0.805 5.440 0.875 ;
        RECT  5.200 0.210 5.270 0.305 ;
        RECT  4.900 0.235 5.200 0.305 ;
        RECT  4.970 0.545 5.180 0.615 ;
        RECT  4.900 0.545 4.970 0.910 ;
        RECT  4.810 0.185 4.900 0.305 ;
        RECT  4.740 0.545 4.900 0.615 ;
        RECT  4.540 0.840 4.900 0.910 ;
        RECT  4.600 0.700 4.800 0.770 ;
        RECT  4.670 0.210 4.740 0.615 ;
        RECT  4.580 0.210 4.670 0.280 ;
        RECT  4.530 0.360 4.600 0.770 ;
        RECT  4.390 0.185 4.460 0.820 ;
        RECT  4.360 0.890 4.430 1.050 ;
        RECT  4.160 0.750 4.390 0.820 ;
        RECT  4.020 0.890 4.360 0.960 ;
        RECT  4.250 0.520 4.320 0.640 ;
        RECT  3.865 0.520 4.250 0.590 ;
        RECT  4.040 0.680 4.160 0.820 ;
        RECT  3.950 0.890 4.020 1.065 ;
        RECT  2.290 0.995 3.950 1.065 ;
        RECT  3.845 0.300 3.865 0.590 ;
        RECT  3.795 0.300 3.845 0.920 ;
        RECT  3.775 0.520 3.795 0.920 ;
        RECT  2.385 0.195 3.690 0.265 ;
        RECT  2.390 0.855 3.690 0.925 ;
        RECT  3.575 0.335 3.645 0.785 ;
        RECT  3.400 0.335 3.575 0.435 ;
        RECT  3.400 0.685 3.575 0.785 ;
        RECT  3.325 0.545 3.390 0.615 ;
        RECT  3.255 0.355 3.325 0.785 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.715 3.255 0.785 ;
        RECT  2.835 0.335 2.905 0.785 ;
        RECT  2.470 0.335 2.835 0.405 ;
        RECT  2.610 0.715 2.835 0.785 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.195 2.385 0.410 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.065 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCND2BWP

MACRO SEDFKCND4BWP
    CLASS CORE ;
    FOREIGN SEDFKCND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.695 0.185 6.765 0.465 ;
        RECT  6.695 0.765 6.765 1.065 ;
        RECT  6.615 0.355 6.695 0.465 ;
        RECT  6.615 0.765 6.695 0.905 ;
        RECT  6.425 0.355 6.615 0.905 ;
        RECT  6.405 0.355 6.425 1.065 ;
        RECT  6.335 0.185 6.405 0.465 ;
        RECT  6.335 0.765 6.405 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.710 6.070 0.800 ;
        RECT  5.915 0.355 6.050 0.455 ;
        RECT  5.705 0.355 5.915 0.800 ;
        RECT  5.550 0.355 5.705 0.455 ;
        RECT  5.590 0.710 5.705 0.800 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 -0.115 7.000 0.115 ;
        RECT  6.870 -0.115 6.950 0.465 ;
        RECT  6.585 -0.115 6.870 0.115 ;
        RECT  6.515 -0.115 6.585 0.285 ;
        RECT  6.240 -0.115 6.515 0.115 ;
        RECT  6.120 -0.115 6.240 0.145 ;
        RECT  5.860 -0.115 6.120 0.115 ;
        RECT  5.740 -0.115 5.860 0.145 ;
        RECT  5.480 -0.115 5.740 0.115 ;
        RECT  5.360 -0.115 5.480 0.145 ;
        RECT  5.100 -0.115 5.360 0.115 ;
        RECT  4.980 -0.115 5.100 0.145 ;
        RECT  4.220 -0.115 4.980 0.115 ;
        RECT  4.100 -0.115 4.220 0.125 ;
        RECT  3.320 -0.115 4.100 0.115 ;
        RECT  3.200 -0.115 3.320 0.130 ;
        RECT  2.960 -0.115 3.200 0.115 ;
        RECT  2.840 -0.115 2.960 0.130 ;
        RECT  2.010 -0.115 2.840 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 1.145 7.000 1.375 ;
        RECT  6.870 0.685 6.950 1.375 ;
        RECT  6.585 1.145 6.870 1.375 ;
        RECT  6.515 0.975 6.585 1.375 ;
        RECT  6.250 1.145 6.515 1.375 ;
        RECT  6.130 1.010 6.250 1.375 ;
        RECT  5.890 1.145 6.130 1.375 ;
        RECT  5.770 1.010 5.890 1.375 ;
        RECT  5.520 1.145 5.770 1.375 ;
        RECT  5.400 1.130 5.520 1.375 ;
        RECT  5.120 1.145 5.400 1.375 ;
        RECT  5.000 1.130 5.120 1.375 ;
        RECT  4.280 1.145 5.000 1.375 ;
        RECT  4.160 1.015 4.280 1.375 ;
        RECT  3.320 1.145 4.160 1.375 ;
        RECT  3.200 1.130 3.320 1.375 ;
        RECT  2.100 1.145 3.200 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.695 0.185 6.765 0.465 ;
        RECT  6.695 0.765 6.765 1.065 ;
        RECT  6.685 0.355 6.695 0.465 ;
        RECT  6.685 0.765 6.695 0.905 ;
        RECT  5.985 0.710 6.070 0.800 ;
        RECT  5.985 0.355 6.050 0.455 ;
        RECT  5.550 0.355 5.635 0.455 ;
        RECT  5.590 0.710 5.635 0.800 ;
        RECT  6.210 0.545 6.320 0.615 ;
        RECT  6.140 0.215 6.210 0.940 ;
        RECT  4.870 0.215 6.140 0.285 ;
        RECT  5.650 0.870 6.140 0.940 ;
        RECT  5.580 0.870 5.650 1.060 ;
        RECT  5.440 0.545 5.620 0.615 ;
        RECT  4.450 0.990 5.580 1.060 ;
        RECT  5.370 0.370 5.440 0.815 ;
        RECT  5.010 0.370 5.370 0.440 ;
        RECT  5.220 0.695 5.370 0.815 ;
        RECT  5.150 0.545 5.290 0.615 ;
        RECT  5.080 0.545 5.150 0.920 ;
        RECT  4.590 0.850 5.080 0.920 ;
        RECT  4.940 0.370 5.010 0.630 ;
        RECT  4.910 0.530 4.940 0.630 ;
        RECT  4.800 0.215 4.870 0.430 ;
        RECT  4.730 0.685 4.830 0.755 ;
        RECT  4.660 0.195 4.730 0.755 ;
        RECT  4.540 0.195 4.660 0.265 ;
        RECT  4.520 0.345 4.590 0.920 ;
        RECT  4.420 0.185 4.540 0.265 ;
        RECT  4.380 0.345 4.450 0.790 ;
        RECT  4.380 0.870 4.450 1.060 ;
        RECT  4.000 0.195 4.420 0.265 ;
        RECT  4.140 0.345 4.380 0.415 ;
        RECT  3.900 0.870 4.380 0.940 ;
        RECT  4.240 0.510 4.310 0.780 ;
        RECT  3.770 0.710 4.240 0.780 ;
        RECT  4.070 0.345 4.140 0.630 ;
        RECT  3.930 0.195 4.000 0.615 ;
        RECT  3.850 0.545 3.930 0.615 ;
        RECT  3.830 0.870 3.900 1.060 ;
        RECT  3.790 0.260 3.860 0.440 ;
        RECT  2.290 0.990 3.830 1.060 ;
        RECT  3.770 0.370 3.790 0.440 ;
        RECT  3.700 0.370 3.770 0.780 ;
        RECT  2.385 0.200 3.710 0.270 ;
        RECT  2.390 0.850 3.700 0.920 ;
        RECT  3.535 0.350 3.605 0.780 ;
        RECT  3.410 0.350 3.535 0.420 ;
        RECT  3.400 0.680 3.535 0.780 ;
        RECT  3.325 0.540 3.380 0.610 ;
        RECT  3.255 0.355 3.325 0.780 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.710 3.255 0.780 ;
        RECT  2.835 0.345 2.905 0.780 ;
        RECT  2.470 0.345 2.835 0.415 ;
        RECT  2.610 0.710 2.835 0.780 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.200 2.385 0.420 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.060 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCND4BWP

MACRO SEDFKCNQD0BWP
    CLASS CORE ;
    FOREIGN SEDFKCNQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0280 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.490 1.540 0.610 ;
        RECT  1.435 0.490 1.505 0.765 ;
        END
    END SE
    PIN Q
        ANTENNAGATEAREA 0.0230 ;
        ANTENNADIFFAREA 0.0379 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.060 0.195 5.145 1.060 ;
        RECT  5.055 0.195 5.060 0.445 ;
        RECT  4.305 0.990 5.060 1.060 ;
        RECT  4.720 0.375 5.055 0.445 ;
        RECT  4.235 0.890 4.305 1.060 ;
        RECT  3.885 0.890 4.235 0.960 ;
        RECT  3.815 0.890 3.885 1.065 ;
        RECT  0.970 0.995 3.815 1.065 ;
        RECT  0.850 0.995 0.970 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0236 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 3.045 0.630 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.640 ;
        RECT  1.245 0.520 1.295 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 -0.115 5.180 0.115 ;
        RECT  4.865 -0.115 4.935 0.305 ;
        RECT  4.105 -0.115 4.865 0.115 ;
        RECT  4.035 -0.115 4.105 0.420 ;
        RECT  3.175 -0.115 4.035 0.115 ;
        RECT  3.055 -0.115 3.175 0.125 ;
        RECT  2.605 -0.115 3.055 0.115 ;
        RECT  2.485 -0.115 2.605 0.120 ;
        RECT  1.845 -0.115 2.485 0.115 ;
        RECT  1.775 -0.115 1.845 0.420 ;
        RECT  1.480 -0.115 1.775 0.115 ;
        RECT  1.360 -0.115 1.480 0.275 ;
        RECT  0.125 -0.115 1.360 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.960 1.145 5.180 1.375 ;
        RECT  4.840 1.140 4.960 1.375 ;
        RECT  4.120 1.145 4.840 1.375 ;
        RECT  3.995 1.030 4.120 1.375 ;
        RECT  3.175 1.145 3.995 1.375 ;
        RECT  3.055 1.135 3.175 1.375 ;
        RECT  2.605 1.145 3.055 1.375 ;
        RECT  2.485 1.135 2.605 1.375 ;
        RECT  1.840 1.145 2.485 1.375 ;
        RECT  1.720 1.135 1.840 1.375 ;
        RECT  1.480 1.145 1.720 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  1.120 1.145 1.360 1.375 ;
        RECT  1.000 1.135 1.120 1.375 ;
        RECT  0.330 1.145 1.000 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.920 0.520 4.990 0.910 ;
        RECT  4.605 0.520 4.920 0.590 ;
        RECT  4.390 0.840 4.920 0.910 ;
        RECT  4.465 0.690 4.670 0.760 ;
        RECT  4.535 0.200 4.605 0.590 ;
        RECT  4.440 0.200 4.535 0.270 ;
        RECT  4.395 0.350 4.465 0.760 ;
        RECT  4.250 0.205 4.320 0.820 ;
        RECT  4.240 0.205 4.250 0.325 ;
        RECT  4.020 0.750 4.250 0.820 ;
        RECT  4.110 0.520 4.180 0.640 ;
        RECT  3.715 0.520 4.110 0.590 ;
        RECT  3.900 0.680 4.020 0.820 ;
        RECT  3.705 0.300 3.715 0.590 ;
        RECT  3.635 0.300 3.705 0.920 ;
        RECT  2.205 0.195 3.550 0.265 ;
        RECT  2.110 0.855 3.550 0.925 ;
        RECT  3.345 0.335 3.415 0.785 ;
        RECT  3.260 0.335 3.345 0.435 ;
        RECT  3.260 0.680 3.345 0.785 ;
        RECT  3.185 0.540 3.250 0.610 ;
        RECT  3.115 0.355 3.185 0.785 ;
        RECT  2.870 0.355 3.115 0.425 ;
        RECT  2.870 0.715 3.115 0.785 ;
        RECT  2.475 0.345 2.790 0.415 ;
        RECT  2.475 0.715 2.790 0.785 ;
        RECT  2.405 0.345 2.475 0.785 ;
        RECT  2.230 0.505 2.300 0.760 ;
        RECT  1.680 0.505 2.230 0.575 ;
        RECT  2.135 0.195 2.205 0.420 ;
        RECT  1.970 0.675 2.130 0.745 ;
        RECT  1.900 0.675 1.970 0.925 ;
        RECT  1.175 0.855 1.900 0.925 ;
        RECT  1.610 0.190 1.680 0.780 ;
        RECT  1.595 0.190 1.610 0.310 ;
        RECT  1.580 0.680 1.610 0.780 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  1.105 0.335 1.175 0.925 ;
        RECT  0.790 0.335 1.105 0.405 ;
        RECT  0.590 0.855 1.105 0.925 ;
        RECT  0.870 0.505 0.990 0.775 ;
        RECT  0.385 0.705 0.870 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCNQD0BWP

MACRO SEDFKCNQD1BWP
    CLASS CORE ;
    FOREIGN SEDFKCNQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.615 0.195 5.705 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.470 -0.115 5.740 0.115 ;
        RECT  5.350 -0.115 5.470 0.145 ;
        RECT  5.080 -0.115 5.350 0.115 ;
        RECT  4.960 -0.115 5.080 0.145 ;
        RECT  4.225 -0.115 4.960 0.115 ;
        RECT  4.155 -0.115 4.225 0.420 ;
        RECT  3.315 -0.115 4.155 0.115 ;
        RECT  3.180 -0.115 3.315 0.125 ;
        RECT  2.980 -0.115 3.180 0.115 ;
        RECT  2.860 -0.115 2.980 0.125 ;
        RECT  2.010 -0.115 2.860 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.470 1.145 5.740 1.375 ;
        RECT  5.350 1.120 5.470 1.375 ;
        RECT  5.080 1.145 5.350 1.375 ;
        RECT  4.960 1.120 5.080 1.375 ;
        RECT  4.240 1.145 4.960 1.375 ;
        RECT  4.115 1.030 4.240 1.375 ;
        RECT  3.315 1.145 4.115 1.375 ;
        RECT  3.195 1.135 3.315 1.375 ;
        RECT  2.940 1.145 3.195 1.375 ;
        RECT  2.820 1.135 2.940 1.375 ;
        RECT  2.100 1.145 2.820 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.475 0.235 5.545 1.050 ;
        RECT  4.880 0.235 5.475 0.305 ;
        RECT  4.410 0.980 5.475 1.050 ;
        RECT  5.250 0.530 5.400 0.630 ;
        RECT  5.180 0.375 5.250 0.895 ;
        RECT  4.960 0.375 5.180 0.445 ;
        RECT  5.040 0.520 5.110 0.910 ;
        RECT  5.020 0.520 5.040 0.630 ;
        RECT  4.520 0.840 5.040 0.910 ;
        RECT  4.720 0.560 5.020 0.630 ;
        RECT  4.840 0.375 4.960 0.465 ;
        RECT  4.790 0.185 4.880 0.305 ;
        RECT  4.580 0.700 4.780 0.770 ;
        RECT  4.650 0.210 4.720 0.630 ;
        RECT  4.560 0.210 4.650 0.280 ;
        RECT  4.510 0.360 4.580 0.770 ;
        RECT  4.370 0.185 4.440 0.820 ;
        RECT  4.340 0.890 4.410 1.050 ;
        RECT  4.140 0.750 4.370 0.820 ;
        RECT  4.020 0.890 4.340 0.960 ;
        RECT  4.230 0.520 4.300 0.640 ;
        RECT  3.865 0.520 4.230 0.590 ;
        RECT  4.020 0.680 4.140 0.820 ;
        RECT  3.950 0.890 4.020 1.065 ;
        RECT  2.290 0.995 3.950 1.065 ;
        RECT  3.845 0.300 3.865 0.590 ;
        RECT  3.795 0.300 3.845 0.920 ;
        RECT  3.775 0.520 3.795 0.920 ;
        RECT  2.385 0.195 3.690 0.265 ;
        RECT  2.390 0.855 3.690 0.925 ;
        RECT  3.575 0.335 3.645 0.785 ;
        RECT  3.400 0.335 3.575 0.435 ;
        RECT  3.400 0.685 3.575 0.785 ;
        RECT  3.325 0.545 3.390 0.615 ;
        RECT  3.255 0.355 3.325 0.785 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.715 3.255 0.785 ;
        RECT  2.835 0.335 2.905 0.785 ;
        RECT  2.470 0.335 2.835 0.405 ;
        RECT  2.610 0.715 2.835 0.785 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.195 2.385 0.410 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.065 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCNQD1BWP

MACRO SEDFKCNQD2BWP
    CLASS CORE ;
    FOREIGN SEDFKCNQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0120 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.645 0.355 5.705 0.815 ;
        RECT  5.635 0.185 5.645 1.035 ;
        RECT  5.575 0.185 5.635 0.465 ;
        RECT  5.575 0.745 5.635 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 -0.115 5.880 0.115 ;
        RECT  5.750 -0.115 5.830 0.300 ;
        RECT  5.470 -0.115 5.750 0.115 ;
        RECT  5.350 -0.115 5.470 0.140 ;
        RECT  5.080 -0.115 5.350 0.115 ;
        RECT  4.960 -0.115 5.080 0.145 ;
        RECT  4.225 -0.115 4.960 0.115 ;
        RECT  4.155 -0.115 4.225 0.420 ;
        RECT  3.315 -0.115 4.155 0.115 ;
        RECT  3.195 -0.115 3.315 0.125 ;
        RECT  2.980 -0.115 3.195 0.115 ;
        RECT  2.860 -0.115 2.980 0.125 ;
        RECT  2.010 -0.115 2.860 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.145 5.880 1.375 ;
        RECT  5.750 0.905 5.830 1.375 ;
        RECT  5.470 1.145 5.750 1.375 ;
        RECT  5.350 1.120 5.470 1.375 ;
        RECT  5.080 1.145 5.350 1.375 ;
        RECT  4.960 1.120 5.080 1.375 ;
        RECT  4.240 1.145 4.960 1.375 ;
        RECT  4.115 1.030 4.240 1.375 ;
        RECT  3.315 1.145 4.115 1.375 ;
        RECT  3.195 1.135 3.315 1.375 ;
        RECT  2.940 1.145 3.195 1.375 ;
        RECT  2.820 1.135 2.940 1.375 ;
        RECT  2.100 1.145 2.820 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.235 5.495 1.050 ;
        RECT  4.880 0.235 5.425 0.305 ;
        RECT  4.410 0.980 5.425 1.050 ;
        RECT  5.285 0.385 5.355 0.875 ;
        RECT  4.840 0.385 5.285 0.455 ;
        RECT  5.150 0.805 5.285 0.875 ;
        RECT  4.940 0.545 5.160 0.615 ;
        RECT  4.870 0.545 4.940 0.910 ;
        RECT  4.790 0.185 4.880 0.305 ;
        RECT  4.720 0.545 4.870 0.615 ;
        RECT  4.520 0.840 4.870 0.910 ;
        RECT  4.580 0.700 4.780 0.770 ;
        RECT  4.650 0.210 4.720 0.615 ;
        RECT  4.560 0.210 4.650 0.280 ;
        RECT  4.510 0.360 4.580 0.770 ;
        RECT  4.370 0.185 4.440 0.820 ;
        RECT  4.340 0.890 4.410 1.050 ;
        RECT  4.140 0.750 4.370 0.820 ;
        RECT  4.020 0.890 4.340 0.960 ;
        RECT  4.220 0.520 4.300 0.640 ;
        RECT  3.865 0.520 4.220 0.590 ;
        RECT  4.020 0.680 4.140 0.820 ;
        RECT  3.950 0.890 4.020 1.065 ;
        RECT  2.290 0.995 3.950 1.065 ;
        RECT  3.845 0.300 3.865 0.590 ;
        RECT  3.795 0.300 3.845 0.920 ;
        RECT  3.775 0.520 3.795 0.920 ;
        RECT  2.385 0.195 3.690 0.265 ;
        RECT  2.390 0.855 3.690 0.925 ;
        RECT  3.575 0.335 3.645 0.785 ;
        RECT  3.400 0.335 3.575 0.435 ;
        RECT  3.400 0.685 3.575 0.785 ;
        RECT  3.325 0.545 3.390 0.615 ;
        RECT  3.255 0.355 3.325 0.785 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.715 3.255 0.785 ;
        RECT  2.835 0.335 2.905 0.785 ;
        RECT  2.470 0.335 2.835 0.405 ;
        RECT  2.610 0.715 2.835 0.785 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.195 2.385 0.410 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.065 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCNQD2BWP

MACRO SEDFKCNQD4BWP
    CLASS CORE ;
    FOREIGN SEDFKCNQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.630 2.205 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.995 0.185 6.065 0.465 ;
        RECT  5.995 0.765 6.065 1.065 ;
        RECT  5.915 0.355 5.995 0.465 ;
        RECT  5.915 0.765 5.995 0.905 ;
        RECT  5.705 0.355 5.915 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.765 5.705 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0264 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0224 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.495 3.185 0.640 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.310 0.640 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.465 ;
        RECT  5.910 -0.115 6.170 0.115 ;
        RECT  5.790 -0.115 5.910 0.275 ;
        RECT  5.540 -0.115 5.790 0.115 ;
        RECT  5.420 -0.115 5.540 0.145 ;
        RECT  5.160 -0.115 5.420 0.115 ;
        RECT  5.040 -0.115 5.160 0.145 ;
        RECT  4.235 -0.115 5.040 0.115 ;
        RECT  4.165 -0.115 4.235 0.420 ;
        RECT  3.320 -0.115 4.165 0.115 ;
        RECT  3.200 -0.115 3.320 0.130 ;
        RECT  2.960 -0.115 3.200 0.115 ;
        RECT  2.840 -0.115 2.960 0.130 ;
        RECT  2.010 -0.115 2.840 0.115 ;
        RECT  1.890 -0.115 2.010 0.420 ;
        RECT  1.470 -0.115 1.890 0.115 ;
        RECT  1.350 -0.115 1.470 0.260 ;
        RECT  0.125 -0.115 1.350 0.115 ;
        RECT  0.055 -0.115 0.125 0.340 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.675 6.250 1.375 ;
        RECT  5.885 1.145 6.170 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  5.540 1.145 5.815 1.375 ;
        RECT  5.420 1.120 5.540 1.375 ;
        RECT  5.140 1.145 5.420 1.375 ;
        RECT  5.010 1.120 5.140 1.375 ;
        RECT  4.280 1.145 5.010 1.375 ;
        RECT  4.155 1.030 4.280 1.375 ;
        RECT  3.320 1.145 4.155 1.375 ;
        RECT  3.200 1.130 3.320 1.375 ;
        RECT  2.925 1.145 3.200 1.375 ;
        RECT  2.805 1.135 2.925 1.375 ;
        RECT  2.100 1.145 2.805 1.375 ;
        RECT  2.030 1.010 2.100 1.375 ;
        RECT  1.460 1.145 2.030 1.375 ;
        RECT  1.340 1.130 1.460 1.375 ;
        RECT  1.110 1.145 1.340 1.375 ;
        RECT  0.990 1.135 1.110 1.375 ;
        RECT  0.330 1.145 0.990 1.375 ;
        RECT  0.210 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.995 0.185 6.065 0.465 ;
        RECT  5.995 0.765 6.065 1.065 ;
        RECT  5.985 0.355 5.995 0.465 ;
        RECT  5.985 0.765 5.995 0.905 ;
        RECT  5.555 0.515 5.580 0.640 ;
        RECT  5.485 0.220 5.555 1.000 ;
        RECT  4.880 0.220 5.485 0.290 ;
        RECT  5.230 0.930 5.485 1.000 ;
        RECT  5.345 0.390 5.415 0.850 ;
        RECT  4.810 0.390 5.345 0.460 ;
        RECT  5.140 0.780 5.345 0.850 ;
        RECT  4.990 0.545 5.265 0.615 ;
        RECT  5.070 0.780 5.140 1.050 ;
        RECT  4.440 0.980 5.070 1.050 ;
        RECT  4.920 0.545 4.990 0.910 ;
        RECT  4.740 0.545 4.920 0.615 ;
        RECT  4.570 0.840 4.920 0.910 ;
        RECT  4.600 0.700 4.840 0.770 ;
        RECT  4.670 0.200 4.740 0.615 ;
        RECT  4.570 0.200 4.670 0.270 ;
        RECT  4.530 0.350 4.600 0.770 ;
        RECT  4.390 0.205 4.460 0.820 ;
        RECT  4.370 0.890 4.440 1.050 ;
        RECT  4.140 0.750 4.390 0.820 ;
        RECT  4.040 0.890 4.370 0.960 ;
        RECT  4.245 0.520 4.315 0.640 ;
        RECT  3.865 0.520 4.245 0.590 ;
        RECT  4.020 0.680 4.140 0.820 ;
        RECT  3.970 0.890 4.040 1.060 ;
        RECT  2.290 0.990 3.970 1.060 ;
        RECT  3.845 0.300 3.865 0.590 ;
        RECT  3.795 0.300 3.845 0.920 ;
        RECT  3.775 0.520 3.795 0.920 ;
        RECT  2.385 0.200 3.690 0.270 ;
        RECT  2.390 0.850 3.690 0.920 ;
        RECT  3.575 0.355 3.645 0.780 ;
        RECT  3.400 0.355 3.575 0.455 ;
        RECT  3.400 0.680 3.575 0.780 ;
        RECT  3.325 0.540 3.380 0.610 ;
        RECT  3.255 0.355 3.325 0.780 ;
        RECT  3.010 0.355 3.255 0.425 ;
        RECT  3.010 0.710 3.255 0.780 ;
        RECT  2.835 0.345 2.905 0.780 ;
        RECT  2.470 0.345 2.835 0.415 ;
        RECT  2.610 0.710 2.835 0.780 ;
        RECT  2.345 0.490 2.415 0.760 ;
        RECT  2.315 0.200 2.385 0.420 ;
        RECT  1.805 0.490 2.345 0.560 ;
        RECT  2.220 0.855 2.290 1.060 ;
        RECT  1.960 0.855 2.220 0.925 ;
        RECT  1.890 0.855 1.960 1.060 ;
        RECT  0.960 0.990 1.890 1.060 ;
        RECT  1.735 0.330 1.805 0.910 ;
        RECT  1.640 0.185 1.760 0.255 ;
        RECT  1.570 0.185 1.640 0.910 ;
        RECT  1.555 0.330 1.570 0.450 ;
        RECT  1.555 0.790 1.570 0.910 ;
        RECT  1.460 0.520 1.500 0.640 ;
        RECT  1.390 0.335 1.460 0.915 ;
        RECT  0.790 0.335 1.390 0.405 ;
        RECT  0.590 0.845 1.390 0.915 ;
        RECT  0.390 0.195 1.270 0.265 ;
        RECT  0.860 0.505 0.980 0.775 ;
        RECT  0.840 0.990 0.960 1.070 ;
        RECT  0.385 0.705 0.860 0.775 ;
        RECT  0.315 0.340 0.385 0.915 ;
        RECT  0.305 0.340 0.315 0.410 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.235 0.220 0.305 0.410 ;
        RECT  0.055 0.845 0.125 1.050 ;
    END
END SEDFKCNQD4BWP

MACRO SEDFQD0BWP
    CLASS CORE ;
    FOREIGN SEDFQD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0276 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.915 0.350 5.005 0.905 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 -0.115 5.040 0.115 ;
        RECT  4.740 -0.115 4.810 0.480 ;
        RECT  4.415 -0.115 4.740 0.115 ;
        RECT  4.345 -0.115 4.415 0.270 ;
        RECT  1.420 -0.115 4.345 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.740 0.760 4.810 1.375 ;
        RECT  3.680 1.145 4.740 1.375 ;
        RECT  3.560 1.020 3.680 1.375 ;
        RECT  0.330 1.145 3.560 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.600 0.350 4.670 1.060 ;
        RECT  4.335 0.350 4.600 0.420 ;
        RECT  3.860 0.990 4.600 1.060 ;
        RECT  4.460 0.520 4.530 0.920 ;
        RECT  4.010 0.850 4.460 0.920 ;
        RECT  4.265 0.350 4.335 0.600 ;
        RECT  4.160 0.685 4.240 0.755 ;
        RECT  4.090 0.195 4.160 0.755 ;
        RECT  3.975 0.195 4.090 0.265 ;
        RECT  3.940 0.340 4.010 0.920 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.855 0.410 3.870 0.810 ;
        RECT  3.790 0.880 3.860 1.060 ;
        RECT  3.800 0.335 3.855 0.810 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.800 0.455 ;
        RECT  3.535 0.740 3.800 0.810 ;
        RECT  3.435 0.880 3.790 0.950 ;
        RECT  3.675 0.530 3.720 0.650 ;
        RECT  3.605 0.340 3.675 0.650 ;
        RECT  3.285 0.340 3.605 0.410 ;
        RECT  3.465 0.520 3.535 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.640 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.570 0.675 0.640 ;
        RECT  0.345 0.570 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQD0BWP

MACRO SEDFQD1BWP
    CLASS CORE ;
    FOREIGN SEDFQD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0302 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.915 0.195 5.005 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 -0.115 5.040 0.115 ;
        RECT  4.740 -0.115 4.810 0.475 ;
        RECT  4.415 -0.115 4.740 0.115 ;
        RECT  4.345 -0.115 4.415 0.270 ;
        RECT  1.420 -0.115 4.345 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.740 0.680 4.810 1.375 ;
        RECT  3.680 1.145 4.740 1.375 ;
        RECT  3.560 1.020 3.680 1.375 ;
        RECT  0.330 1.145 3.560 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.600 0.350 4.670 1.060 ;
        RECT  4.335 0.350 4.600 0.420 ;
        RECT  3.860 0.990 4.600 1.060 ;
        RECT  4.460 0.520 4.530 0.920 ;
        RECT  4.010 0.850 4.460 0.920 ;
        RECT  4.265 0.350 4.335 0.590 ;
        RECT  4.160 0.685 4.240 0.755 ;
        RECT  4.090 0.195 4.160 0.755 ;
        RECT  3.975 0.195 4.090 0.265 ;
        RECT  3.940 0.340 4.010 0.920 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.850 0.410 3.870 0.810 ;
        RECT  3.790 0.880 3.860 1.060 ;
        RECT  3.800 0.335 3.850 0.810 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.800 0.460 ;
        RECT  3.535 0.740 3.800 0.810 ;
        RECT  3.435 0.880 3.790 0.950 ;
        RECT  3.675 0.520 3.720 0.640 ;
        RECT  3.605 0.340 3.675 0.640 ;
        RECT  3.285 0.340 3.605 0.410 ;
        RECT  3.465 0.520 3.535 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.545 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.545 1.765 0.615 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQD1BWP

MACRO SEDFQD2BWP
    CLASS CORE ;
    FOREIGN SEDFQD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0302 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.355 5.145 0.820 ;
        RECT  5.075 0.185 5.085 1.035 ;
        RECT  5.015 0.185 5.075 0.465 ;
        RECT  5.015 0.735 5.075 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.300 ;
        RECT  4.930 -0.115 5.190 0.115 ;
        RECT  4.810 -0.115 4.930 0.280 ;
        RECT  4.455 -0.115 4.810 0.115 ;
        RECT  4.385 -0.115 4.455 0.280 ;
        RECT  1.420 -0.115 4.385 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.905 5.270 1.375 ;
        RECT  4.930 1.145 5.190 1.375 ;
        RECT  4.810 1.010 4.930 1.375 ;
        RECT  3.700 1.145 4.810 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  0.330 1.145 3.580 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.365 4.935 0.910 ;
        RECT  4.355 0.365 4.865 0.435 ;
        RECT  4.645 0.840 4.865 0.910 ;
        RECT  4.505 0.545 4.775 0.615 ;
        RECT  4.575 0.840 4.645 1.050 ;
        RECT  3.880 0.980 4.575 1.050 ;
        RECT  4.435 0.545 4.505 0.910 ;
        RECT  4.030 0.840 4.435 0.910 ;
        RECT  4.285 0.365 4.355 0.620 ;
        RECT  4.180 0.700 4.240 0.770 ;
        RECT  4.110 0.195 4.180 0.770 ;
        RECT  3.975 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.910 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.050 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.820 0.455 ;
        RECT  3.550 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.690 0.525 3.740 0.645 ;
        RECT  3.620 0.340 3.690 0.645 ;
        RECT  3.285 0.340 3.620 0.410 ;
        RECT  3.480 0.520 3.550 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.545 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.545 1.765 0.615 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQD2BWP

MACRO SEDFQD4BWP
    CLASS CORE ;
    FOREIGN SEDFQD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0302 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.715 0.185 5.785 0.465 ;
        RECT  5.715 0.765 5.785 1.065 ;
        RECT  5.635 0.355 5.715 0.465 ;
        RECT  5.635 0.765 5.715 0.905 ;
        RECT  5.425 0.355 5.635 0.905 ;
        RECT  5.355 0.185 5.425 0.465 ;
        RECT  5.355 0.765 5.425 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 -0.115 6.020 0.115 ;
        RECT  5.890 -0.115 5.970 0.465 ;
        RECT  5.630 -0.115 5.890 0.115 ;
        RECT  5.510 -0.115 5.630 0.275 ;
        RECT  5.270 -0.115 5.510 0.115 ;
        RECT  5.150 -0.115 5.270 0.280 ;
        RECT  4.835 -0.115 5.150 0.115 ;
        RECT  4.765 -0.115 4.835 0.290 ;
        RECT  1.420 -0.115 4.765 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.970 1.145 6.020 1.375 ;
        RECT  5.890 0.685 5.970 1.375 ;
        RECT  5.605 1.145 5.890 1.375 ;
        RECT  5.535 0.975 5.605 1.375 ;
        RECT  5.270 1.145 5.535 1.375 ;
        RECT  5.150 1.005 5.270 1.375 ;
        RECT  4.090 1.145 5.150 1.375 ;
        RECT  3.970 1.040 4.090 1.375 ;
        RECT  3.700 1.145 3.970 1.375 ;
        RECT  3.580 1.040 3.700 1.375 ;
        RECT  0.330 1.145 3.580 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.715 0.185 5.785 0.465 ;
        RECT  5.715 0.765 5.785 1.065 ;
        RECT  5.705 0.355 5.715 0.465 ;
        RECT  5.705 0.765 5.715 0.905 ;
        RECT  5.205 0.365 5.275 0.935 ;
        RECT  4.775 0.365 5.205 0.435 ;
        RECT  5.045 0.865 5.205 0.935 ;
        RECT  4.975 0.520 5.045 0.790 ;
        RECT  4.975 0.865 5.045 1.050 ;
        RECT  4.810 0.720 4.975 0.790 ;
        RECT  4.255 0.980 4.975 1.050 ;
        RECT  4.740 0.720 4.810 0.910 ;
        RECT  4.705 0.365 4.775 0.640 ;
        RECT  4.410 0.840 4.740 0.910 ;
        RECT  4.550 0.700 4.620 0.770 ;
        RECT  4.480 0.200 4.550 0.770 ;
        RECT  4.350 0.200 4.480 0.270 ;
        RECT  4.340 0.340 4.410 0.910 ;
        RECT  4.210 0.185 4.350 0.270 ;
        RECT  4.310 0.340 4.340 0.460 ;
        RECT  4.230 0.750 4.270 0.820 ;
        RECT  4.185 0.900 4.255 1.050 ;
        RECT  4.160 0.350 4.230 0.820 ;
        RECT  3.295 0.200 4.210 0.270 ;
        RECT  3.435 0.900 4.185 0.970 ;
        RECT  3.750 0.350 4.160 0.420 ;
        RECT  3.580 0.750 4.160 0.820 ;
        RECT  3.285 0.540 3.950 0.610 ;
        RECT  3.460 0.680 3.580 0.820 ;
        RECT  3.365 0.900 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.200 3.110 0.270 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.200 1.775 0.460 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.690 1.680 0.760 ;
        RECT  1.460 0.690 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQD4BWP

MACRO SEDFQND0BWP
    CLASS CORE ;
    FOREIGN SEDFQND0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0272 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.320 5.005 0.905 ;
        RECT  4.915 0.320 4.935 0.440 ;
        RECT  4.915 0.765 4.935 0.905 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0260 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 -0.115 5.040 0.115 ;
        RECT  4.740 -0.115 4.810 0.440 ;
        RECT  4.415 -0.115 4.740 0.115 ;
        RECT  4.345 -0.115 4.415 0.270 ;
        RECT  1.420 -0.115 4.345 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.740 0.760 4.810 1.375 ;
        RECT  3.680 1.145 4.740 1.375 ;
        RECT  3.560 1.020 3.680 1.375 ;
        RECT  0.330 1.145 3.560 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.670 0.520 4.865 0.640 ;
        RECT  4.600 0.350 4.670 1.060 ;
        RECT  4.335 0.350 4.600 0.420 ;
        RECT  3.860 0.990 4.600 1.060 ;
        RECT  4.460 0.520 4.530 0.920 ;
        RECT  4.010 0.850 4.460 0.920 ;
        RECT  4.265 0.350 4.335 0.590 ;
        RECT  4.160 0.685 4.240 0.755 ;
        RECT  4.090 0.195 4.160 0.755 ;
        RECT  3.975 0.195 4.090 0.265 ;
        RECT  3.940 0.345 4.010 0.920 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.800 0.335 3.870 0.810 ;
        RECT  3.790 0.880 3.860 1.060 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.800 0.455 ;
        RECT  3.535 0.740 3.800 0.810 ;
        RECT  3.435 0.880 3.790 0.950 ;
        RECT  3.675 0.520 3.730 0.640 ;
        RECT  3.605 0.340 3.675 0.640 ;
        RECT  3.285 0.340 3.605 0.410 ;
        RECT  3.465 0.520 3.535 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.540 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.540 1.765 0.610 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.640 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.570 0.675 0.640 ;
        RECT  0.345 0.570 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQND0BWP

MACRO SEDFQND1BWP
    CLASS CORE ;
    FOREIGN SEDFQND1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.045 ;
        RECT  4.915 0.185 4.935 0.465 ;
        RECT  4.915 0.745 4.935 1.045 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 -0.115 5.040 0.115 ;
        RECT  4.740 -0.115 4.810 0.465 ;
        RECT  4.415 -0.115 4.740 0.115 ;
        RECT  4.345 -0.115 4.415 0.270 ;
        RECT  1.420 -0.115 4.345 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.740 0.740 4.810 1.375 ;
        RECT  3.680 1.145 4.740 1.375 ;
        RECT  3.560 1.020 3.680 1.375 ;
        RECT  0.330 1.145 3.560 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.670 0.545 4.865 0.615 ;
        RECT  4.600 0.350 4.670 1.060 ;
        RECT  4.335 0.350 4.600 0.420 ;
        RECT  3.860 0.990 4.600 1.060 ;
        RECT  4.460 0.520 4.530 0.920 ;
        RECT  4.010 0.850 4.460 0.920 ;
        RECT  4.265 0.350 4.335 0.590 ;
        RECT  4.160 0.685 4.240 0.755 ;
        RECT  4.090 0.195 4.160 0.755 ;
        RECT  3.975 0.195 4.090 0.265 ;
        RECT  3.940 0.350 4.010 0.920 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.800 0.335 3.870 0.810 ;
        RECT  3.790 0.880 3.860 1.060 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.800 0.455 ;
        RECT  3.535 0.740 3.800 0.810 ;
        RECT  3.435 0.880 3.790 0.950 ;
        RECT  3.675 0.520 3.730 0.640 ;
        RECT  3.605 0.340 3.675 0.640 ;
        RECT  3.285 0.340 3.605 0.410 ;
        RECT  3.465 0.520 3.535 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.545 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.545 1.765 0.615 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQND1BWP

MACRO SEDFQND2BWP
    CLASS CORE ;
    FOREIGN SEDFQND2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.355 5.145 0.820 ;
        RECT  5.075 0.185 5.085 1.035 ;
        RECT  5.015 0.185 5.075 0.465 ;
        RECT  5.015 0.735 5.075 1.035 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.300 ;
        RECT  4.930 -0.115 5.190 0.115 ;
        RECT  4.810 -0.115 4.930 0.280 ;
        RECT  4.455 -0.115 4.810 0.115 ;
        RECT  4.385 -0.115 4.455 0.280 ;
        RECT  1.420 -0.115 4.385 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.905 5.270 1.375 ;
        RECT  4.930 1.145 5.190 1.375 ;
        RECT  4.810 1.005 4.930 1.375 ;
        RECT  3.700 1.145 4.810 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  0.330 1.145 3.580 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.855 0.365 4.925 0.910 ;
        RECT  4.355 0.365 4.855 0.435 ;
        RECT  4.645 0.840 4.855 0.910 ;
        RECT  4.575 0.840 4.645 1.050 ;
        RECT  3.880 0.980 4.575 1.050 ;
        RECT  4.505 0.545 4.570 0.615 ;
        RECT  4.435 0.545 4.505 0.910 ;
        RECT  4.030 0.840 4.435 0.910 ;
        RECT  4.285 0.365 4.355 0.620 ;
        RECT  4.180 0.700 4.240 0.770 ;
        RECT  4.110 0.195 4.180 0.770 ;
        RECT  3.975 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.910 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.050 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.820 0.455 ;
        RECT  3.550 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.690 0.520 3.730 0.640 ;
        RECT  3.620 0.340 3.690 0.640 ;
        RECT  3.285 0.340 3.620 0.410 ;
        RECT  3.480 0.520 3.550 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.195 3.110 0.265 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.535 1.835 0.780 ;
        RECT  1.705 0.195 1.775 0.455 ;
        RECT  1.390 0.535 1.765 0.605 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQND2BWP

MACRO SEDFQND4BWP
    CLASS CORE ;
    FOREIGN SEDFQND4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.190 0.630 ;
        RECT  1.990 0.495 2.065 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0298 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.225 0.630 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.295 0.185 5.365 0.465 ;
        RECT  5.295 0.755 5.365 1.065 ;
        RECT  5.215 0.355 5.295 0.465 ;
        RECT  5.215 0.755 5.295 0.905 ;
        RECT  5.005 0.355 5.215 0.905 ;
        RECT  4.935 0.185 5.005 0.465 ;
        RECT  4.935 0.755 5.005 1.065 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0316 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.350 0.245 0.670 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0172 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.385 0.570 0.485 ;
        RECT  0.455 0.215 0.525 0.485 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.625 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.550 0.465 ;
        RECT  5.210 -0.115 5.470 0.115 ;
        RECT  5.090 -0.115 5.210 0.275 ;
        RECT  4.850 -0.115 5.090 0.115 ;
        RECT  4.730 -0.115 4.850 0.285 ;
        RECT  4.490 -0.115 4.730 0.115 ;
        RECT  4.370 -0.115 4.490 0.285 ;
        RECT  1.420 -0.115 4.370 0.115 ;
        RECT  1.300 -0.115 1.420 0.275 ;
        RECT  0.330 -0.115 1.300 0.115 ;
        RECT  0.210 -0.115 0.330 0.260 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 1.145 5.600 1.375 ;
        RECT  5.470 0.680 5.550 1.375 ;
        RECT  5.185 1.145 5.470 1.375 ;
        RECT  5.115 0.985 5.185 1.375 ;
        RECT  4.850 1.145 5.115 1.375 ;
        RECT  4.730 1.005 4.850 1.375 ;
        RECT  3.700 1.145 4.730 1.375 ;
        RECT  3.580 1.020 3.700 1.375 ;
        RECT  0.330 1.145 3.580 1.375 ;
        RECT  0.210 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.295 0.185 5.365 0.465 ;
        RECT  5.295 0.755 5.365 1.065 ;
        RECT  5.285 0.355 5.295 0.465 ;
        RECT  5.285 0.755 5.295 0.905 ;
        RECT  4.855 0.520 4.890 0.640 ;
        RECT  4.785 0.370 4.855 0.930 ;
        RECT  4.645 0.370 4.785 0.440 ;
        RECT  4.645 0.860 4.785 0.930 ;
        RECT  4.575 0.185 4.645 0.440 ;
        RECT  4.575 0.860 4.645 1.050 ;
        RECT  4.535 0.520 4.605 0.790 ;
        RECT  4.345 0.370 4.575 0.440 ;
        RECT  3.880 0.980 4.575 1.050 ;
        RECT  4.410 0.720 4.535 0.790 ;
        RECT  4.340 0.720 4.410 0.910 ;
        RECT  4.275 0.370 4.345 0.610 ;
        RECT  4.030 0.840 4.340 0.910 ;
        RECT  4.180 0.700 4.240 0.770 ;
        RECT  4.110 0.195 4.180 0.770 ;
        RECT  3.975 0.195 4.110 0.265 ;
        RECT  3.960 0.350 4.030 0.910 ;
        RECT  3.835 0.185 3.975 0.265 ;
        RECT  3.820 0.335 3.890 0.810 ;
        RECT  3.810 0.880 3.880 1.050 ;
        RECT  3.295 0.195 3.835 0.265 ;
        RECT  3.760 0.335 3.820 0.455 ;
        RECT  3.550 0.740 3.820 0.810 ;
        RECT  3.435 0.880 3.810 0.950 ;
        RECT  3.690 0.520 3.730 0.640 ;
        RECT  3.620 0.340 3.690 0.640 ;
        RECT  3.285 0.340 3.620 0.410 ;
        RECT  3.480 0.520 3.550 0.810 ;
        RECT  3.365 0.880 3.435 1.065 ;
        RECT  0.940 0.995 3.365 1.065 ;
        RECT  3.215 0.340 3.285 0.910 ;
        RECT  1.670 0.855 3.130 0.925 ;
        RECT  1.775 0.200 3.110 0.270 ;
        RECT  3.005 0.340 3.075 0.785 ;
        RECT  2.835 0.340 3.005 0.460 ;
        RECT  2.840 0.685 3.005 0.785 ;
        RECT  2.765 0.545 2.830 0.615 ;
        RECT  2.695 0.345 2.765 0.785 ;
        RECT  2.430 0.345 2.695 0.415 ;
        RECT  2.410 0.695 2.695 0.785 ;
        RECT  2.270 0.355 2.340 0.785 ;
        RECT  1.940 0.355 2.270 0.425 ;
        RECT  2.240 0.685 2.270 0.785 ;
        RECT  1.765 0.540 1.835 0.780 ;
        RECT  1.705 0.200 1.775 0.460 ;
        RECT  1.390 0.540 1.765 0.610 ;
        RECT  1.530 0.695 1.680 0.765 ;
        RECT  1.460 0.695 1.530 0.925 ;
        RECT  0.900 0.855 1.460 0.925 ;
        RECT  1.320 0.345 1.390 0.785 ;
        RECT  1.110 0.345 1.320 0.415 ;
        RECT  1.110 0.715 1.320 0.785 ;
        RECT  0.820 0.995 0.940 1.075 ;
        RECT  0.830 0.235 0.900 0.925 ;
        RECT  0.685 0.235 0.830 0.305 ;
        RECT  0.570 0.805 0.830 0.875 ;
        RECT  0.675 0.390 0.745 0.630 ;
        RECT  0.595 0.185 0.685 0.305 ;
        RECT  0.415 0.560 0.675 0.630 ;
        RECT  0.345 0.560 0.415 0.820 ;
        RECT  0.125 0.750 0.345 0.820 ;
        RECT  0.105 0.185 0.140 0.285 ;
        RECT  0.105 0.750 0.125 0.950 ;
        RECT  0.055 0.185 0.105 0.950 ;
        RECT  0.035 0.185 0.055 0.820 ;
    END
END SEDFQND4BWP

MACRO SEDFQNXD0BWP
    CLASS CORE ;
    FOREIGN SEDFQNXD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0246 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 0.215 5.565 1.045 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0362 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.360 -0.115 5.600 0.115 ;
        RECT  5.240 -0.115 5.360 0.125 ;
        RECT  5.060 -0.115 5.240 0.115 ;
        RECT  4.940 -0.115 5.060 0.125 ;
        RECT  4.160 -0.115 4.940 0.115 ;
        RECT  4.040 -0.115 4.160 0.125 ;
        RECT  3.430 -0.115 4.040 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  3.080 -0.115 3.360 0.115 ;
        RECT  2.960 -0.115 3.080 0.140 ;
        RECT  2.455 -0.115 2.960 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.360 1.145 5.600 1.375 ;
        RECT  5.240 1.135 5.360 1.375 ;
        RECT  5.060 1.145 5.240 1.375 ;
        RECT  4.940 1.135 5.060 1.375 ;
        RECT  4.160 1.145 4.940 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  3.080 1.145 3.640 1.375 ;
        RECT  2.960 1.140 3.080 1.375 ;
        RECT  2.700 1.145 2.960 1.375 ;
        RECT  2.580 1.135 2.700 1.375 ;
        RECT  2.320 1.145 2.580 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.480 1.145 0.735 1.375 ;
        RECT  0.360 1.140 0.480 1.375 ;
        RECT  0.125 1.145 0.360 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.340 0.195 5.410 1.065 ;
        RECT  4.820 0.195 5.340 0.265 ;
        RECT  4.360 0.995 5.340 1.065 ;
        RECT  5.200 0.345 5.270 0.925 ;
        RECT  4.960 0.345 5.200 0.415 ;
        RECT  5.100 0.825 5.200 0.925 ;
        RECT  5.030 0.520 5.100 0.755 ;
        RECT  4.960 0.685 5.030 0.925 ;
        RECT  4.890 0.345 4.960 0.615 ;
        RECT  4.520 0.855 4.960 0.925 ;
        RECT  4.820 0.545 4.890 0.615 ;
        RECT  4.750 0.195 4.820 0.440 ;
        RECT  4.680 0.715 4.760 0.785 ;
        RECT  4.610 0.195 4.680 0.785 ;
        RECT  4.480 0.195 4.610 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.730 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.635 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.465 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.355 0.335 2.465 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.355 0.405 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.255 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.145 0.195 1.255 0.410 ;
        RECT  0.820 0.340 1.145 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.670 0.500 0.675 0.910 ;
        RECT  0.605 0.340 0.670 0.910 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.605 0.590 ;
        RECT  0.485 0.500 0.590 0.590 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.405 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.215 0.835 0.330 0.935 ;
        RECT  0.190 0.195 0.260 0.630 ;
        RECT  0.100 0.530 0.190 0.630 ;
    END
END SEDFQNXD0BWP

MACRO SEDFQNXD1BWP
    CLASS CORE ;
    FOREIGN SEDFQNXD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.070 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.360 -0.115 5.600 0.115 ;
        RECT  5.240 -0.115 5.360 0.125 ;
        RECT  5.060 -0.115 5.240 0.115 ;
        RECT  4.940 -0.115 5.060 0.125 ;
        RECT  4.160 -0.115 4.940 0.115 ;
        RECT  4.040 -0.115 4.160 0.125 ;
        RECT  3.430 -0.115 4.040 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  3.080 -0.115 3.360 0.115 ;
        RECT  2.960 -0.115 3.080 0.140 ;
        RECT  2.455 -0.115 2.960 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.360 1.145 5.600 1.375 ;
        RECT  5.240 1.135 5.360 1.375 ;
        RECT  5.060 1.145 5.240 1.375 ;
        RECT  4.940 1.135 5.060 1.375 ;
        RECT  4.160 1.145 4.940 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  3.080 1.145 3.640 1.375 ;
        RECT  2.960 1.140 3.080 1.375 ;
        RECT  2.700 1.145 2.960 1.375 ;
        RECT  2.580 1.135 2.700 1.375 ;
        RECT  2.320 1.145 2.580 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.480 1.145 0.735 1.375 ;
        RECT  0.360 1.140 0.480 1.375 ;
        RECT  0.125 1.145 0.360 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.335 0.195 5.405 1.065 ;
        RECT  4.800 0.195 5.335 0.265 ;
        RECT  4.360 0.995 5.335 1.065 ;
        RECT  5.195 0.360 5.265 0.925 ;
        RECT  4.940 0.360 5.195 0.430 ;
        RECT  5.100 0.825 5.195 0.925 ;
        RECT  5.030 0.520 5.080 0.755 ;
        RECT  5.010 0.520 5.030 0.925 ;
        RECT  4.960 0.685 5.010 0.925 ;
        RECT  4.520 0.855 4.960 0.925 ;
        RECT  4.870 0.360 4.940 0.615 ;
        RECT  4.800 0.545 4.870 0.615 ;
        RECT  4.730 0.195 4.800 0.455 ;
        RECT  4.660 0.715 4.760 0.785 ;
        RECT  4.590 0.195 4.660 0.785 ;
        RECT  4.480 0.195 4.590 0.265 ;
        RECT  4.450 0.345 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.910 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.910 4.290 0.980 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.345 4.190 0.630 ;
        RECT  3.895 0.345 4.120 0.415 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.345 3.895 0.840 ;
        RECT  3.710 0.345 3.825 0.415 ;
        RECT  3.710 0.770 3.825 0.840 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.910 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.465 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.355 0.335 2.465 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.355 0.405 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.255 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.145 0.195 1.255 0.410 ;
        RECT  0.820 0.340 1.145 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.670 0.500 0.675 0.920 ;
        RECT  0.605 0.340 0.670 0.920 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.605 0.590 ;
        RECT  0.485 0.500 0.590 0.590 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.430 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.830 0.330 0.940 ;
        RECT  0.190 0.195 0.260 0.620 ;
        RECT  0.100 0.540 0.190 0.620 ;
    END
END SEDFQNXD1BWP

MACRO SEDFQNXD2BWP
    CLASS CORE ;
    FOREIGN SEDFQNXD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.505 0.355 5.565 0.815 ;
        RECT  5.495 0.195 5.505 1.035 ;
        RECT  5.435 0.195 5.495 0.475 ;
        RECT  5.435 0.735 5.495 1.035 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.930 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.300 ;
        RECT  3.390 -0.115 5.610 0.115 ;
        RECT  3.320 -0.115 3.390 0.300 ;
        RECT  2.455 -0.115 3.320 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.895 5.690 1.375 ;
        RECT  4.120 1.145 5.610 1.375 ;
        RECT  4.000 1.060 4.120 1.375 ;
        RECT  3.720 1.145 4.000 1.375 ;
        RECT  3.600 1.060 3.720 1.375 ;
        RECT  2.320 1.145 3.600 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.295 0.195 5.365 1.065 ;
        RECT  4.760 0.195 5.295 0.265 ;
        RECT  4.780 0.995 5.295 1.065 ;
        RECT  5.155 0.360 5.225 0.925 ;
        RECT  4.900 0.360 5.155 0.430 ;
        RECT  5.060 0.825 5.155 0.925 ;
        RECT  4.990 0.520 5.040 0.755 ;
        RECT  4.970 0.520 4.990 0.920 ;
        RECT  4.920 0.685 4.970 0.920 ;
        RECT  4.480 0.850 4.920 0.920 ;
        RECT  4.830 0.360 4.900 0.615 ;
        RECT  4.760 0.545 4.830 0.615 ;
        RECT  4.660 0.990 4.780 1.065 ;
        RECT  4.690 0.195 4.760 0.455 ;
        RECT  4.620 0.710 4.720 0.780 ;
        RECT  4.320 0.995 4.660 1.065 ;
        RECT  4.550 0.195 4.620 0.780 ;
        RECT  4.440 0.195 4.550 0.265 ;
        RECT  4.410 0.345 4.480 0.920 ;
        RECT  4.320 0.185 4.440 0.265 ;
        RECT  4.270 0.335 4.340 0.825 ;
        RECT  3.900 0.195 4.320 0.265 ;
        RECT  4.250 0.920 4.320 1.065 ;
        RECT  4.220 0.335 4.270 0.435 ;
        RECT  4.010 0.755 4.270 0.825 ;
        RECT  3.530 0.920 4.250 0.990 ;
        RECT  4.150 0.510 4.200 0.630 ;
        RECT  4.080 0.355 4.150 0.630 ;
        RECT  3.855 0.355 4.080 0.425 ;
        RECT  3.940 0.560 4.010 0.825 ;
        RECT  3.780 0.185 3.900 0.265 ;
        RECT  3.785 0.355 3.855 0.850 ;
        RECT  3.670 0.355 3.785 0.425 ;
        RECT  3.670 0.780 3.785 0.850 ;
        RECT  3.560 0.195 3.780 0.265 ;
        RECT  3.590 0.525 3.700 0.595 ;
        RECT  3.520 0.525 3.590 0.825 ;
        RECT  3.490 0.195 3.560 0.450 ;
        RECT  3.460 0.920 3.530 1.065 ;
        RECT  3.390 0.755 3.520 0.825 ;
        RECT  3.445 0.380 3.490 0.450 ;
        RECT  2.510 0.995 3.460 1.065 ;
        RECT  3.375 0.380 3.445 0.645 ;
        RECT  3.320 0.755 3.390 0.925 ;
        RECT  3.250 0.380 3.375 0.450 ;
        RECT  2.650 0.855 3.320 0.925 ;
        RECT  3.180 0.195 3.250 0.785 ;
        RECT  3.140 0.195 3.180 0.320 ;
        RECT  3.160 0.665 3.180 0.785 ;
        RECT  3.070 0.480 3.110 0.600 ;
        RECT  3.000 0.215 3.070 0.785 ;
        RECT  2.730 0.215 3.000 0.285 ;
        RECT  2.750 0.715 3.000 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.615 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.615 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.600 0.340 0.670 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.600 0.570 ;
        RECT  0.470 0.500 0.590 0.570 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.420 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.525 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.455 0.190 0.640 ;
    END
END SEDFQNXD2BWP

MACRO SEDFQNXD4BWP
    CLASS CORE ;
    FOREIGN SEDFQNXD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.995 0.185 6.065 0.465 ;
        RECT  5.995 0.765 6.065 1.065 ;
        RECT  5.915 0.355 5.995 0.465 ;
        RECT  5.915 0.765 5.995 0.905 ;
        RECT  5.705 0.355 5.915 0.905 ;
        RECT  5.635 0.185 5.705 0.465 ;
        RECT  5.635 0.765 5.705 1.065 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.640 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.470 ;
        RECT  5.910 -0.115 6.170 0.115 ;
        RECT  5.790 -0.115 5.910 0.275 ;
        RECT  3.430 -0.115 5.790 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.675 6.250 1.375 ;
        RECT  5.885 1.145 6.170 1.375 ;
        RECT  5.815 0.975 5.885 1.375 ;
        RECT  4.180 1.145 5.815 1.375 ;
        RECT  4.060 1.060 4.180 1.375 ;
        RECT  3.760 1.145 4.060 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.995 0.185 6.065 0.465 ;
        RECT  5.995 0.765 6.065 1.065 ;
        RECT  5.985 0.355 5.995 0.465 ;
        RECT  5.985 0.765 5.995 0.905 ;
        RECT  5.555 0.520 5.580 0.640 ;
        RECT  5.485 0.210 5.555 1.000 ;
        RECT  4.840 0.210 5.485 0.280 ;
        RECT  5.180 0.930 5.485 1.000 ;
        RECT  5.345 0.375 5.415 0.850 ;
        RECT  4.770 0.375 5.345 0.445 ;
        RECT  5.090 0.780 5.345 0.850 ;
        RECT  4.940 0.545 5.230 0.615 ;
        RECT  5.020 0.780 5.090 1.065 ;
        RECT  4.860 0.995 5.020 1.065 ;
        RECT  4.870 0.545 4.940 0.920 ;
        RECT  4.560 0.850 4.870 0.920 ;
        RECT  4.740 0.990 4.860 1.065 ;
        RECT  4.700 0.700 4.800 0.770 ;
        RECT  4.410 0.995 4.740 1.065 ;
        RECT  4.630 0.195 4.700 0.770 ;
        RECT  4.530 0.195 4.630 0.265 ;
        RECT  4.490 0.350 4.560 0.920 ;
        RECT  4.410 0.185 4.530 0.265 ;
        RECT  4.350 0.345 4.420 0.825 ;
        RECT  3.940 0.195 4.410 0.265 ;
        RECT  4.340 0.920 4.410 1.065 ;
        RECT  4.290 0.345 4.350 0.415 ;
        RECT  4.055 0.755 4.350 0.825 ;
        RECT  3.570 0.920 4.340 0.990 ;
        RECT  4.195 0.510 4.280 0.630 ;
        RECT  4.125 0.345 4.195 0.630 ;
        RECT  3.895 0.345 4.125 0.415 ;
        RECT  3.985 0.500 4.055 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.345 3.895 0.850 ;
        RECT  3.710 0.345 3.825 0.415 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.520 3.150 0.640 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.620 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.620 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.600 0.340 0.670 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.600 0.570 ;
        RECT  0.470 0.500 0.590 0.570 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.420 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.520 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.450 0.190 0.640 ;
    END
END SEDFQNXD4BWP

MACRO SEDFQXD0BWP
    CLASS CORE ;
    FOREIGN SEDFQXD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0246 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 0.215 5.565 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0362 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 -0.115 5.600 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.970 -0.115 2.385 0.115 ;
        RECT  0.900 -0.115 0.970 0.260 ;
        RECT  0.120 -0.115 0.900 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.145 5.600 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.340 0.195 5.410 1.065 ;
        RECT  4.830 0.195 5.340 0.265 ;
        RECT  4.360 0.995 5.340 1.065 ;
        RECT  5.200 0.345 5.270 0.925 ;
        RECT  4.970 0.345 5.200 0.415 ;
        RECT  5.100 0.825 5.200 0.925 ;
        RECT  5.055 0.520 5.125 0.755 ;
        RECT  5.030 0.685 5.055 0.755 ;
        RECT  4.960 0.685 5.030 0.925 ;
        RECT  4.900 0.345 4.970 0.615 ;
        RECT  4.520 0.855 4.960 0.925 ;
        RECT  4.820 0.545 4.900 0.615 ;
        RECT  4.760 0.195 4.830 0.440 ;
        RECT  4.690 0.715 4.760 0.785 ;
        RECT  4.620 0.195 4.690 0.785 ;
        RECT  4.480 0.195 4.620 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.730 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.625 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.625 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.825 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.755 0.195 0.825 0.410 ;
        RECT  0.260 0.195 0.755 0.265 ;
        RECT  0.605 0.335 0.675 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.470 0.495 0.605 0.565 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.405 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.540 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.470 0.190 0.640 ;
    END
END SEDFQXD0BWP

MACRO SEDFQXD1BWP
    CLASS CORE ;
    FOREIGN SEDFQXD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 -0.115 5.600 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.145 5.600 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.335 0.195 5.405 1.065 ;
        RECT  4.830 0.195 5.335 0.265 ;
        RECT  4.820 0.995 5.335 1.065 ;
        RECT  5.195 0.345 5.265 0.925 ;
        RECT  4.970 0.345 5.195 0.415 ;
        RECT  5.100 0.825 5.195 0.925 ;
        RECT  5.055 0.520 5.125 0.755 ;
        RECT  5.030 0.685 5.055 0.755 ;
        RECT  4.960 0.685 5.030 0.915 ;
        RECT  4.900 0.345 4.970 0.615 ;
        RECT  4.520 0.845 4.960 0.915 ;
        RECT  4.820 0.545 4.900 0.615 ;
        RECT  4.760 0.195 4.830 0.440 ;
        RECT  4.700 0.990 4.820 1.065 ;
        RECT  4.690 0.705 4.760 0.775 ;
        RECT  4.360 0.995 4.700 1.065 ;
        RECT  4.620 0.195 4.690 0.775 ;
        RECT  4.480 0.195 4.620 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.915 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.620 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.620 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.600 0.340 0.670 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.600 0.570 ;
        RECT  0.470 0.500 0.590 0.570 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.420 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.510 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.440 0.190 0.640 ;
    END
END SEDFQXD1BWP

MACRO SEDFQXD2BWP
    CLASS CORE ;
    FOREIGN SEDFQXD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.505 0.355 5.565 0.815 ;
        RECT  5.495 0.195 5.505 1.035 ;
        RECT  5.435 0.195 5.495 0.475 ;
        RECT  5.435 0.735 5.495 1.035 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.930 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.300 ;
        RECT  3.390 -0.115 5.610 0.115 ;
        RECT  3.320 -0.115 3.390 0.300 ;
        RECT  2.455 -0.115 3.320 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.235 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.895 5.690 1.375 ;
        RECT  4.120 1.145 5.610 1.375 ;
        RECT  4.000 1.060 4.120 1.375 ;
        RECT  3.720 1.145 4.000 1.375 ;
        RECT  3.600 1.060 3.720 1.375 ;
        RECT  2.320 1.145 3.600 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.295 0.195 5.365 1.065 ;
        RECT  4.785 0.195 5.295 0.265 ;
        RECT  4.780 0.995 5.295 1.065 ;
        RECT  5.155 0.345 5.225 0.925 ;
        RECT  4.930 0.345 5.155 0.415 ;
        RECT  5.060 0.825 5.155 0.925 ;
        RECT  5.015 0.520 5.085 0.755 ;
        RECT  4.990 0.685 5.015 0.755 ;
        RECT  4.920 0.685 4.990 0.920 ;
        RECT  4.860 0.345 4.930 0.615 ;
        RECT  4.480 0.850 4.920 0.920 ;
        RECT  4.780 0.545 4.860 0.615 ;
        RECT  4.715 0.195 4.785 0.440 ;
        RECT  4.660 0.990 4.780 1.065 ;
        RECT  4.645 0.710 4.720 0.780 ;
        RECT  4.320 0.995 4.660 1.065 ;
        RECT  4.575 0.195 4.645 0.780 ;
        RECT  4.440 0.195 4.575 0.265 ;
        RECT  4.480 0.335 4.500 0.465 ;
        RECT  4.410 0.335 4.480 0.920 ;
        RECT  4.320 0.185 4.440 0.265 ;
        RECT  4.270 0.335 4.340 0.825 ;
        RECT  3.900 0.195 4.320 0.265 ;
        RECT  4.250 0.920 4.320 1.065 ;
        RECT  4.220 0.335 4.270 0.435 ;
        RECT  4.010 0.755 4.270 0.825 ;
        RECT  3.530 0.920 4.250 0.990 ;
        RECT  4.150 0.510 4.200 0.630 ;
        RECT  4.080 0.355 4.150 0.630 ;
        RECT  3.855 0.355 4.080 0.425 ;
        RECT  3.940 0.560 4.010 0.825 ;
        RECT  3.780 0.185 3.900 0.265 ;
        RECT  3.785 0.355 3.855 0.850 ;
        RECT  3.670 0.355 3.785 0.425 ;
        RECT  3.670 0.780 3.785 0.850 ;
        RECT  3.560 0.195 3.780 0.265 ;
        RECT  3.590 0.525 3.700 0.595 ;
        RECT  3.520 0.525 3.590 0.825 ;
        RECT  3.490 0.195 3.560 0.450 ;
        RECT  3.460 0.920 3.530 1.065 ;
        RECT  3.390 0.755 3.520 0.825 ;
        RECT  3.445 0.380 3.490 0.450 ;
        RECT  2.510 0.995 3.460 1.065 ;
        RECT  3.375 0.380 3.445 0.645 ;
        RECT  3.320 0.755 3.390 0.925 ;
        RECT  3.250 0.380 3.375 0.450 ;
        RECT  2.650 0.855 3.320 0.925 ;
        RECT  3.180 0.195 3.250 0.785 ;
        RECT  3.140 0.195 3.180 0.320 ;
        RECT  3.160 0.665 3.180 0.785 ;
        RECT  3.070 0.480 3.110 0.600 ;
        RECT  3.000 0.215 3.070 0.785 ;
        RECT  2.730 0.215 3.000 0.285 ;
        RECT  2.750 0.715 3.000 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.620 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.620 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.600 0.340 0.670 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.600 0.570 ;
        RECT  0.470 0.500 0.590 0.570 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.420 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.485 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.415 0.190 0.640 ;
    END
END SEDFQXD2BWP

MACRO SEDFQXD4BWP
    CLASS CORE ;
    FOREIGN SEDFQXD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.275 0.185 6.345 0.465 ;
        RECT  6.275 0.765 6.345 1.065 ;
        RECT  6.195 0.355 6.275 0.465 ;
        RECT  6.195 0.765 6.275 0.905 ;
        RECT  5.985 0.355 6.195 0.905 ;
        RECT  5.915 0.185 5.985 0.465 ;
        RECT  5.915 0.765 5.985 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0202 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.640 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 -0.115 6.580 0.115 ;
        RECT  6.450 -0.115 6.530 0.465 ;
        RECT  6.190 -0.115 6.450 0.115 ;
        RECT  6.070 -0.115 6.190 0.275 ;
        RECT  3.430 -0.115 6.070 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.580 1.375 ;
        RECT  6.450 0.675 6.530 1.375 ;
        RECT  6.165 1.145 6.450 1.375 ;
        RECT  6.095 0.975 6.165 1.375 ;
        RECT  4.590 1.145 6.095 1.375 ;
        RECT  4.470 1.040 4.590 1.375 ;
        RECT  4.180 1.145 4.470 1.375 ;
        RECT  4.060 1.060 4.180 1.375 ;
        RECT  3.760 1.145 4.060 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.275 0.185 6.345 0.465 ;
        RECT  6.275 0.765 6.345 1.065 ;
        RECT  6.265 0.355 6.275 0.465 ;
        RECT  6.265 0.765 6.275 0.905 ;
        RECT  5.760 0.195 5.830 1.065 ;
        RECT  5.210 0.195 5.760 0.265 ;
        RECT  4.730 0.995 5.760 1.065 ;
        RECT  5.620 0.365 5.690 0.920 ;
        RECT  5.370 0.365 5.620 0.435 ;
        RECT  5.540 0.820 5.620 0.920 ;
        RECT  5.470 0.520 5.525 0.750 ;
        RECT  5.455 0.520 5.470 0.925 ;
        RECT  5.400 0.680 5.455 0.925 ;
        RECT  4.920 0.855 5.400 0.925 ;
        RECT  5.300 0.365 5.370 0.615 ;
        RECT  5.220 0.545 5.300 0.615 ;
        RECT  5.140 0.195 5.210 0.460 ;
        RECT  5.070 0.705 5.140 0.775 ;
        RECT  5.000 0.195 5.070 0.775 ;
        RECT  4.870 0.195 5.000 0.265 ;
        RECT  4.850 0.350 4.920 0.925 ;
        RECT  4.750 0.190 4.870 0.265 ;
        RECT  4.710 0.345 4.780 0.830 ;
        RECT  3.940 0.195 4.750 0.265 ;
        RECT  4.660 0.900 4.730 1.065 ;
        RECT  4.270 0.345 4.710 0.415 ;
        RECT  4.055 0.760 4.710 0.830 ;
        RECT  4.045 0.900 4.660 0.970 ;
        RECT  4.200 0.545 4.380 0.615 ;
        RECT  4.130 0.345 4.200 0.615 ;
        RECT  3.895 0.345 4.130 0.415 ;
        RECT  3.985 0.500 4.055 0.830 ;
        RECT  3.975 0.900 4.045 0.990 ;
        RECT  3.570 0.920 3.975 0.990 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.345 3.895 0.850 ;
        RECT  3.710 0.345 3.825 0.415 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.520 3.150 0.640 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.615 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.615 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.600 0.340 0.670 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.590 0.340 0.600 0.570 ;
        RECT  0.470 0.500 0.590 0.570 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.420 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 1.060 ;
        RECT  0.195 0.195 0.260 0.520 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.450 0.190 0.640 ;
    END
END SEDFQXD4BWP

MACRO SEDFXD0BWP
    CLASS CORE ;
    FOREIGN SEDFXD0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0246 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0578 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.005 0.715 5.070 0.785 ;
        RECT  5.005 0.355 5.045 0.495 ;
        RECT  4.935 0.355 5.005 0.785 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.900 0.215 5.985 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0358 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0140 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.905 -0.115 6.020 0.115 ;
        RECT  4.835 -0.115 4.905 0.280 ;
        RECT  3.430 -0.115 4.835 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.125 -0.115 0.890 0.115 ;
        RECT  0.055 -0.115 0.125 0.230 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.145 6.020 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.760 0.215 5.830 1.060 ;
        RECT  5.220 0.215 5.760 0.285 ;
        RECT  5.490 0.990 5.760 1.060 ;
        RECT  5.620 0.370 5.690 0.920 ;
        RECT  5.300 0.370 5.620 0.440 ;
        RECT  5.405 0.850 5.620 0.920 ;
        RECT  5.465 0.520 5.535 0.780 ;
        RECT  5.230 0.710 5.465 0.780 ;
        RECT  5.335 0.850 5.405 1.065 ;
        RECT  4.360 0.995 5.335 1.065 ;
        RECT  5.220 0.545 5.290 0.615 ;
        RECT  5.160 0.710 5.230 0.925 ;
        RECT  5.150 0.215 5.220 0.615 ;
        RECT  4.520 0.855 5.160 0.925 ;
        RECT  4.690 0.715 4.760 0.785 ;
        RECT  4.620 0.195 4.690 0.785 ;
        RECT  4.480 0.195 4.620 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.730 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.470 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.350 0.335 2.470 0.700 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.350 0.405 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.295 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.295 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.275 0.195 0.750 0.265 ;
        RECT  0.670 0.515 0.675 0.920 ;
        RECT  0.605 0.335 0.670 0.920 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.600 0.335 0.605 0.570 ;
        RECT  0.485 0.500 0.600 0.570 ;
        RECT  0.415 0.990 0.520 1.060 ;
        RECT  0.415 0.335 0.510 0.405 ;
        RECT  0.345 0.335 0.415 1.060 ;
        RECT  0.235 0.815 0.345 0.940 ;
        RECT  0.205 0.195 0.275 0.525 ;
        RECT  0.195 0.455 0.205 0.525 ;
        RECT  0.125 0.455 0.195 0.640 ;
    END
END SEDFXD0BWP

MACRO SEDFXD1BWP
    CLASS CORE ;
    FOREIGN SEDFXD1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.350 5.425 0.470 ;
        RECT  5.335 0.775 5.425 1.065 ;
        RECT  5.285 0.775 5.335 0.905 ;
        RECT  5.215 0.350 5.285 0.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.895 0.195 5.985 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 -0.115 6.020 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.775 1.145 6.020 1.375 ;
        RECT  5.705 0.745 5.775 1.375 ;
        RECT  4.160 1.145 5.705 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.210 5.775 0.640 ;
        RECT  4.900 0.210 5.705 0.280 ;
        RECT  5.515 0.370 5.585 0.825 ;
        RECT  5.370 0.545 5.515 0.615 ;
        RECT  4.975 0.370 5.045 1.065 ;
        RECT  4.360 0.995 4.975 1.065 ;
        RECT  4.830 0.210 4.900 0.925 ;
        RECT  4.520 0.855 4.830 0.925 ;
        RECT  4.690 0.695 4.760 0.785 ;
        RECT  4.620 0.195 4.690 0.785 ;
        RECT  4.480 0.195 4.620 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.615 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.615 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.605 0.340 0.675 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.585 0.340 0.605 0.575 ;
        RECT  0.470 0.505 0.585 0.575 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.335 0.510 0.425 ;
        RECT  0.330 0.335 0.400 1.060 ;
        RECT  0.235 0.815 0.330 0.945 ;
        RECT  0.195 0.195 0.260 0.545 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.475 0.190 0.640 ;
    END
END SEDFXD1BWP

MACRO SEDFXD2BWP
    CLASS CORE ;
    FOREIGN SEDFXD2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.425 0.350 5.490 0.420 ;
        RECT  5.425 0.735 5.465 1.045 ;
        RECT  5.355 0.350 5.425 1.045 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.205 0.355 6.265 0.815 ;
        RECT  6.195 0.185 6.205 1.045 ;
        RECT  6.135 0.185 6.195 0.465 ;
        RECT  6.135 0.735 6.195 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.630 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.390 -0.115 6.440 0.115 ;
        RECT  6.310 -0.115 6.390 0.300 ;
        RECT  3.430 -0.115 6.310 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.390 1.145 6.440 1.375 ;
        RECT  6.310 0.895 6.390 1.375 ;
        RECT  6.015 1.145 6.310 1.375 ;
        RECT  5.945 0.745 6.015 1.375 ;
        RECT  5.645 1.145 5.945 1.375 ;
        RECT  5.575 0.735 5.645 1.375 ;
        RECT  5.275 1.145 5.575 1.375 ;
        RECT  5.205 0.675 5.275 1.375 ;
        RECT  4.160 1.145 5.205 1.375 ;
        RECT  4.040 1.060 4.160 1.375 ;
        RECT  3.760 1.145 4.040 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.945 0.210 6.015 0.640 ;
        RECT  4.900 0.210 5.945 0.280 ;
        RECT  5.755 0.360 5.825 1.035 ;
        RECT  5.505 0.545 5.755 0.615 ;
        RECT  4.975 0.370 5.045 1.065 ;
        RECT  4.360 0.995 4.975 1.065 ;
        RECT  4.830 0.210 4.900 0.925 ;
        RECT  4.520 0.855 4.830 0.925 ;
        RECT  4.690 0.695 4.760 0.785 ;
        RECT  4.620 0.195 4.690 0.785 ;
        RECT  4.480 0.195 4.620 0.265 ;
        RECT  4.520 0.335 4.540 0.465 ;
        RECT  4.450 0.335 4.520 0.925 ;
        RECT  4.360 0.185 4.480 0.265 ;
        RECT  4.310 0.335 4.380 0.825 ;
        RECT  3.940 0.195 4.360 0.265 ;
        RECT  4.290 0.920 4.360 1.065 ;
        RECT  4.260 0.335 4.310 0.435 ;
        RECT  4.050 0.755 4.310 0.825 ;
        RECT  3.570 0.920 4.290 0.990 ;
        RECT  4.190 0.510 4.240 0.630 ;
        RECT  4.120 0.355 4.190 0.630 ;
        RECT  3.895 0.355 4.120 0.425 ;
        RECT  3.980 0.560 4.050 0.825 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.355 3.895 0.850 ;
        RECT  3.710 0.355 3.825 0.425 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.480 3.150 0.600 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.620 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.620 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.835 1.585 0.905 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.605 0.335 0.675 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.585 0.335 0.605 0.575 ;
        RECT  0.505 0.505 0.585 0.575 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.345 0.510 0.425 ;
        RECT  0.330 0.345 0.400 1.060 ;
        RECT  0.235 0.815 0.330 0.945 ;
        RECT  0.195 0.195 0.260 0.560 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.490 0.190 0.640 ;
    END
END SEDFXD2BWP

MACRO SEDFXD4BWP
    CLASS CORE ;
    FOREIGN SEDFXD4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.0116 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.495 2.220 0.710 ;
        RECT  1.995 0.495 2.120 0.635 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0274 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.765 0.625 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.350 6.240 0.450 ;
        RECT  6.155 0.765 6.225 1.065 ;
        RECT  6.055 0.765 6.155 0.905 ;
        RECT  5.845 0.350 6.055 0.905 ;
        RECT  5.750 0.350 5.845 0.450 ;
        RECT  5.775 0.765 5.845 1.065 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.255 0.185 7.325 0.465 ;
        RECT  7.255 0.765 7.325 1.065 ;
        RECT  7.175 0.355 7.255 0.465 ;
        RECT  7.175 0.765 7.255 0.865 ;
        RECT  6.965 0.355 7.175 0.865 ;
        RECT  6.895 0.185 6.965 0.465 ;
        RECT  6.895 0.765 6.965 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.0390 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.995 1.420 1.065 ;
        RECT  0.875 0.545 0.945 1.065 ;
        RECT  0.775 0.545 0.875 0.615 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0204 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.505 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.925 0.640 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.510 -0.115 7.560 0.115 ;
        RECT  7.430 -0.115 7.510 0.465 ;
        RECT  7.170 -0.115 7.430 0.115 ;
        RECT  7.050 -0.115 7.170 0.275 ;
        RECT  3.430 -0.115 7.050 0.115 ;
        RECT  3.360 -0.115 3.430 0.300 ;
        RECT  2.455 -0.115 3.360 0.115 ;
        RECT  2.385 -0.115 2.455 0.250 ;
        RECT  0.960 -0.115 2.385 0.115 ;
        RECT  0.890 -0.115 0.960 0.260 ;
        RECT  0.120 -0.115 0.890 0.115 ;
        RECT  0.050 -0.115 0.120 0.230 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.510 1.145 7.560 1.375 ;
        RECT  7.430 0.680 7.510 1.375 ;
        RECT  7.145 1.145 7.430 1.375 ;
        RECT  7.075 0.935 7.145 1.375 ;
        RECT  6.775 1.145 7.075 1.375 ;
        RECT  6.705 0.735 6.775 1.375 ;
        RECT  6.405 1.145 6.705 1.375 ;
        RECT  6.335 0.735 6.405 1.375 ;
        RECT  6.035 1.145 6.335 1.375 ;
        RECT  5.965 0.975 6.035 1.375 ;
        RECT  5.655 1.145 5.965 1.375 ;
        RECT  5.585 0.675 5.655 1.375 ;
        RECT  4.590 1.145 5.585 1.375 ;
        RECT  4.470 1.040 4.590 1.375 ;
        RECT  4.180 1.145 4.470 1.375 ;
        RECT  4.060 1.060 4.180 1.375 ;
        RECT  3.760 1.145 4.060 1.375 ;
        RECT  3.640 1.060 3.760 1.375 ;
        RECT  2.320 1.145 3.640 1.375 ;
        RECT  2.200 1.060 2.320 1.375 ;
        RECT  0.805 1.145 2.200 1.375 ;
        RECT  0.735 1.030 0.805 1.375 ;
        RECT  0.125 1.145 0.735 1.375 ;
        RECT  0.055 0.825 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.255 0.185 7.325 0.465 ;
        RECT  7.255 0.765 7.325 1.065 ;
        RECT  7.245 0.355 7.255 0.465 ;
        RECT  7.245 0.765 7.255 0.865 ;
        RECT  6.125 0.350 6.240 0.450 ;
        RECT  6.155 0.765 6.225 1.065 ;
        RECT  6.125 0.765 6.155 0.905 ;
        RECT  5.750 0.350 5.775 0.450 ;
        RECT  6.705 0.210 6.775 0.640 ;
        RECT  5.280 0.210 6.705 0.280 ;
        RECT  6.515 0.350 6.585 1.070 ;
        RECT  6.210 0.545 6.515 0.615 ;
        RECT  5.355 0.380 5.430 1.065 ;
        RECT  4.730 0.995 5.355 1.065 ;
        RECT  5.210 0.210 5.280 0.925 ;
        RECT  4.920 0.855 5.210 0.925 ;
        RECT  5.080 0.705 5.140 0.775 ;
        RECT  5.010 0.195 5.080 0.775 ;
        RECT  4.870 0.195 5.010 0.265 ;
        RECT  4.850 0.350 4.920 0.925 ;
        RECT  4.750 0.190 4.870 0.265 ;
        RECT  4.710 0.345 4.780 0.820 ;
        RECT  3.940 0.195 4.750 0.265 ;
        RECT  4.660 0.900 4.730 1.065 ;
        RECT  4.270 0.345 4.710 0.415 ;
        RECT  4.055 0.750 4.710 0.820 ;
        RECT  4.015 0.900 4.660 0.970 ;
        RECT  4.200 0.545 4.380 0.615 ;
        RECT  4.130 0.345 4.200 0.615 ;
        RECT  3.895 0.345 4.130 0.415 ;
        RECT  3.985 0.500 4.055 0.820 ;
        RECT  3.945 0.900 4.015 0.990 ;
        RECT  3.570 0.920 3.945 0.990 ;
        RECT  3.820 0.185 3.940 0.265 ;
        RECT  3.825 0.345 3.895 0.850 ;
        RECT  3.710 0.345 3.825 0.415 ;
        RECT  3.710 0.780 3.825 0.850 ;
        RECT  3.600 0.195 3.820 0.265 ;
        RECT  3.630 0.525 3.740 0.595 ;
        RECT  3.560 0.525 3.630 0.825 ;
        RECT  3.530 0.195 3.600 0.450 ;
        RECT  3.500 0.920 3.570 1.065 ;
        RECT  3.430 0.755 3.560 0.825 ;
        RECT  3.485 0.380 3.530 0.450 ;
        RECT  2.510 0.995 3.500 1.065 ;
        RECT  3.415 0.380 3.485 0.645 ;
        RECT  3.360 0.755 3.430 0.925 ;
        RECT  3.290 0.380 3.415 0.450 ;
        RECT  2.650 0.855 3.360 0.925 ;
        RECT  3.220 0.195 3.290 0.785 ;
        RECT  3.175 0.195 3.220 0.320 ;
        RECT  3.170 0.715 3.220 0.785 ;
        RECT  3.085 0.520 3.150 0.640 ;
        RECT  3.015 0.215 3.085 0.785 ;
        RECT  2.770 0.215 3.015 0.285 ;
        RECT  2.750 0.715 3.015 0.785 ;
        RECT  2.460 0.335 2.670 0.405 ;
        RECT  2.580 0.780 2.650 0.925 ;
        RECT  1.925 0.780 2.580 0.850 ;
        RECT  2.440 0.920 2.510 1.065 ;
        RECT  2.460 0.610 2.470 0.710 ;
        RECT  2.360 0.335 2.460 0.710 ;
        RECT  1.655 0.920 2.440 0.990 ;
        RECT  2.260 0.335 2.360 0.405 ;
        RECT  2.350 0.610 2.360 0.710 ;
        RECT  2.190 0.195 2.260 0.405 ;
        RECT  2.030 0.195 2.190 0.265 ;
        RECT  1.925 0.355 2.110 0.425 ;
        RECT  1.910 0.185 2.030 0.265 ;
        RECT  1.855 0.335 1.925 0.850 ;
        RECT  1.260 0.195 1.910 0.265 ;
        RECT  1.425 0.335 1.855 0.405 ;
        RECT  1.810 0.780 1.855 0.850 ;
        RECT  1.655 0.475 1.775 0.545 ;
        RECT  1.585 0.475 1.655 0.990 ;
        RECT  1.410 0.840 1.585 0.910 ;
        RECT  1.355 0.335 1.425 0.550 ;
        RECT  1.085 0.480 1.355 0.550 ;
        RECT  1.085 0.835 1.310 0.905 ;
        RECT  1.160 0.195 1.260 0.270 ;
        RECT  1.090 0.195 1.160 0.410 ;
        RECT  0.820 0.340 1.090 0.410 ;
        RECT  1.015 0.480 1.085 0.905 ;
        RECT  0.750 0.195 0.820 0.410 ;
        RECT  0.260 0.195 0.750 0.265 ;
        RECT  0.605 0.335 0.675 0.900 ;
        RECT  0.520 0.990 0.640 1.075 ;
        RECT  0.585 0.335 0.605 0.575 ;
        RECT  0.500 0.505 0.585 0.575 ;
        RECT  0.400 0.990 0.520 1.060 ;
        RECT  0.400 0.345 0.510 0.435 ;
        RECT  0.330 0.345 0.400 1.060 ;
        RECT  0.235 0.815 0.330 0.945 ;
        RECT  0.195 0.195 0.260 0.545 ;
        RECT  0.190 0.195 0.195 0.640 ;
        RECT  0.125 0.475 0.190 0.640 ;
    END
END SEDFXD4BWP

MACRO TAPCELLBWP
    CLASS CORE ;
    FOREIGN TAPCELLBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.410 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.780 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
END TAPCELLBWP

MACRO TIEHBWP
    CLASS CORE ;
    FOREIGN TIEHBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0451 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.735 0.385 1.045 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.115 0.420 0.115 ;
        RECT  0.115 -0.115 0.185 0.465 ;
        RECT  0.000 -0.115 0.115 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.145 0.420 1.375 ;
        RECT  0.115 0.745 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 0.185 0.365 0.615 ;
        RECT  0.200 0.545 0.295 0.615 ;
    END
END TIEHBWP

MACRO TIELBWP
    CLASS CORE ;
    FOREIGN TIELBWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0341 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.185 0.385 0.485 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 -0.115 0.420 0.115 ;
        RECT  0.115 -0.115 0.185 0.465 ;
        RECT  0.000 -0.115 0.115 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.145 0.420 1.375 ;
        RECT  0.115 0.745 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 0.555 0.365 1.045 ;
        RECT  0.190 0.555 0.295 0.625 ;
    END
END TIELBWP

MACRO XNR2D0BWP
    CLASS CORE ;
    FOREIGN XNR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.195 1.365 1.045 ;
        RECT  1.275 0.195 1.295 0.355 ;
        RECT  1.275 0.840 1.295 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.350 1.085 0.630 ;
        RECT  0.980 0.510 1.015 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0318 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.170 0.270 ;
        RECT  0.260 -0.115 1.070 0.115 ;
        RECT  0.260 0.345 0.380 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.145 1.400 1.375 ;
        RECT  1.070 1.010 1.170 1.375 ;
        RECT  0.330 1.145 1.070 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.500 1.225 0.770 ;
        RECT  1.155 0.500 1.190 0.920 ;
        RECT  1.120 0.700 1.155 0.920 ;
        RECT  0.765 0.850 1.120 0.920 ;
        RECT  0.910 0.200 0.990 0.270 ;
        RECT  0.910 0.710 0.990 0.780 ;
        RECT  0.770 0.995 0.930 1.075 ;
        RECT  0.840 0.200 0.910 0.780 ;
        RECT  0.370 0.200 0.840 0.270 ;
        RECT  0.560 0.995 0.770 1.065 ;
        RECT  0.685 0.350 0.765 0.920 ;
        RECT  0.490 0.860 0.560 1.065 ;
        RECT  0.485 0.350 0.555 0.790 ;
        RECT  0.125 0.860 0.490 0.930 ;
        RECT  0.405 0.720 0.485 0.790 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR2D0BWP

MACRO XNR2D1BWP
    CLASS CORE ;
    FOREIGN XNR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.185 1.365 1.060 ;
        RECT  1.275 0.185 1.295 0.465 ;
        RECT  1.270 0.900 1.295 1.060 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.350 1.085 0.630 ;
        RECT  0.960 0.510 1.015 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.170 0.270 ;
        RECT  0.260 -0.115 1.070 0.115 ;
        RECT  0.260 0.345 0.340 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.145 1.400 1.375 ;
        RECT  1.070 0.995 1.170 1.375 ;
        RECT  0.330 1.145 1.070 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.190 0.515 1.225 0.770 ;
        RECT  1.155 0.515 1.190 0.915 ;
        RECT  1.120 0.700 1.155 0.915 ;
        RECT  0.740 0.845 1.120 0.915 ;
        RECT  0.890 0.705 1.000 0.775 ;
        RECT  0.890 0.210 0.990 0.280 ;
        RECT  0.740 0.995 0.900 1.075 ;
        RECT  0.820 0.210 0.890 0.775 ;
        RECT  0.490 0.210 0.820 0.280 ;
        RECT  0.670 0.350 0.740 0.915 ;
        RECT  0.560 0.995 0.740 1.065 ;
        RECT  0.490 0.860 0.560 1.065 ;
        RECT  0.485 0.350 0.555 0.775 ;
        RECT  0.370 0.200 0.490 0.280 ;
        RECT  0.125 0.860 0.490 0.930 ;
        RECT  0.405 0.705 0.485 0.775 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR2D1BWP

MACRO XNR2D2BWP
    CLASS CORE ;
    FOREIGN XNR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.395 1.505 0.910 ;
        RECT  1.305 0.395 1.435 0.465 ;
        RECT  1.200 0.840 1.435 0.910 ;
        RECT  1.235 0.185 1.305 0.465 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.630 ;
        RECT  0.970 0.530 1.015 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.315 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.350 0.350 0.420 ;
        RECT  0.190 -0.115 0.260 0.420 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.145 1.540 1.375 ;
        RECT  1.410 0.990 1.490 1.375 ;
        RECT  1.140 1.145 1.410 1.375 ;
        RECT  1.040 1.000 1.140 1.375 ;
        RECT  0.330 1.145 1.040 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.540 1.340 0.620 ;
        RECT  1.155 0.540 1.225 0.770 ;
        RECT  1.120 0.700 1.155 0.770 ;
        RECT  1.050 0.700 1.120 0.910 ;
        RECT  0.725 0.840 1.050 0.910 ;
        RECT  0.885 0.700 0.970 0.770 ;
        RECT  0.885 0.210 0.960 0.280 ;
        RECT  0.815 0.210 0.885 0.770 ;
        RECT  0.710 0.995 0.870 1.075 ;
        RECT  0.470 0.210 0.815 0.280 ;
        RECT  0.655 0.350 0.725 0.910 ;
        RECT  0.560 0.995 0.710 1.065 ;
        RECT  0.490 0.860 0.560 1.065 ;
        RECT  0.475 0.350 0.545 0.790 ;
        RECT  0.125 0.860 0.490 0.930 ;
        RECT  0.395 0.720 0.475 0.790 ;
        RECT  0.350 0.195 0.470 0.280 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR2D2BWP

MACRO XNR2D4BWP
    CLASS CORE ;
    FOREIGN XNR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.195 2.705 0.480 ;
        RECT  2.695 0.775 2.705 1.055 ;
        RECT  2.635 0.195 2.695 1.055 ;
        RECT  2.485 0.355 2.635 0.905 ;
        RECT  2.345 0.355 2.485 0.480 ;
        RECT  2.345 0.775 2.485 0.905 ;
        RECT  2.275 0.195 2.345 0.480 ;
        RECT  2.275 0.775 2.345 1.055 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0720 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 0.495 2.065 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.485 ;
        RECT  2.540 -0.115 2.810 0.115 ;
        RECT  2.440 -0.115 2.540 0.275 ;
        RECT  0.670 -0.115 2.440 0.115 ;
        RECT  0.590 -0.115 0.670 0.450 ;
        RECT  0.330 -0.115 0.590 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.665 2.890 1.375 ;
        RECT  2.540 1.145 2.810 1.375 ;
        RECT  2.440 0.985 2.540 1.375 ;
        RECT  0.310 1.145 2.440 1.375 ;
        RECT  0.230 0.885 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.480 ;
        RECT  2.345 0.775 2.415 0.905 ;
        RECT  2.275 0.195 2.345 0.480 ;
        RECT  2.275 0.775 2.345 1.055 ;
        RECT  2.205 0.550 2.395 0.620 ;
        RECT  2.135 0.195 2.205 1.050 ;
        RECT  1.430 0.195 2.135 0.265 ;
        RECT  1.690 0.980 2.135 1.050 ;
        RECT  1.850 0.340 2.010 0.410 ;
        RECT  1.850 0.840 2.010 0.910 ;
        RECT  1.780 0.340 1.850 0.910 ;
        RECT  1.640 0.335 1.710 0.910 ;
        RECT  1.510 0.335 1.640 0.405 ;
        RECT  1.610 0.840 1.640 0.910 ;
        RECT  1.530 0.840 1.610 1.050 ;
        RECT  1.400 0.510 1.570 0.580 ;
        RECT  0.490 0.980 1.530 1.050 ;
        RECT  1.350 0.195 1.430 0.405 ;
        RECT  1.350 0.700 1.430 0.910 ;
        RECT  1.330 0.510 1.400 0.620 ;
        RECT  1.010 0.335 1.350 0.405 ;
        RECT  1.010 0.700 1.350 0.770 ;
        RECT  1.090 0.540 1.330 0.620 ;
        RECT  0.870 0.195 1.270 0.265 ;
        RECT  0.870 0.840 1.270 0.910 ;
        RECT  0.940 0.335 1.010 0.770 ;
        RECT  0.800 0.195 0.870 0.910 ;
        RECT  0.770 0.195 0.800 0.340 ;
        RECT  0.490 0.520 0.730 0.640 ;
        RECT  0.410 0.185 0.490 1.050 ;
        RECT  0.130 0.330 0.410 0.405 ;
        RECT  0.130 0.725 0.410 0.795 ;
        RECT  0.050 0.245 0.130 0.405 ;
        RECT  0.050 0.725 0.130 1.045 ;
    END
END XNR2D4BWP

MACRO XNR3D0BWP
    CLASS CORE ;
    FOREIGN XNR3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.210 2.485 1.045 ;
        RECT  2.395 0.210 2.415 0.370 ;
        RECT  2.395 0.885 2.415 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.165 0.215 2.205 0.485 ;
        RECT  2.135 0.215 2.165 0.640 ;
        RECT  2.095 0.415 2.135 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.630 1.085 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 2.520 0.115 ;
        RECT  1.380 -0.115 1.460 0.465 ;
        RECT  1.090 -0.115 1.380 0.115 ;
        RECT  1.010 -0.115 1.090 0.330 ;
        RECT  0.310 -0.115 1.010 0.115 ;
        RECT  0.230 -0.115 0.310 0.350 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.530 1.145 2.520 1.375 ;
        RECT  1.460 0.835 1.530 1.375 ;
        RECT  1.345 0.835 1.460 0.905 ;
        RECT  0.330 1.145 1.460 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.325 0.510 2.345 0.670 ;
        RECT  2.275 0.510 2.325 1.050 ;
        RECT  2.255 0.600 2.275 1.050 ;
        RECT  1.880 0.980 2.255 1.050 ;
        RECT  2.020 0.840 2.090 0.910 ;
        RECT  1.950 0.205 2.020 0.910 ;
        RECT  1.600 0.205 1.950 0.275 ;
        RECT  1.810 0.365 1.880 1.050 ;
        RECT  1.720 0.365 1.810 0.435 ;
        RECT  1.795 0.870 1.810 1.050 ;
        RECT  1.670 0.520 1.740 0.765 ;
        RECT  1.270 0.695 1.670 0.765 ;
        RECT  1.530 0.205 1.600 0.615 ;
        RECT  1.420 0.545 1.530 0.615 ;
        RECT  0.765 0.995 1.380 1.065 ;
        RECT  1.265 0.330 1.270 0.765 ;
        RECT  1.190 0.330 1.265 0.900 ;
        RECT  0.835 0.195 0.905 0.910 ;
        RECT  0.485 0.195 0.835 0.265 ;
        RECT  0.695 0.340 0.765 1.065 ;
        RECT  0.570 0.340 0.695 0.410 ;
        RECT  0.590 0.900 0.695 0.980 ;
        RECT  0.555 0.500 0.625 0.800 ;
        RECT  0.445 0.730 0.555 0.800 ;
        RECT  0.415 0.195 0.485 0.620 ;
        RECT  0.375 0.730 0.445 0.930 ;
        RECT  0.340 0.540 0.415 0.620 ;
        RECT  0.130 0.860 0.375 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D0BWP

MACRO XNR3D1BWP
    CLASS CORE ;
    FOREIGN XNR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.045 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.730 2.415 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.165 0.215 2.205 0.485 ;
        RECT  2.135 0.215 2.165 0.640 ;
        RECT  2.095 0.415 2.135 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.495 1.085 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.455 -0.115 2.520 0.115 ;
        RECT  1.385 -0.115 1.455 0.465 ;
        RECT  1.090 -0.115 1.385 0.115 ;
        RECT  1.010 -0.115 1.090 0.420 ;
        RECT  0.310 -0.115 1.010 0.115 ;
        RECT  0.230 -0.115 0.310 0.355 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.145 2.520 1.375 ;
        RECT  1.450 0.835 1.520 1.375 ;
        RECT  1.350 0.835 1.450 0.905 ;
        RECT  0.330 1.145 1.450 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.325 0.515 2.345 0.670 ;
        RECT  2.275 0.515 2.325 1.050 ;
        RECT  2.255 0.600 2.275 1.050 ;
        RECT  1.880 0.980 2.255 1.050 ;
        RECT  2.020 0.840 2.090 0.910 ;
        RECT  1.950 0.205 2.020 0.910 ;
        RECT  1.600 0.205 1.950 0.275 ;
        RECT  1.810 0.365 1.880 1.050 ;
        RECT  1.720 0.365 1.810 0.435 ;
        RECT  1.790 0.880 1.810 1.050 ;
        RECT  1.670 0.520 1.740 0.765 ;
        RECT  1.270 0.695 1.670 0.765 ;
        RECT  1.530 0.205 1.600 0.615 ;
        RECT  1.420 0.545 1.530 0.615 ;
        RECT  0.765 0.995 1.380 1.065 ;
        RECT  1.190 0.330 1.270 0.900 ;
        RECT  0.835 0.195 0.905 0.915 ;
        RECT  0.485 0.195 0.835 0.265 ;
        RECT  0.695 0.340 0.765 1.065 ;
        RECT  0.590 0.340 0.695 0.410 ;
        RECT  0.590 0.900 0.695 0.980 ;
        RECT  0.555 0.490 0.625 0.800 ;
        RECT  0.445 0.730 0.555 0.800 ;
        RECT  0.415 0.195 0.485 0.620 ;
        RECT  0.375 0.730 0.445 0.930 ;
        RECT  0.325 0.540 0.415 0.620 ;
        RECT  0.130 0.860 0.375 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D1BWP

MACRO XNR3D2BWP
    CLASS CORE ;
    FOREIGN XNR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.355 3.045 0.905 ;
        RECT  2.975 0.185 2.985 1.035 ;
        RECT  2.915 0.185 2.975 0.465 ;
        RECT  2.915 0.735 2.975 1.035 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.665 0.640 ;
        RECT  2.555 0.495 2.625 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.355 1.085 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.300 ;
        RECT  1.500 -0.115 3.095 0.115 ;
        RECT  1.430 -0.115 1.500 0.390 ;
        RECT  1.110 -0.115 1.430 0.115 ;
        RECT  1.030 -0.115 1.110 0.275 ;
        RECT  0.260 -0.115 1.030 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.965 3.170 1.375 ;
        RECT  2.800 1.145 3.090 1.375 ;
        RECT  2.720 0.800 2.800 1.375 ;
        RECT  1.510 1.145 2.720 1.375 ;
        RECT  1.440 0.780 1.510 1.375 ;
        RECT  0.330 1.145 1.440 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.830 0.520 2.870 0.640 ;
        RECT  2.760 0.210 2.830 0.640 ;
        RECT  2.345 0.210 2.760 0.280 ;
        RECT  2.485 0.350 2.640 0.420 ;
        RECT  2.485 0.905 2.620 0.985 ;
        RECT  2.415 0.350 2.485 1.065 ;
        RECT  1.650 0.995 2.415 1.065 ;
        RECT  2.275 0.210 2.345 0.925 ;
        RECT  2.000 0.210 2.275 0.280 ;
        RECT  1.870 0.855 2.275 0.925 ;
        RECT  2.090 0.350 2.170 0.785 ;
        RECT  1.790 0.715 2.090 0.785 ;
        RECT  1.930 0.210 2.000 0.445 ;
        RECT  1.870 0.375 1.930 0.445 ;
        RECT  1.760 0.185 1.860 0.290 ;
        RECT  1.720 0.370 1.790 0.915 ;
        RECT  1.650 0.220 1.760 0.290 ;
        RECT  1.580 0.220 1.650 0.530 ;
        RECT  1.580 0.600 1.650 1.065 ;
        RECT  1.310 0.460 1.580 0.530 ;
        RECT  1.500 0.600 1.580 0.670 ;
        RECT  1.050 0.995 1.370 1.065 ;
        RECT  1.220 0.300 1.310 0.900 ;
        RECT  0.970 0.845 1.050 1.065 ;
        RECT  0.710 0.845 0.970 0.915 ;
        RECT  0.820 0.195 0.920 0.775 ;
        RECT  0.700 0.995 0.860 1.075 ;
        RECT  0.340 0.195 0.820 0.270 ;
        RECT  0.630 0.350 0.710 0.915 ;
        RECT  0.550 0.995 0.700 1.065 ;
        RECT  0.480 0.860 0.550 1.065 ;
        RECT  0.450 0.350 0.530 0.780 ;
        RECT  0.125 0.860 0.480 0.930 ;
        RECT  0.390 0.710 0.450 0.780 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR3D2BWP

MACRO XNR3D4BWP
    CLASS CORE ;
    FOREIGN XNR3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.485 ;
        RECT  3.955 0.745 3.965 1.065 ;
        RECT  3.895 0.185 3.955 1.065 ;
        RECT  3.745 0.355 3.895 0.905 ;
        RECT  3.605 0.355 3.745 0.485 ;
        RECT  3.605 0.745 3.745 0.905 ;
        RECT  3.535 0.185 3.605 0.485 ;
        RECT  3.535 0.745 3.605 1.065 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.945 0.355 3.045 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.110 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 -0.115 4.200 0.115 ;
        RECT  4.075 -0.115 4.145 0.485 ;
        RECT  3.800 -0.115 4.075 0.115 ;
        RECT  3.700 -0.115 3.800 0.275 ;
        RECT  1.490 -0.115 3.700 0.115 ;
        RECT  1.410 -0.115 1.490 0.485 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.270 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 1.145 4.200 1.375 ;
        RECT  4.075 0.685 4.145 1.375 ;
        RECT  3.800 1.145 4.075 1.375 ;
        RECT  3.700 0.985 3.800 1.375 ;
        RECT  3.440 1.145 3.700 1.375 ;
        RECT  3.340 1.010 3.440 1.375 ;
        RECT  3.080 1.145 3.340 1.375 ;
        RECT  2.980 1.010 3.080 1.375 ;
        RECT  2.360 1.145 2.980 1.375 ;
        RECT  2.260 0.990 2.360 1.375 ;
        RECT  1.140 1.145 2.260 1.375 ;
        RECT  1.040 0.990 1.140 1.375 ;
        RECT  0.330 1.145 1.040 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.355 3.675 0.485 ;
        RECT  3.605 0.745 3.675 0.905 ;
        RECT  3.535 0.185 3.605 0.485 ;
        RECT  3.535 0.745 3.605 1.065 ;
        RECT  3.450 0.555 3.540 0.625 ;
        RECT  3.380 0.210 3.450 0.940 ;
        RECT  2.300 0.210 3.380 0.280 ;
        RECT  2.890 0.870 3.380 0.940 ;
        RECT  3.230 0.730 3.290 0.800 ;
        RECT  3.150 0.360 3.230 0.800 ;
        RECT  2.845 0.730 3.150 0.800 ;
        RECT  2.820 0.870 2.890 1.065 ;
        RECT  2.775 0.350 2.845 0.800 ;
        RECT  2.590 0.995 2.820 1.065 ;
        RECT  2.710 0.730 2.775 0.800 ;
        RECT  2.640 0.730 2.710 0.920 ;
        RECT  2.550 0.565 2.650 0.635 ;
        RECT  2.330 0.850 2.640 0.920 ;
        RECT  2.480 0.470 2.550 0.780 ;
        RECT  2.465 0.470 2.480 0.545 ;
        RECT  2.410 0.710 2.480 0.780 ;
        RECT  2.395 0.350 2.465 0.545 ;
        RECT  1.990 0.475 2.395 0.545 ;
        RECT  2.260 0.615 2.330 0.920 ;
        RECT  2.230 0.210 2.300 0.405 ;
        RECT  2.090 0.615 2.260 0.685 ;
        RECT  1.845 0.335 2.230 0.405 ;
        RECT  1.670 0.840 2.180 0.910 ;
        RECT  1.670 0.195 2.100 0.265 ;
        RECT  1.915 0.475 1.990 0.610 ;
        RECT  1.845 0.700 1.960 0.770 ;
        RECT  1.800 0.980 1.960 1.075 ;
        RECT  1.775 0.335 1.845 0.770 ;
        RECT  1.470 0.980 1.800 1.050 ;
        RECT  1.590 0.195 1.670 0.910 ;
        RECT  1.400 0.845 1.470 1.050 ;
        RECT  0.725 0.845 1.400 0.915 ;
        RECT  1.310 0.705 1.350 0.775 ;
        RECT  1.230 0.195 1.310 0.775 ;
        RECT  0.930 0.705 1.230 0.775 ;
        RECT  0.850 0.200 0.930 0.775 ;
        RECT  0.720 0.995 0.880 1.075 ;
        RECT  0.350 0.200 0.850 0.270 ;
        RECT  0.655 0.350 0.725 0.915 ;
        RECT  0.560 0.995 0.720 1.065 ;
        RECT  0.490 0.860 0.560 1.065 ;
        RECT  0.475 0.350 0.545 0.790 ;
        RECT  0.125 0.860 0.490 0.930 ;
        RECT  0.395 0.720 0.475 0.790 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR3D4BWP

MACRO XNR4D0BWP
    CLASS CORE ;
    FOREIGN XNR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.215 2.410 0.295 ;
        RECT  2.345 0.715 2.410 0.785 ;
        RECT  2.275 0.215 2.345 0.785 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.100 0.655 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.355 2.640 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.495 3.465 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.410 -0.115 3.640 0.115 ;
        RECT  3.340 -0.115 3.410 0.415 ;
        RECT  2.600 -0.115 3.340 0.115 ;
        RECT  2.480 -0.115 2.600 0.275 ;
        RECT  1.480 -0.115 2.480 0.115 ;
        RECT  1.410 -0.115 1.480 0.445 ;
        RECT  1.130 -0.115 1.410 0.115 ;
        RECT  1.050 -0.115 1.130 0.280 ;
        RECT  0.260 -0.115 1.050 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.390 1.145 3.640 1.375 ;
        RECT  3.290 0.990 3.390 1.375 ;
        RECT  1.530 1.145 3.290 1.375 ;
        RECT  1.430 0.985 1.530 1.375 ;
        RECT  0.330 1.145 1.430 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.535 0.290 3.605 1.000 ;
        RECT  3.510 0.290 3.535 0.430 ;
        RECT  3.515 0.850 3.535 1.000 ;
        RECT  3.080 0.850 3.515 0.920 ;
        RECT  3.200 0.200 3.270 0.660 ;
        RECT  2.800 0.200 3.200 0.270 ;
        RECT  3.010 0.530 3.080 0.920 ;
        RECT  2.940 0.350 2.955 0.470 ;
        RECT  2.870 0.350 2.940 1.065 ;
        RECT  2.530 0.995 2.870 1.065 ;
        RECT  2.730 0.200 2.800 0.915 ;
        RECT  2.670 0.200 2.730 0.280 ;
        RECT  2.650 0.845 2.730 0.915 ;
        RECT  2.460 0.855 2.530 1.065 ;
        RECT  2.205 0.855 2.460 0.925 ;
        RECT  2.050 0.995 2.380 1.065 ;
        RECT  2.130 0.195 2.205 0.925 ;
        RECT  1.620 0.195 2.130 0.265 ;
        RECT  1.980 0.335 2.050 1.065 ;
        RECT  1.910 0.335 1.980 0.405 ;
        RECT  1.870 0.995 1.980 1.065 ;
        RECT  1.840 0.510 1.910 0.915 ;
        RECT  1.305 0.845 1.840 0.915 ;
        RECT  1.700 0.335 1.770 0.775 ;
        RECT  1.630 0.705 1.700 0.775 ;
        RECT  1.550 0.195 1.620 0.615 ;
        RECT  1.480 0.545 1.550 0.615 ;
        RECT  0.750 0.995 1.340 1.065 ;
        RECT  1.235 0.315 1.305 0.915 ;
        RECT  0.870 0.195 0.940 0.925 ;
        RECT  0.450 0.195 0.870 0.265 ;
        RECT  0.830 0.825 0.870 0.925 ;
        RECT  0.680 0.340 0.750 1.065 ;
        RECT  0.670 0.340 0.680 0.885 ;
        RECT  0.635 0.755 0.670 0.885 ;
        RECT  0.490 0.985 0.610 1.055 ;
        RECT  0.430 0.355 0.510 0.800 ;
        RECT  0.420 0.870 0.490 1.055 ;
        RECT  0.330 0.185 0.450 0.285 ;
        RECT  0.130 0.870 0.420 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.305 0.120 0.445 ;
        RECT  0.035 0.305 0.105 1.050 ;
    END
END XNR4D0BWP

MACRO XNR4D1BWP
    CLASS CORE ;
    FOREIGN XNR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.0862 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.715 2.450 0.785 ;
        RECT  2.345 0.215 2.410 0.440 ;
        RECT  2.270 0.215 2.345 0.785 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0310 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0284 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.010 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.520 2.655 0.640 ;
        RECT  2.550 0.355 2.625 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.495 3.465 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.410 -0.115 3.640 0.115 ;
        RECT  3.340 -0.115 3.410 0.415 ;
        RECT  2.610 -0.115 3.340 0.115 ;
        RECT  2.510 -0.115 2.610 0.275 ;
        RECT  1.480 -0.115 2.510 0.115 ;
        RECT  1.410 -0.115 1.480 0.445 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.390 1.145 3.640 1.375 ;
        RECT  3.290 0.990 3.390 1.375 ;
        RECT  1.520 1.145 3.290 1.375 ;
        RECT  1.440 0.985 1.520 1.375 ;
        RECT  0.330 1.145 1.440 1.375 ;
        RECT  0.210 1.030 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.535 0.290 3.605 1.000 ;
        RECT  3.515 0.290 3.535 0.430 ;
        RECT  3.515 0.850 3.535 1.000 ;
        RECT  3.100 0.850 3.515 0.920 ;
        RECT  3.200 0.200 3.270 0.660 ;
        RECT  2.820 0.200 3.200 0.270 ;
        RECT  3.030 0.530 3.100 0.920 ;
        RECT  2.960 0.350 3.030 0.430 ;
        RECT  2.890 0.350 2.960 1.045 ;
        RECT  2.530 0.975 2.890 1.045 ;
        RECT  2.750 0.200 2.820 0.905 ;
        RECT  2.700 0.345 2.750 0.415 ;
        RECT  2.670 0.835 2.750 0.905 ;
        RECT  2.460 0.855 2.530 1.045 ;
        RECT  2.200 0.855 2.460 0.925 ;
        RECT  2.180 0.995 2.340 1.075 ;
        RECT  2.130 0.195 2.200 0.925 ;
        RECT  2.050 0.995 2.180 1.065 ;
        RECT  1.620 0.195 2.130 0.265 ;
        RECT  1.980 0.335 2.050 1.065 ;
        RECT  1.910 0.335 1.980 0.405 ;
        RECT  1.870 0.995 1.980 1.065 ;
        RECT  1.840 0.520 1.910 0.915 ;
        RECT  1.310 0.845 1.840 0.915 ;
        RECT  1.700 0.335 1.770 0.775 ;
        RECT  1.630 0.705 1.700 0.775 ;
        RECT  1.620 0.545 1.630 0.615 ;
        RECT  1.550 0.195 1.620 0.615 ;
        RECT  1.510 0.545 1.550 0.615 ;
        RECT  1.220 0.995 1.360 1.075 ;
        RECT  1.230 0.305 1.310 0.915 ;
        RECT  0.780 0.995 1.220 1.065 ;
        RECT  1.080 0.355 1.150 0.915 ;
        RECT  0.950 0.355 1.080 0.425 ;
        RECT  0.850 0.845 1.080 0.915 ;
        RECT  0.870 0.200 0.950 0.425 ;
        RECT  0.330 0.200 0.870 0.270 ;
        RECT  0.710 0.350 0.780 1.065 ;
        RECT  0.690 0.350 0.710 0.905 ;
        RECT  0.645 0.745 0.690 0.905 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.430 0.350 0.510 0.820 ;
        RECT  0.420 0.890 0.490 1.055 ;
        RECT  0.130 0.890 0.420 0.960 ;
        RECT  0.105 0.890 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D1BWP

MACRO XNR4D2BWP
    CLASS CORE ;
    FOREIGN XNR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.770 ;
        RECT  2.550 0.355 2.555 0.475 ;
        RECT  2.470 0.650 2.555 0.770 ;
        RECT  2.470 0.195 2.550 0.475 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0306 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.010 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.520 2.795 0.640 ;
        RECT  2.695 0.355 2.765 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0306 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.495 3.605 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.780 0.115 ;
        RECT  3.520 -0.115 3.590 0.425 ;
        RECT  2.740 -0.115 3.520 0.115 ;
        RECT  3.430 0.355 3.520 0.425 ;
        RECT  2.640 -0.115 2.740 0.275 ;
        RECT  2.370 -0.115 2.640 0.115 ;
        RECT  2.290 -0.115 2.370 0.290 ;
        RECT  1.480 -0.115 2.290 0.115 ;
        RECT  1.410 -0.115 1.480 0.465 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.145 3.780 1.375 ;
        RECT  3.450 1.010 3.570 1.375 ;
        RECT  2.370 1.145 3.450 1.375 ;
        RECT  2.290 0.980 2.370 1.375 ;
        RECT  1.540 1.145 2.290 1.375 ;
        RECT  1.420 0.985 1.540 1.375 ;
        RECT  0.330 1.145 1.420 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.290 3.745 1.050 ;
        RECT  3.660 0.290 3.675 0.440 ;
        RECT  3.650 0.870 3.675 1.050 ;
        RECT  3.305 0.870 3.650 0.940 ;
        RECT  2.950 0.200 3.450 0.270 ;
        RECT  3.270 0.365 3.350 0.800 ;
        RECT  3.235 0.870 3.305 1.055 ;
        RECT  3.160 0.985 3.235 1.055 ;
        RECT  3.090 0.700 3.145 0.830 ;
        RECT  3.020 0.365 3.090 1.050 ;
        RECT  2.520 0.980 3.020 1.050 ;
        RECT  2.880 0.200 2.950 0.910 ;
        RECT  2.835 0.320 2.880 0.440 ;
        RECT  2.810 0.840 2.880 0.910 ;
        RECT  2.450 0.840 2.520 1.050 ;
        RECT  2.390 0.840 2.450 0.910 ;
        RECT  2.320 0.380 2.390 0.910 ;
        RECT  2.180 0.380 2.320 0.450 ;
        RECT  2.180 0.840 2.320 0.910 ;
        RECT  2.040 0.520 2.240 0.640 ;
        RECT  2.110 0.200 2.180 0.450 ;
        RECT  2.110 0.840 2.180 1.050 ;
        RECT  1.620 0.200 2.110 0.270 ;
        RECT  1.970 0.350 2.040 1.055 ;
        RECT  1.870 0.350 1.970 0.420 ;
        RECT  1.860 0.985 1.970 1.055 ;
        RECT  1.830 0.525 1.900 0.915 ;
        RECT  1.310 0.845 1.830 0.915 ;
        RECT  1.690 0.350 1.760 0.775 ;
        RECT  1.610 0.705 1.690 0.775 ;
        RECT  1.550 0.200 1.620 0.630 ;
        RECT  1.510 0.530 1.550 0.630 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  1.230 0.325 1.310 0.915 ;
        RECT  0.780 0.995 1.220 1.065 ;
        RECT  1.080 0.355 1.150 0.915 ;
        RECT  0.950 0.355 1.080 0.425 ;
        RECT  0.850 0.845 1.080 0.915 ;
        RECT  0.870 0.200 0.950 0.425 ;
        RECT  0.330 0.200 0.870 0.270 ;
        RECT  0.710 0.350 0.780 1.065 ;
        RECT  0.690 0.350 0.710 0.905 ;
        RECT  0.645 0.745 0.690 0.905 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.510 0.710 0.520 0.810 ;
        RECT  0.430 0.350 0.510 0.810 ;
        RECT  0.420 0.880 0.490 1.055 ;
        RECT  0.420 0.710 0.430 0.810 ;
        RECT  0.130 0.880 0.420 0.950 ;
        RECT  0.105 0.880 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D2BWP

MACRO XNR4D4BWP
    CLASS CORE ;
    FOREIGN XNR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.2160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.650 3.120 0.790 ;
        RECT  3.030 0.195 3.110 0.485 ;
        RECT  2.975 0.345 3.030 0.485 ;
        RECT  2.765 0.345 2.975 0.790 ;
        RECT  2.720 0.345 2.765 0.485 ;
        RECT  2.640 0.650 2.765 0.790 ;
        RECT  2.640 0.195 2.720 0.485 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0306 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.495 1.090 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.520 3.355 0.640 ;
        RECT  3.255 0.355 3.325 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0306 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.495 4.165 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.340 0.115 ;
        RECT  4.080 -0.115 4.150 0.425 ;
        RECT  3.300 -0.115 4.080 0.115 ;
        RECT  4.010 0.355 4.080 0.425 ;
        RECT  3.200 -0.115 3.300 0.275 ;
        RECT  2.930 -0.115 3.200 0.115 ;
        RECT  2.830 -0.115 2.930 0.275 ;
        RECT  2.530 -0.115 2.830 0.115 ;
        RECT  2.460 -0.115 2.530 0.290 ;
        RECT  1.140 -0.115 2.460 0.115 ;
        RECT  1.040 -0.115 1.140 0.420 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.145 4.340 1.375 ;
        RECT  4.010 1.010 4.130 1.375 ;
        RECT  2.940 1.145 4.010 1.375 ;
        RECT  2.820 1.010 2.940 1.375 ;
        RECT  2.550 1.145 2.820 1.375 ;
        RECT  2.430 1.010 2.550 1.375 ;
        RECT  2.090 1.145 2.430 1.375 ;
        RECT  1.970 1.010 2.090 1.375 ;
        RECT  0.330 1.145 1.970 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.045 0.650 3.120 0.790 ;
        RECT  3.045 0.195 3.110 0.485 ;
        RECT  2.640 0.195 2.695 0.485 ;
        RECT  2.640 0.650 2.695 0.790 ;
        RECT  4.235 0.300 4.305 1.050 ;
        RECT  4.220 0.300 4.235 0.440 ;
        RECT  4.210 0.870 4.235 1.050 ;
        RECT  3.865 0.870 4.210 0.940 ;
        RECT  3.510 0.200 4.010 0.270 ;
        RECT  3.830 0.350 3.910 0.800 ;
        RECT  3.795 0.870 3.865 1.055 ;
        RECT  3.720 0.985 3.795 1.055 ;
        RECT  3.650 0.700 3.705 0.830 ;
        RECT  3.580 0.350 3.650 1.050 ;
        RECT  3.260 0.980 3.580 1.050 ;
        RECT  3.440 0.200 3.510 0.910 ;
        RECT  3.395 0.320 3.440 0.440 ;
        RECT  3.370 0.840 3.440 0.910 ;
        RECT  3.180 0.870 3.260 1.050 ;
        RECT  2.560 0.870 3.180 0.940 ;
        RECT  2.490 0.370 2.560 0.940 ;
        RECT  2.390 0.370 2.490 0.440 ;
        RECT  2.340 0.520 2.410 0.940 ;
        RECT  2.320 0.210 2.390 0.440 ;
        RECT  1.690 0.870 2.340 0.940 ;
        RECT  2.065 0.210 2.320 0.280 ;
        RECT  2.240 0.710 2.270 0.800 ;
        RECT  2.170 0.350 2.240 0.800 ;
        RECT  1.865 0.730 2.170 0.800 ;
        RECT  1.985 0.210 2.065 0.660 ;
        RECT  1.520 0.210 1.985 0.280 ;
        RECT  1.790 0.350 1.865 0.800 ;
        RECT  1.610 0.350 1.690 1.060 ;
        RECT  1.450 0.210 1.520 1.020 ;
        RECT  1.410 0.325 1.450 0.445 ;
        RECT  1.390 0.940 1.450 1.020 ;
        RECT  1.310 0.530 1.380 0.650 ;
        RECT  1.235 0.350 1.310 0.880 ;
        RECT  0.780 0.980 1.310 1.050 ;
        RECT  0.920 0.840 0.990 0.910 ;
        RECT  0.920 0.320 0.960 0.420 ;
        RECT  0.850 0.200 0.920 0.910 ;
        RECT  0.340 0.200 0.850 0.270 ;
        RECT  0.710 0.350 0.780 1.050 ;
        RECT  0.690 0.350 0.710 0.910 ;
        RECT  0.635 0.840 0.690 0.910 ;
        RECT  0.550 0.990 0.640 1.060 ;
        RECT  0.480 0.870 0.550 1.060 ;
        RECT  0.465 0.345 0.540 0.800 ;
        RECT  0.130 0.870 0.480 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D4BWP

MACRO XOR2D0BWP
    CLASS CORE ;
    FOREIGN XOR2D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.365 1.070 ;
        RECT  1.275 0.345 1.295 0.465 ;
        RECT  1.260 0.970 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.085 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 -0.115 1.400 0.115 ;
        RECT  1.080 -0.115 1.160 0.425 ;
        RECT  0.260 -0.115 1.080 0.115 ;
        RECT  0.260 0.355 0.330 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 1.400 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.165 0.530 1.225 0.905 ;
        RECT  1.155 0.530 1.165 1.050 ;
        RECT  1.095 0.835 1.155 1.050 ;
        RECT  0.775 0.980 1.095 1.050 ;
        RECT  0.915 0.840 1.005 0.910 ;
        RECT  0.915 0.330 1.000 0.400 ;
        RECT  0.845 0.200 0.915 0.910 ;
        RECT  0.330 0.200 0.845 0.270 ;
        RECT  0.705 0.350 0.775 1.050 ;
        RECT  0.685 0.350 0.705 0.790 ;
        RECT  0.650 0.700 0.685 0.790 ;
        RECT  0.545 0.860 0.635 1.070 ;
        RECT  0.510 0.365 0.580 0.780 ;
        RECT  0.125 0.860 0.545 0.930 ;
        RECT  0.415 0.365 0.510 0.435 ;
        RECT  0.450 0.700 0.510 0.780 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.315 0.120 0.450 ;
        RECT  0.035 0.315 0.105 1.040 ;
    END
END XOR2D0BWP

MACRO XOR2D1BWP
    CLASS CORE ;
    FOREIGN XOR2D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.200 1.365 1.070 ;
        RECT  1.275 0.200 1.295 0.460 ;
        RECT  1.260 0.970 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.985 0.520 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0340 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 -0.115 1.400 0.115 ;
        RECT  1.080 -0.115 1.160 0.275 ;
        RECT  0.260 -0.115 1.080 0.115 ;
        RECT  0.260 0.355 0.330 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.145 1.400 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.520 1.225 0.835 ;
        RECT  1.145 0.765 1.155 0.835 ;
        RECT  1.075 0.765 1.145 1.050 ;
        RECT  0.775 0.980 1.075 1.050 ;
        RECT  0.915 0.840 0.995 0.910 ;
        RECT  0.915 0.305 0.945 0.425 ;
        RECT  0.845 0.200 0.915 0.910 ;
        RECT  0.330 0.200 0.845 0.270 ;
        RECT  0.705 0.350 0.775 1.050 ;
        RECT  0.685 0.350 0.705 0.790 ;
        RECT  0.650 0.700 0.685 0.790 ;
        RECT  0.545 0.860 0.635 1.070 ;
        RECT  0.510 0.365 0.580 0.780 ;
        RECT  0.125 0.860 0.545 0.930 ;
        RECT  0.415 0.365 0.510 0.435 ;
        RECT  0.440 0.700 0.510 0.780 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.305 0.120 0.445 ;
        RECT  0.035 0.305 0.105 1.040 ;
    END
END XOR2D1BWP

MACRO XOR2D2BWP
    CLASS CORE ;
    FOREIGN XOR2D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.395 1.505 0.920 ;
        RECT  1.310 0.395 1.435 0.465 ;
        RECT  1.210 0.850 1.435 0.920 ;
        RECT  1.230 0.185 1.310 0.465 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.990 0.510 1.015 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.410 -0.115 1.490 0.315 ;
        RECT  1.150 -0.115 1.410 0.115 ;
        RECT  1.030 -0.115 1.150 0.255 ;
        RECT  0.260 -0.115 1.030 0.115 ;
        RECT  0.260 0.355 0.340 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.990 1.500 1.375 ;
        RECT  1.150 1.145 1.400 1.375 ;
        RECT  1.030 1.010 1.150 1.375 ;
        RECT  0.330 1.145 1.030 1.375 ;
        RECT  0.210 1.020 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.545 1.320 0.615 ;
        RECT  1.155 0.545 1.225 0.780 ;
        RECT  1.130 0.710 1.155 0.780 ;
        RECT  1.060 0.710 1.130 0.930 ;
        RECT  0.765 0.860 1.060 0.930 ;
        RECT  0.920 0.720 0.970 0.790 ;
        RECT  0.920 0.300 0.945 0.420 ;
        RECT  0.850 0.200 0.920 0.790 ;
        RECT  0.330 0.200 0.850 0.270 ;
        RECT  0.695 0.350 0.765 0.930 ;
        RECT  0.645 0.690 0.695 0.810 ;
        RECT  0.550 0.990 0.650 1.060 ;
        RECT  0.490 0.365 0.560 0.810 ;
        RECT  0.480 0.880 0.550 1.060 ;
        RECT  0.430 0.365 0.490 0.435 ;
        RECT  0.395 0.730 0.490 0.810 ;
        RECT  0.125 0.880 0.480 0.950 ;
        RECT  0.105 0.880 0.125 1.055 ;
        RECT  0.105 0.300 0.120 0.450 ;
        RECT  0.035 0.300 0.105 1.055 ;
    END
END XOR2D2BWP

MACRO XOR2D4BWP
    CLASS CORE ;
    FOREIGN XOR2D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.195 2.705 0.480 ;
        RECT  2.695 0.775 2.705 1.055 ;
        RECT  2.635 0.195 2.695 1.055 ;
        RECT  2.485 0.355 2.635 0.905 ;
        RECT  2.345 0.355 2.485 0.480 ;
        RECT  2.345 0.775 2.485 0.905 ;
        RECT  2.275 0.195 2.345 0.480 ;
        RECT  2.275 0.775 2.345 1.055 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0568 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.065 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.485 ;
        RECT  2.540 -0.115 2.810 0.115 ;
        RECT  2.440 -0.115 2.540 0.275 ;
        RECT  0.670 -0.115 2.440 0.115 ;
        RECT  0.590 -0.115 0.670 0.450 ;
        RECT  0.330 -0.115 0.590 0.115 ;
        RECT  0.210 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.210 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.665 2.890 1.375 ;
        RECT  2.540 1.145 2.810 1.375 ;
        RECT  2.440 0.985 2.540 1.375 ;
        RECT  0.310 1.145 2.440 1.375 ;
        RECT  0.230 0.995 0.310 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.415 0.480 ;
        RECT  2.345 0.775 2.415 0.905 ;
        RECT  2.275 0.195 2.345 0.480 ;
        RECT  2.275 0.775 2.345 1.055 ;
        RECT  2.205 0.550 2.395 0.620 ;
        RECT  2.135 0.200 2.205 1.050 ;
        RECT  1.960 0.200 2.135 0.270 ;
        RECT  1.690 0.980 2.135 1.050 ;
        RECT  1.850 0.340 2.010 0.410 ;
        RECT  1.850 0.840 2.010 0.910 ;
        RECT  1.890 0.195 1.960 0.270 ;
        RECT  1.430 0.195 1.890 0.265 ;
        RECT  1.780 0.340 1.850 0.910 ;
        RECT  1.640 0.335 1.710 0.860 ;
        RECT  1.510 0.335 1.640 0.405 ;
        RECT  1.605 0.790 1.640 0.860 ;
        RECT  1.535 0.790 1.605 1.050 ;
        RECT  1.400 0.510 1.570 0.580 ;
        RECT  0.490 0.980 1.535 1.050 ;
        RECT  1.350 0.195 1.430 0.405 ;
        RECT  1.350 0.700 1.430 0.910 ;
        RECT  1.330 0.510 1.400 0.620 ;
        RECT  1.010 0.335 1.350 0.405 ;
        RECT  1.010 0.700 1.350 0.770 ;
        RECT  1.090 0.540 1.330 0.620 ;
        RECT  0.870 0.195 1.270 0.265 ;
        RECT  0.870 0.840 1.270 0.910 ;
        RECT  0.940 0.335 1.010 0.770 ;
        RECT  0.800 0.195 0.870 0.910 ;
        RECT  0.770 0.195 0.800 0.340 ;
        RECT  0.490 0.520 0.730 0.640 ;
        RECT  0.410 0.185 0.490 1.050 ;
        RECT  0.130 0.330 0.410 0.405 ;
        RECT  0.130 0.845 0.410 0.915 ;
        RECT  0.050 0.245 0.130 0.405 ;
        RECT  0.050 0.845 0.130 1.005 ;
    END
END XOR2D4BWP

MACRO XOR3D0BWP
    CLASS CORE ;
    FOREIGN XOR3D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.215 2.485 1.045 ;
        RECT  2.395 0.215 2.415 0.385 ;
        RECT  2.400 0.840 2.415 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 0.215 2.205 0.485 ;
        RECT  2.135 0.215 2.170 0.660 ;
        RECT  2.100 0.415 2.135 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.495 1.095 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 2.520 0.115 ;
        RECT  1.390 -0.115 1.460 0.465 ;
        RECT  1.120 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.120 0.415 ;
        RECT  0.310 -0.115 1.020 0.115 ;
        RECT  0.230 -0.115 0.310 0.330 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.550 1.145 2.520 1.375 ;
        RECT  1.480 0.835 1.550 1.375 ;
        RECT  1.370 0.835 1.480 0.905 ;
        RECT  0.330 1.145 1.480 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.330 0.515 2.345 0.650 ;
        RECT  2.275 0.515 2.330 1.055 ;
        RECT  2.260 0.590 2.275 1.055 ;
        RECT  1.890 0.985 2.260 1.055 ;
        RECT  1.960 0.205 2.030 0.905 ;
        RECT  1.600 0.205 1.960 0.275 ;
        RECT  1.820 0.365 1.890 1.055 ;
        RECT  1.710 0.365 1.820 0.435 ;
        RECT  1.770 0.850 1.820 1.055 ;
        RECT  1.680 0.520 1.750 0.765 ;
        RECT  1.290 0.695 1.680 0.765 ;
        RECT  1.530 0.205 1.600 0.615 ;
        RECT  1.420 0.545 1.530 0.615 ;
        RECT  0.750 0.995 1.400 1.065 ;
        RECT  1.210 0.330 1.290 0.900 ;
        RECT  0.915 0.845 0.960 0.915 ;
        RECT  0.845 0.195 0.915 0.915 ;
        RECT  0.490 0.195 0.845 0.265 ;
        RECT  0.820 0.845 0.845 0.915 ;
        RECT  0.675 0.335 0.750 1.065 ;
        RECT  0.610 0.335 0.675 0.415 ;
        RECT  0.610 0.870 0.675 0.940 ;
        RECT  0.535 0.550 0.605 0.790 ;
        RECT  0.425 0.720 0.535 0.790 ;
        RECT  0.425 0.195 0.490 0.480 ;
        RECT  0.420 0.195 0.425 0.640 ;
        RECT  0.345 0.720 0.425 0.930 ;
        RECT  0.355 0.410 0.420 0.640 ;
        RECT  0.130 0.860 0.345 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XOR3D0BWP

MACRO XOR3D1BWP
    CLASS CORE ;
    FOREIGN XOR3D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.045 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.400 0.725 2.415 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 0.215 2.205 0.485 ;
        RECT  2.135 0.215 2.170 0.660 ;
        RECT  2.100 0.415 2.135 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0338 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.970 0.495 1.015 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.460 -0.115 2.520 0.115 ;
        RECT  1.390 -0.115 1.460 0.465 ;
        RECT  1.120 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.120 0.415 ;
        RECT  0.310 -0.115 1.020 0.115 ;
        RECT  0.230 -0.115 0.310 0.330 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.550 1.145 2.520 1.375 ;
        RECT  1.480 0.835 1.550 1.375 ;
        RECT  1.370 0.835 1.480 0.905 ;
        RECT  0.330 1.145 1.480 1.375 ;
        RECT  0.210 1.000 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.330 0.515 2.345 0.650 ;
        RECT  2.275 0.515 2.330 1.055 ;
        RECT  2.260 0.590 2.275 1.055 ;
        RECT  1.890 0.985 2.260 1.055 ;
        RECT  1.960 0.205 2.030 0.905 ;
        RECT  1.600 0.205 1.960 0.275 ;
        RECT  1.820 0.365 1.890 1.055 ;
        RECT  1.710 0.365 1.820 0.435 ;
        RECT  1.770 0.850 1.820 1.055 ;
        RECT  1.680 0.520 1.750 0.765 ;
        RECT  1.290 0.695 1.680 0.765 ;
        RECT  1.530 0.205 1.600 0.620 ;
        RECT  1.420 0.550 1.530 0.620 ;
        RECT  0.760 0.995 1.400 1.065 ;
        RECT  1.210 0.330 1.290 0.900 ;
        RECT  0.830 0.195 0.900 0.915 ;
        RECT  0.490 0.195 0.830 0.265 ;
        RECT  0.685 0.335 0.760 1.065 ;
        RECT  0.610 0.335 0.685 0.415 ;
        RECT  0.675 0.870 0.685 1.065 ;
        RECT  0.610 0.870 0.675 0.940 ;
        RECT  0.545 0.545 0.615 0.790 ;
        RECT  0.425 0.720 0.545 0.790 ;
        RECT  0.425 0.195 0.490 0.470 ;
        RECT  0.420 0.195 0.425 0.640 ;
        RECT  0.345 0.720 0.425 0.930 ;
        RECT  0.355 0.400 0.420 0.640 ;
        RECT  0.130 0.860 0.345 0.930 ;
        RECT  0.105 0.195 0.130 0.355 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END XOR3D1BWP

MACRO XOR3D2BWP
    CLASS CORE ;
    FOREIGN XOR3D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.765 ;
        RECT  2.590 0.355 2.695 0.465 ;
        RECT  2.570 0.695 2.695 0.765 ;
        RECT  2.500 0.185 2.590 0.465 ;
        RECT  2.480 0.695 2.570 1.055 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.735 2.350 1.050 ;
        RECT  2.275 0.520 2.290 1.050 ;
        RECT  2.220 0.520 2.275 0.805 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.100 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.280 ;
        RECT  1.560 -0.115 2.670 0.115 ;
        RECT  1.440 -0.115 1.560 0.200 ;
        RECT  1.130 -0.115 1.440 0.115 ;
        RECT  1.050 -0.115 1.130 0.285 ;
        RECT  0.260 -0.115 1.050 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.885 2.750 1.375 ;
        RECT  1.500 1.145 2.670 1.375 ;
        RECT  1.430 0.780 1.500 1.375 ;
        RECT  0.330 1.145 1.430 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.430 0.545 2.610 0.615 ;
        RECT  2.360 0.220 2.430 0.615 ;
        RECT  2.010 0.220 2.360 0.290 ;
        RECT  2.150 0.360 2.230 0.430 ;
        RECT  2.150 0.885 2.175 1.065 ;
        RECT  2.080 0.360 2.150 1.065 ;
        RECT  1.640 0.995 2.080 1.065 ;
        RECT  1.940 0.220 2.010 0.915 ;
        RECT  1.880 0.350 1.940 0.510 ;
        RECT  1.870 0.835 1.940 0.915 ;
        RECT  1.750 0.200 1.860 0.270 ;
        RECT  1.720 0.410 1.790 0.920 ;
        RECT  1.680 0.200 1.750 0.340 ;
        RECT  1.630 0.410 1.720 0.480 ;
        RECT  1.330 0.270 1.680 0.340 ;
        RECT  1.570 0.560 1.640 1.065 ;
        RECT  1.480 0.560 1.570 0.635 ;
        RECT  0.765 0.995 1.350 1.065 ;
        RECT  1.250 0.270 1.330 0.900 ;
        RECT  0.920 0.855 0.990 0.925 ;
        RECT  0.920 0.200 0.940 0.480 ;
        RECT  0.850 0.200 0.920 0.925 ;
        RECT  0.340 0.200 0.850 0.270 ;
        RECT  0.695 0.345 0.765 1.065 ;
        RECT  0.655 0.785 0.695 0.915 ;
        RECT  0.540 0.990 0.620 1.060 ;
        RECT  0.470 0.870 0.540 1.060 ;
        RECT  0.450 0.345 0.530 0.800 ;
        RECT  0.125 0.870 0.470 0.940 ;
        RECT  0.105 0.870 0.125 1.050 ;
        RECT  0.105 0.300 0.120 0.450 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR3D2BWP

MACRO XOR3D4BWP
    CLASS CORE ;
    FOREIGN XOR3D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 3.965 0.485 ;
        RECT  3.955 0.745 3.965 1.065 ;
        RECT  3.895 0.185 3.955 1.065 ;
        RECT  3.745 0.355 3.895 0.905 ;
        RECT  3.605 0.355 3.745 0.485 ;
        RECT  3.605 0.745 3.745 0.905 ;
        RECT  3.535 0.185 3.605 0.485 ;
        RECT  3.535 0.745 3.605 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.355 3.070 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0864 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.115 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 -0.115 4.200 0.115 ;
        RECT  4.075 -0.115 4.145 0.485 ;
        RECT  3.800 -0.115 4.075 0.115 ;
        RECT  3.700 -0.115 3.800 0.275 ;
        RECT  1.490 -0.115 3.700 0.115 ;
        RECT  1.410 -0.115 1.490 0.485 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.270 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 1.145 4.200 1.375 ;
        RECT  4.075 0.755 4.145 1.375 ;
        RECT  3.800 1.145 4.075 1.375 ;
        RECT  3.700 0.985 3.800 1.375 ;
        RECT  3.440 1.145 3.700 1.375 ;
        RECT  3.340 1.010 3.440 1.375 ;
        RECT  3.080 1.145 3.340 1.375 ;
        RECT  2.980 1.010 3.080 1.375 ;
        RECT  2.360 1.145 2.980 1.375 ;
        RECT  2.260 0.990 2.360 1.375 ;
        RECT  1.130 1.145 2.260 1.375 ;
        RECT  1.030 0.990 1.130 1.375 ;
        RECT  0.330 1.145 1.030 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.355 3.675 0.485 ;
        RECT  3.605 0.745 3.675 0.905 ;
        RECT  3.535 0.185 3.605 0.485 ;
        RECT  3.535 0.745 3.605 1.065 ;
        RECT  3.450 0.555 3.540 0.625 ;
        RECT  3.380 0.210 3.450 0.940 ;
        RECT  2.300 0.210 3.380 0.280 ;
        RECT  2.890 0.870 3.380 0.940 ;
        RECT  3.230 0.730 3.290 0.800 ;
        RECT  3.150 0.350 3.230 0.800 ;
        RECT  2.850 0.730 3.150 0.800 ;
        RECT  2.820 0.870 2.890 1.065 ;
        RECT  2.770 0.350 2.850 0.800 ;
        RECT  2.590 0.995 2.820 1.065 ;
        RECT  2.710 0.730 2.770 0.800 ;
        RECT  2.640 0.730 2.710 0.920 ;
        RECT  2.550 0.565 2.650 0.635 ;
        RECT  2.330 0.850 2.640 0.920 ;
        RECT  2.480 0.470 2.550 0.780 ;
        RECT  2.465 0.470 2.480 0.545 ;
        RECT  2.410 0.710 2.480 0.780 ;
        RECT  2.395 0.350 2.465 0.545 ;
        RECT  1.990 0.475 2.395 0.545 ;
        RECT  2.260 0.615 2.330 0.920 ;
        RECT  2.230 0.210 2.300 0.405 ;
        RECT  2.090 0.615 2.260 0.685 ;
        RECT  1.845 0.335 2.230 0.405 ;
        RECT  1.670 0.840 2.180 0.910 ;
        RECT  1.670 0.195 2.100 0.265 ;
        RECT  1.915 0.475 1.990 0.610 ;
        RECT  1.845 0.700 1.960 0.770 ;
        RECT  1.800 0.980 1.960 1.075 ;
        RECT  1.775 0.335 1.845 0.770 ;
        RECT  1.470 0.980 1.800 1.050 ;
        RECT  1.590 0.195 1.670 0.910 ;
        RECT  1.400 0.845 1.470 1.050 ;
        RECT  0.760 0.845 1.400 0.915 ;
        RECT  1.305 0.705 1.350 0.775 ;
        RECT  1.235 0.195 1.305 0.775 ;
        RECT  0.945 0.705 1.235 0.775 ;
        RECT  0.875 0.200 0.945 0.775 ;
        RECT  0.340 0.200 0.875 0.270 ;
        RECT  0.830 0.685 0.875 0.775 ;
        RECT  0.690 0.345 0.760 0.915 ;
        RECT  0.600 0.840 0.690 0.915 ;
        RECT  0.520 0.990 0.630 1.060 ;
        RECT  0.440 0.345 0.520 0.800 ;
        RECT  0.450 0.870 0.520 1.060 ;
        RECT  0.125 0.870 0.450 0.940 ;
        RECT  0.105 0.870 0.125 1.050 ;
        RECT  0.105 0.320 0.120 0.450 ;
        RECT  0.035 0.320 0.105 1.050 ;
    END
END XOR3D4BWP

MACRO XOR4D0BWP
    CLASS CORE ;
    FOREIGN XOR4D0BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0664 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.345 0.905 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.990 0.520 1.015 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0144 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.520 2.650 0.640 ;
        RECT  2.555 0.355 2.625 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.495 3.465 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.640 0.115 ;
        RECT  3.380 -0.115 3.450 0.425 ;
        RECT  1.480 -0.115 3.380 0.115 ;
        RECT  3.290 0.355 3.380 0.425 ;
        RECT  1.410 -0.115 1.480 0.460 ;
        RECT  1.150 -0.115 1.410 0.115 ;
        RECT  1.030 -0.115 1.150 0.275 ;
        RECT  0.260 -0.115 1.030 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.145 3.640 1.375 ;
        RECT  3.310 1.010 3.430 1.375 ;
        RECT  1.540 1.145 3.310 1.375 ;
        RECT  1.420 0.985 1.540 1.375 ;
        RECT  0.330 1.145 1.420 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.535 0.300 3.605 1.050 ;
        RECT  3.520 0.300 3.535 0.440 ;
        RECT  3.510 0.870 3.535 1.050 ;
        RECT  3.165 0.870 3.510 0.940 ;
        RECT  2.810 0.200 3.310 0.270 ;
        RECT  3.095 0.870 3.165 1.055 ;
        RECT  3.020 0.985 3.095 1.055 ;
        RECT  2.950 0.710 3.050 0.790 ;
        RECT  2.880 0.350 2.950 1.060 ;
        RECT  2.485 0.990 2.880 1.060 ;
        RECT  2.740 0.200 2.810 0.910 ;
        RECT  2.695 0.315 2.740 0.435 ;
        RECT  2.670 0.840 2.740 0.910 ;
        RECT  2.415 0.200 2.485 1.060 ;
        RECT  1.620 0.200 2.415 0.270 ;
        RECT  2.180 0.990 2.415 1.060 ;
        RECT  2.040 0.530 2.205 0.650 ;
        RECT  2.110 0.890 2.180 1.060 ;
        RECT  1.970 0.360 2.040 1.055 ;
        RECT  1.850 0.360 1.970 0.440 ;
        RECT  1.850 0.985 1.970 1.055 ;
        RECT  1.830 0.520 1.900 0.915 ;
        RECT  1.310 0.845 1.830 0.915 ;
        RECT  1.690 0.360 1.760 0.775 ;
        RECT  1.610 0.700 1.690 0.775 ;
        RECT  1.550 0.200 1.620 0.620 ;
        RECT  1.480 0.540 1.550 0.620 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  1.220 0.345 1.310 0.915 ;
        RECT  0.780 0.995 1.220 1.065 ;
        RECT  0.920 0.845 0.990 0.915 ;
        RECT  0.920 0.200 0.945 0.320 ;
        RECT  0.850 0.200 0.920 0.915 ;
        RECT  0.330 0.200 0.850 0.270 ;
        RECT  0.710 0.350 0.780 1.065 ;
        RECT  0.690 0.350 0.710 0.875 ;
        RECT  0.645 0.745 0.690 0.875 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.430 0.350 0.510 0.800 ;
        RECT  0.420 0.870 0.490 1.055 ;
        RECT  0.130 0.870 0.420 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D0BWP

MACRO XOR4D1BWP
    CLASS CORE ;
    FOREIGN XOR4D1BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.0985 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.345 0.905 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.010 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.520 2.650 0.640 ;
        RECT  2.555 0.355 2.625 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.495 3.465 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.640 0.115 ;
        RECT  3.380 -0.115 3.450 0.425 ;
        RECT  1.480 -0.115 3.380 0.115 ;
        RECT  3.290 0.355 3.380 0.425 ;
        RECT  1.410 -0.115 1.480 0.460 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.145 3.640 1.375 ;
        RECT  3.310 1.010 3.430 1.375 ;
        RECT  1.540 1.145 3.310 1.375 ;
        RECT  1.420 0.985 1.540 1.375 ;
        RECT  0.330 1.145 1.420 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.535 0.300 3.605 1.050 ;
        RECT  3.520 0.300 3.535 0.440 ;
        RECT  3.510 0.870 3.535 1.050 ;
        RECT  3.165 0.870 3.510 0.940 ;
        RECT  2.810 0.200 3.310 0.270 ;
        RECT  3.095 0.870 3.165 1.055 ;
        RECT  3.020 0.985 3.095 1.055 ;
        RECT  2.950 0.710 3.050 0.790 ;
        RECT  2.880 0.350 2.950 1.060 ;
        RECT  2.485 0.990 2.880 1.060 ;
        RECT  2.740 0.200 2.810 0.910 ;
        RECT  2.695 0.300 2.740 0.420 ;
        RECT  2.670 0.840 2.740 0.910 ;
        RECT  2.415 0.200 2.485 1.060 ;
        RECT  1.620 0.200 2.415 0.270 ;
        RECT  2.180 0.990 2.415 1.060 ;
        RECT  2.040 0.510 2.205 0.630 ;
        RECT  2.110 0.890 2.180 1.060 ;
        RECT  1.970 0.360 2.040 1.055 ;
        RECT  1.850 0.360 1.970 0.440 ;
        RECT  1.850 0.985 1.970 1.055 ;
        RECT  1.830 0.520 1.900 0.915 ;
        RECT  1.310 0.845 1.830 0.915 ;
        RECT  1.690 0.360 1.760 0.775 ;
        RECT  1.610 0.700 1.690 0.775 ;
        RECT  1.550 0.200 1.620 0.620 ;
        RECT  1.480 0.540 1.550 0.620 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  1.230 0.185 1.310 0.915 ;
        RECT  0.780 0.995 1.220 1.065 ;
        RECT  1.080 0.345 1.150 0.915 ;
        RECT  0.950 0.345 1.080 0.415 ;
        RECT  0.850 0.845 1.080 0.915 ;
        RECT  0.870 0.200 0.950 0.415 ;
        RECT  0.330 0.200 0.870 0.270 ;
        RECT  0.710 0.350 0.780 1.065 ;
        RECT  0.690 0.350 0.710 0.830 ;
        RECT  0.645 0.700 0.690 0.830 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.430 0.350 0.510 0.800 ;
        RECT  0.420 0.870 0.490 1.055 ;
        RECT  0.130 0.870 0.420 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D1BWP

MACRO XOR4D2BWP
    CLASS CORE ;
    FOREIGN XOR4D2BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.770 ;
        RECT  2.530 0.355 2.555 0.475 ;
        RECT  2.470 0.650 2.555 0.770 ;
        RECT  2.460 0.195 2.530 0.475 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.010 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.520 2.790 0.640 ;
        RECT  2.695 0.355 2.765 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0336 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.495 3.605 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.780 0.115 ;
        RECT  3.520 -0.115 3.590 0.425 ;
        RECT  2.720 -0.115 3.520 0.115 ;
        RECT  3.430 0.355 3.520 0.425 ;
        RECT  2.640 -0.115 2.720 0.275 ;
        RECT  2.350 -0.115 2.640 0.115 ;
        RECT  2.270 -0.115 2.350 0.290 ;
        RECT  1.480 -0.115 2.270 0.115 ;
        RECT  1.410 -0.115 1.480 0.460 ;
        RECT  1.140 -0.115 1.410 0.115 ;
        RECT  1.040 -0.115 1.140 0.275 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.145 3.780 1.375 ;
        RECT  3.450 1.010 3.570 1.375 ;
        RECT  2.370 1.145 3.450 1.375 ;
        RECT  2.290 0.980 2.370 1.375 ;
        RECT  1.540 1.145 2.290 1.375 ;
        RECT  1.420 0.985 1.540 1.375 ;
        RECT  0.330 1.145 1.420 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.300 3.745 1.050 ;
        RECT  3.660 0.300 3.675 0.440 ;
        RECT  3.650 0.870 3.675 1.050 ;
        RECT  3.305 0.870 3.650 0.940 ;
        RECT  2.950 0.200 3.450 0.270 ;
        RECT  3.270 0.345 3.350 0.800 ;
        RECT  3.235 0.870 3.305 1.055 ;
        RECT  3.160 0.985 3.235 1.055 ;
        RECT  3.090 0.700 3.145 0.830 ;
        RECT  3.020 0.350 3.090 1.050 ;
        RECT  2.520 0.980 3.020 1.050 ;
        RECT  2.880 0.200 2.950 0.910 ;
        RECT  2.835 0.300 2.880 0.420 ;
        RECT  2.810 0.840 2.880 0.910 ;
        RECT  2.450 0.840 2.520 1.050 ;
        RECT  2.390 0.840 2.450 0.910 ;
        RECT  2.320 0.370 2.390 0.910 ;
        RECT  2.190 0.370 2.320 0.440 ;
        RECT  2.180 0.730 2.320 0.800 ;
        RECT  2.040 0.520 2.250 0.640 ;
        RECT  2.120 0.210 2.190 0.440 ;
        RECT  2.110 0.730 2.180 1.050 ;
        RECT  1.620 0.210 2.120 0.280 ;
        RECT  1.970 0.360 2.040 1.055 ;
        RECT  1.850 0.360 1.970 0.440 ;
        RECT  1.850 0.985 1.970 1.055 ;
        RECT  1.830 0.520 1.900 0.915 ;
        RECT  1.310 0.845 1.830 0.915 ;
        RECT  1.690 0.360 1.760 0.775 ;
        RECT  1.610 0.700 1.690 0.775 ;
        RECT  1.550 0.210 1.620 0.620 ;
        RECT  1.480 0.540 1.550 0.620 ;
        RECT  1.220 0.995 1.340 1.075 ;
        RECT  1.230 0.185 1.310 0.915 ;
        RECT  0.780 0.995 1.220 1.065 ;
        RECT  1.080 0.345 1.150 0.915 ;
        RECT  0.950 0.345 1.080 0.415 ;
        RECT  0.850 0.845 1.080 0.915 ;
        RECT  0.870 0.200 0.950 0.415 ;
        RECT  0.330 0.200 0.870 0.270 ;
        RECT  0.710 0.350 0.780 1.065 ;
        RECT  0.690 0.350 0.710 0.830 ;
        RECT  0.645 0.700 0.690 0.830 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.430 0.350 0.510 0.800 ;
        RECT  0.420 0.870 0.490 1.055 ;
        RECT  0.130 0.870 0.420 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D2BWP

MACRO XOR4D4BWP
    CLASS CORE ;
    FOREIGN XOR4D4BWP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.2016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.985 0.485 ;
        RECT  2.915 0.775 2.985 1.055 ;
        RECT  2.835 0.775 2.915 0.905 ;
        RECT  2.625 0.355 2.835 0.905 ;
        RECT  2.535 0.355 2.625 0.480 ;
        RECT  2.605 0.775 2.625 0.905 ;
        RECT  2.535 0.775 2.605 1.055 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0332 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0288 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.495 1.090 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0576 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.495 3.475 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0344 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.360 0.495 4.445 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 -0.115 4.620 0.115 ;
        RECT  4.300 -0.115 4.400 0.315 ;
        RECT  1.140 -0.115 4.300 0.115 ;
        RECT  1.040 -0.115 1.140 0.420 ;
        RECT  0.260 -0.115 1.040 0.115 ;
        RECT  0.260 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 1.145 4.620 1.375 ;
        RECT  4.310 0.985 4.380 1.375 ;
        RECT  3.530 1.145 4.310 1.375 ;
        RECT  3.450 0.985 3.530 1.375 ;
        RECT  3.170 1.145 3.450 1.375 ;
        RECT  3.090 0.665 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.710 0.985 2.810 1.375 ;
        RECT  2.090 1.145 2.710 1.375 ;
        RECT  1.970 1.010 2.090 1.375 ;
        RECT  0.330 1.145 1.970 1.375 ;
        RECT  0.210 1.010 0.330 1.375 ;
        RECT  0.000 1.145 0.210 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.355 2.985 0.485 ;
        RECT  2.915 0.775 2.985 1.055 ;
        RECT  2.905 0.775 2.915 0.905 ;
        RECT  2.535 0.355 2.555 0.480 ;
        RECT  2.535 0.775 2.555 1.055 ;
        RECT  4.515 0.195 4.585 1.005 ;
        RECT  4.490 0.195 4.515 0.355 ;
        RECT  4.490 0.845 4.515 1.005 ;
        RECT  4.020 0.845 4.490 0.915 ;
        RECT  3.720 0.990 4.230 1.060 ;
        RECT  4.140 0.375 4.210 0.755 ;
        RECT  4.030 0.375 4.140 0.445 ;
        RECT  4.090 0.685 4.140 0.755 ;
        RECT  3.950 0.540 4.020 0.915 ;
        RECT  3.880 0.210 3.970 0.315 ;
        RECT  3.810 0.210 3.880 0.910 ;
        RECT  2.065 0.210 3.810 0.280 ;
        RECT  3.635 0.350 3.720 1.060 ;
        RECT  3.230 0.350 3.635 0.420 ;
        RECT  3.250 0.845 3.635 0.915 ;
        RECT  2.450 0.550 2.530 0.620 ;
        RECT  2.380 0.550 2.450 0.940 ;
        RECT  1.690 0.870 2.380 0.940 ;
        RECT  2.175 0.350 2.270 0.800 ;
        RECT  1.865 0.730 2.175 0.800 ;
        RECT  1.985 0.210 2.065 0.660 ;
        RECT  1.520 0.210 1.985 0.280 ;
        RECT  1.790 0.350 1.865 0.800 ;
        RECT  1.610 0.350 1.690 1.040 ;
        RECT  1.450 0.210 1.520 0.905 ;
        RECT  1.370 0.210 1.450 0.300 ;
        RECT  1.390 0.835 1.450 0.905 ;
        RECT  1.310 0.530 1.380 0.650 ;
        RECT  0.780 0.980 1.325 1.050 ;
        RECT  1.235 0.350 1.310 0.880 ;
        RECT  0.920 0.840 0.990 0.910 ;
        RECT  0.920 0.310 0.960 0.410 ;
        RECT  0.850 0.200 0.920 0.910 ;
        RECT  0.340 0.200 0.850 0.270 ;
        RECT  0.710 0.350 0.780 1.050 ;
        RECT  0.690 0.350 0.710 0.910 ;
        RECT  0.630 0.840 0.690 0.910 ;
        RECT  0.550 0.990 0.640 1.060 ;
        RECT  0.480 0.870 0.550 1.060 ;
        RECT  0.465 0.350 0.540 0.800 ;
        RECT  0.130 0.870 0.480 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D4BWP

END LIBRARY
