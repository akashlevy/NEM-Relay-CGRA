VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MANUFACTURINGGRID 0.005 ;

MACRO nem_ohmux_invd0_4i_8b
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN nem_ohmux_invd0_4i_8b 0 0 ;
  SIZE 16.4 BY 4.38 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN I0_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.34 2.87 2.51 3.04 ;
    END
  END I0_0
  PIN I0_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.95 2.71 2.12 2.88 ;
    END
  END I0_7
  PIN I0_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.045 2.56 3.215 2.73 ;
    END
  END I0_1
  PIN I0_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.195 2.23 3.365 2.4 ;
    END
  END I0_2
  PIN I0_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.95 1.535 3.12 1.705 ;
    END
  END I0_3
  PIN I0_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.575 1.38 2.745 1.55 ;
    END
  END I0_4
  PIN I0_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.84 1.655 2.01 1.825 ;
    END
  END I0_5
  PIN I0_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.685 1.995 1.855 2.165 ;
    END
  END I0_6
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.365 2.095 2.535 2.265 ;
    END
  END S0
  PIN ZN_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.96 1.265 7.105 1.345 ;
        RECT 7.035 0.515 7.105 1.345 ;
        RECT 6.96 0.515 7.105 0.595 ;
    END
  END ZN_3
  PIN ZN_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.54 1.265 6.685 1.345 ;
        RECT 6.615 0.515 6.685 1.345 ;
        RECT 6.54 0.515 6.685 0.595 ;
    END
  END ZN_6
  PIN ZN_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.12 1.265 6.265 1.345 ;
        RECT 6.195 0.515 6.265 1.345 ;
        RECT 6.12 0.515 6.265 0.595 ;
    END
  END ZN_4
  PIN ZN_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7 1.265 5.845 1.345 ;
        RECT 5.775 0.515 5.845 1.345 ;
        RECT 5.7 0.515 5.845 0.595 ;
    END
  END ZN_5
  PIN ZN_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.96 3.785 7.105 3.865 ;
        RECT 7.035 3.035 7.105 3.865 ;
        RECT 6.96 3.035 7.105 3.115 ;
    END
  END ZN_1
  PIN ZN_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.54 3.785 6.685 3.865 ;
        RECT 6.615 3.035 6.685 3.865 ;
        RECT 6.54 3.035 6.685 3.115 ;
    END
  END ZN_2
  PIN ZN_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.12 3.785 6.265 3.865 ;
        RECT 6.195 3.035 6.265 3.865 ;
        RECT 6.12 3.035 6.265 3.115 ;
    END
  END ZN_0
  PIN ZN_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.7 3.785 5.845 3.865 ;
        RECT 5.775 3.035 5.845 3.865 ;
        RECT 5.7 3.035 5.845 3.115 ;
    END
  END ZN_7
  PIN I3_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.915 1.38 14.085 1.55 ;
    END
  END I3_4
  PIN I1_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.675 2.515 5.845 2.685 ;
    END
  END I1_7
  PIN I3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.385 2.56 14.555 2.73 ;
    END
  END I3_1
  PIN I3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.68 2.87 13.85 3.04 ;
    END
  END I3_0
  PIN I3_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.29 1.535 14.46 1.705 ;
    END
  END I3_3
  PIN I3_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.18 1.655 13.35 1.825 ;
    END
  END I3_5
  PIN I3_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.535 2.23 14.705 2.4 ;
    END
  END I3_2
  PIN I3_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.025 1.995 13.195 2.165 ;
    END
  END I3_6
  PIN S3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.705 2.095 13.875 2.265 ;
    END
  END S3
  PIN VSNEM
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M8 ;
        RECT 0 0 1.28 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 3.78 0 5.06 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 7.56 0 8.84 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 11.34 0 12.62 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 15.12 0 16.4 4.38 ;
    END
  END VSNEM
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 5.46 2.705 7.14 2.935 ;
        RECT 6.8 2.705 6.88 3.145 ;
        RECT 6.38 2.705 6.46 3.145 ;
        RECT 5.96 2.705 6.04 3.145 ;
        RECT 5.54 2.705 5.62 3.145 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.46 0.185 7.14 0.415 ;
        RECT 6.8 0.185 6.88 0.625 ;
        RECT 6.38 0.185 6.46 0.625 ;
        RECT 5.96 0.185 6.04 0.625 ;
        RECT 5.54 0.185 5.62 0.625 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 5.46 3.965 7.14 4.195 ;
        RECT 6.8 3.755 6.88 4.195 ;
        RECT 6.38 3.755 6.46 4.195 ;
        RECT 5.96 3.755 6.04 4.195 ;
        RECT 5.54 3.755 5.62 4.195 ;
    END
    PORT
      LAYER M1 ;
        RECT 5.46 1.445 7.14 1.675 ;
        RECT 6.8 1.235 6.88 1.675 ;
        RECT 6.38 1.235 6.46 1.675 ;
        RECT 5.96 1.235 6.04 1.675 ;
        RECT 5.54 1.235 5.62 1.675 ;
    END
  END VDD
  PIN S2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.925 2.095 10.095 2.265 ;
    END
  END S2
  PIN I2_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.755 2.23 10.925 2.4 ;
    END
  END I2_2
  PIN I2_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.135 1.38 10.305 1.55 ;
    END
  END I2_4
  PIN I2_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.51 1.535 10.68 1.705 ;
    END
  END I2_3
  PIN I2_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.245 1.995 9.415 2.165 ;
    END
  END I2_6
  PIN I2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.605 2.56 10.775 2.73 ;
    END
  END I2_1
  PIN I2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.9 2.87 10.07 3.04 ;
    END
  END I2_0
  PIN I2_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.4 1.655 9.57 1.825 ;
    END
  END I2_5
  PIN I2_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.51 2.71 9.68 2.88 ;
    END
  END I2_7
  PIN I3_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.29 2.71 13.46 2.88 ;
    END
  END I3_7
  PIN I1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.075 2.87 6.245 3.04 ;
    END
  END I1_0
  PIN I1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.825 2.56 6.995 2.73 ;
    END
  END I1_1
  PIN I1_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.975 2.23 7.145 2.4 ;
    END
  END I1_2
  PIN I1_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.73 1.535 6.9 1.705 ;
    END
  END I1_3
  PIN I1_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.355 1.385 6.525 1.555 ;
    END
  END I1_4
  PIN I1_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.62 1.655 5.79 1.825 ;
    END
  END I1_5
  PIN I1_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.465 1.995 5.635 2.165 ;
    END
  END I1_6
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.145 2.095 6.315 2.265 ;
    END
  END S1
  OBS
    LAYER OVERLAP ;
      RECT 0 0 16.4 4.38 ;
    LAYER M1 ;
      RECT 6.755 0.795 6.825 1.065 ;
      RECT 6.755 0.845 6.96 0.915 ;
      RECT 6.755 3.315 6.825 3.585 ;
      RECT 6.755 3.365 6.96 3.435 ;
      RECT 6.335 0.795 6.405 1.065 ;
      RECT 6.335 0.845 6.54 0.915 ;
      RECT 6.335 3.315 6.405 3.585 ;
      RECT 6.335 3.365 6.54 3.435 ;
      RECT 5.915 0.795 5.985 1.065 ;
      RECT 5.915 0.845 6.12 0.915 ;
      RECT 5.915 3.315 5.985 3.585 ;
      RECT 5.915 3.365 6.12 3.435 ;
      RECT 5.495 0.795 5.565 1.065 ;
      RECT 5.495 0.845 5.7 0.915 ;
      RECT 5.495 3.315 5.565 3.585 ;
      RECT 5.495 3.365 5.7 3.435 ;
    LAYER M2 ;
      RECT 6.755 0.675 6.825 1.065 ;
      RECT 6.755 3.195 6.825 3.585 ;
      RECT 6.335 0.675 6.405 1.065 ;
      RECT 6.335 3.195 6.405 3.585 ;
      RECT 5.915 0.675 5.985 1.065 ;
      RECT 5.915 3.195 5.985 3.585 ;
      RECT 5.495 0.675 5.565 1.065 ;
      RECT 5.495 3.195 5.565 3.585 ;
    LAYER M3 ;
      RECT 6.755 0.675 6.825 1.065 ;
      RECT 6.755 3.195 6.825 3.585 ;
      RECT 6.335 0.675 6.405 1.065 ;
      RECT 6.335 3.195 6.405 3.585 ;
      RECT 5.915 0.675 5.985 1.065 ;
      RECT 5.915 3.195 5.985 3.585 ;
      RECT 5.495 0.675 5.565 1.065 ;
      RECT 5.495 3.195 5.565 3.585 ;
    LAYER M4 ;
      RECT 6.755 0.675 6.825 1.065 ;
      RECT 6.755 3.195 6.825 3.585 ;
      RECT 6.335 0.675 6.405 1.065 ;
      RECT 6.335 3.195 6.405 3.585 ;
      RECT 5.915 0.675 5.985 1.065 ;
      RECT 5.915 3.195 5.985 3.585 ;
      RECT 5.495 0.675 5.565 1.065 ;
      RECT 5.495 3.195 5.565 3.585 ;
    LAYER M5 ;
      RECT 6.755 0.675 6.825 1.065 ;
      RECT 6.755 3.195 6.825 3.585 ;
      RECT 6.335 0.675 6.405 1.065 ;
      RECT 6.335 3.195 6.405 3.585 ;
      RECT 5.915 0.675 5.985 1.065 ;
      RECT 5.915 3.195 5.985 3.585 ;
      RECT 5.495 0.675 5.565 1.065 ;
      RECT 5.495 3.195 5.565 3.585 ;
    LAYER M6 ;
      RECT 6.755 0.795 6.825 1.475 ;
      RECT 6.755 2.87 6.825 3.585 ;
      RECT 6.335 0.795 6.405 1.325 ;
      RECT 6.335 2.87 6.405 3.585 ;
      RECT 5.915 0.795 5.985 1.585 ;
      RECT 5.915 2.87 5.985 3.585 ;
      RECT 5.495 0.795 5.565 1.585 ;
      RECT 5.495 2.87 5.565 3.585 ;
    LAYER M7 ;
      RECT 6.725 1.215 6.86 1.455 ;
      RECT 6.75 2.8 6.83 3.14 ;
      RECT 6.235 1.21 6.5 1.315 ;
      RECT 6.335 2.75 6.405 3.14 ;
      RECT 5.91 1.245 5.99 1.585 ;
      RECT 5.915 2.75 5.985 3.14 ;
      RECT 5.49 1.245 5.57 1.585 ;
      RECT 5.495 2.75 5.565 3.14 ;
    LAYER M8 ;
      RECT 14.765 3.335 14.895 3.465 ;
      RECT 14.795 2.15 14.865 3.465 ;
      RECT 14.765 2.15 14.895 2.28 ;
      RECT 14.58 1.37 14.71 1.5 ;
      RECT 14.61 0.505 14.68 1.5 ;
      RECT 14.58 0.505 14.71 0.635 ;
      RECT 14.555 3.735 14.685 3.865 ;
      RECT 14.585 2.885 14.655 3.865 ;
      RECT 14.555 2.885 14.685 3.015 ;
      RECT 13.08 3.535 13.21 3.665 ;
      RECT 13.11 2.87 13.18 3.665 ;
      RECT 13.04 2.87 13.18 3 ;
      RECT 13.05 1.38 13.18 1.51 ;
      RECT 13.08 0.705 13.15 1.51 ;
      RECT 13.05 0.705 13.18 0.835 ;
      RECT 12.835 2.11 12.965 2.24 ;
      RECT 12.865 0.905 12.935 2.24 ;
      RECT 12.835 0.905 12.965 1.035 ;
      RECT 10.985 3.335 11.115 3.465 ;
      RECT 11.015 2.15 11.085 3.465 ;
      RECT 10.985 2.15 11.115 2.28 ;
      RECT 10.8 1.37 10.93 1.5 ;
      RECT 10.83 0.505 10.9 1.5 ;
      RECT 10.8 0.505 10.93 0.635 ;
      RECT 10.775 3.735 10.905 3.865 ;
      RECT 10.805 2.885 10.875 3.865 ;
      RECT 10.775 2.885 10.905 3.015 ;
      RECT 9.3 3.535 9.43 3.665 ;
      RECT 9.33 2.87 9.4 3.665 ;
      RECT 9.26 2.87 9.4 3 ;
      RECT 9.27 1.38 9.4 1.51 ;
      RECT 9.3 0.705 9.37 1.51 ;
      RECT 9.27 0.705 9.4 0.835 ;
      RECT 9.055 2.11 9.185 2.24 ;
      RECT 9.085 0.905 9.155 2.24 ;
      RECT 9.055 0.905 9.185 1.035 ;
      RECT 7.205 3.335 7.335 3.465 ;
      RECT 7.235 2.15 7.305 3.465 ;
      RECT 7.205 2.15 7.335 2.28 ;
      RECT 7.02 1.37 7.15 1.5 ;
      RECT 7.05 0.505 7.12 1.5 ;
      RECT 7.02 0.505 7.15 0.635 ;
      RECT 6.995 3.735 7.125 3.865 ;
      RECT 7.025 2.885 7.095 3.865 ;
      RECT 6.995 2.885 7.125 3.015 ;
      RECT 6.755 0.505 6.825 1.465 ;
      RECT 6.725 0.505 6.855 0.635 ;
      RECT 6.725 3.735 6.855 3.865 ;
      RECT 6.755 2.87 6.825 3.865 ;
      RECT 6.335 0.905 6.405 1.315 ;
      RECT 6.305 0.905 6.435 1.035 ;
      RECT 6.305 3.335 6.435 3.465 ;
      RECT 6.335 2.87 6.405 3.465 ;
      RECT 5.915 1.105 5.985 1.515 ;
      RECT 5.885 1.105 6.015 1.235 ;
      RECT 5.885 3.135 6.015 3.265 ;
      RECT 5.915 2.87 5.985 3.265 ;
      RECT 5.465 3.535 5.595 3.665 ;
      RECT 5.495 2.87 5.565 3.665 ;
      RECT 5.495 2.87 5.625 3 ;
      RECT 5.47 1.38 5.6 1.51 ;
      RECT 5.495 0.705 5.565 1.51 ;
      RECT 5.465 0.705 5.595 0.835 ;
      RECT 5.275 2.11 5.405 2.24 ;
      RECT 5.305 0.905 5.375 2.24 ;
      RECT 5.275 0.905 5.405 1.035 ;
      RECT 3.425 3.335 3.555 3.465 ;
      RECT 3.455 2.15 3.525 3.465 ;
      RECT 3.425 2.15 3.555 2.28 ;
      RECT 3.24 1.37 3.37 1.5 ;
      RECT 3.27 0.505 3.34 1.5 ;
      RECT 3.24 0.505 3.37 0.635 ;
      RECT 3.215 3.735 3.345 3.865 ;
      RECT 3.245 2.885 3.315 3.865 ;
      RECT 3.215 2.885 3.345 3.015 ;
      RECT 1.74 3.535 1.87 3.665 ;
      RECT 1.77 2.87 1.84 3.665 ;
      RECT 1.7 2.87 1.84 3 ;
      RECT 1.71 1.38 1.84 1.51 ;
      RECT 1.74 0.705 1.81 1.51 ;
      RECT 1.71 0.705 1.84 0.835 ;
      RECT 1.495 2.11 1.625 2.24 ;
      RECT 1.525 0.905 1.595 2.24 ;
      RECT 1.495 0.905 1.625 1.035 ;
      RECT 14.525 2.225 14.695 2.395 ;
      RECT 14.385 2.565 14.555 2.735 ;
      RECT 14.29 1.535 14.46 1.705 ;
      RECT 13.9 1.385 14.07 1.555 ;
      RECT 13.705 2.09 13.875 2.26 ;
      RECT 13.68 2.87 13.85 3.04 ;
      RECT 13.29 2.71 13.46 2.88 ;
      RECT 13.18 1.635 13.35 1.805 ;
      RECT 13.035 1.99 13.205 2.16 ;
      RECT 10.745 2.225 10.915 2.395 ;
      RECT 10.605 2.565 10.775 2.735 ;
      RECT 10.51 1.535 10.68 1.705 ;
      RECT 10.12 1.385 10.29 1.555 ;
      RECT 9.925 2.09 10.095 2.26 ;
      RECT 9.9 2.87 10.07 3.04 ;
      RECT 9.51 2.71 9.68 2.88 ;
      RECT 9.4 1.635 9.57 1.805 ;
      RECT 9.255 1.99 9.425 2.16 ;
      RECT 6.965 2.225 7.135 2.395 ;
      RECT 6.825 2.565 6.995 2.735 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 6.075 2.87 6.245 3.04 ;
      RECT 5.745 2.535 5.87 2.79 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 3.185 2.225 3.355 2.395 ;
      RECT 3.045 2.565 3.215 2.735 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 2.34 2.87 2.51 3.04 ;
      RECT 1.95 2.71 2.12 2.88 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.695 1.99 1.865 2.16 ;
    LAYER M9 ;
      RECT 6.12 2.87 6.29 3.04 ;
      RECT 6.115 2.87 6.29 3 ;
      RECT 15.61 0.165 15.91 0.435 ;
      RECT 15.61 3.945 15.91 4.215 ;
      RECT 14.765 2.15 15 2.28 ;
      RECT 1.495 0.505 14.895 0.635 ;
      RECT 1.495 0.705 14.895 0.835 ;
      RECT 1.495 0.905 14.895 1.035 ;
      RECT 1.495 1.105 14.895 1.235 ;
      RECT 1.495 3.135 14.895 3.265 ;
      RECT 1.495 3.335 14.895 3.465 ;
      RECT 1.495 3.535 14.895 3.665 ;
      RECT 1.495 3.735 14.895 3.865 ;
      RECT 14.56 1.35 14.73 1.52 ;
      RECT 14.535 2.865 14.705 3.035 ;
      RECT 14.525 2.225 14.695 2.395 ;
      RECT 14.385 2.565 14.555 2.735 ;
      RECT 14.29 1.535 14.46 1.705 ;
      RECT 13.9 1.385 14.07 1.555 ;
      RECT 13.705 2.09 13.875 2.26 ;
      RECT 13.68 2.87 13.85 3.04 ;
      RECT 13.29 2.71 13.46 2.88 ;
      RECT 13.18 1.635 13.35 1.805 ;
      RECT 13.035 1.99 13.205 2.16 ;
      RECT 13.03 1.36 13.2 1.53 ;
      RECT 13.02 2.85 13.19 3.02 ;
      RECT 12.75 2.11 12.965 2.24 ;
      RECT 11.83 0.165 12.13 0.435 ;
      RECT 11.83 3.945 12.13 4.215 ;
      RECT 10.985 2.15 11.22 2.28 ;
      RECT 10.78 1.35 10.95 1.52 ;
      RECT 10.755 2.865 10.925 3.035 ;
      RECT 10.745 2.225 10.915 2.395 ;
      RECT 10.605 2.565 10.775 2.735 ;
      RECT 10.51 1.535 10.68 1.705 ;
      RECT 10.12 1.385 10.29 1.555 ;
      RECT 9.925 2.09 10.095 2.26 ;
      RECT 9.9 2.87 10.07 3.04 ;
      RECT 9.51 2.71 9.68 2.88 ;
      RECT 9.4 1.635 9.57 1.805 ;
      RECT 9.255 1.99 9.425 2.16 ;
      RECT 9.25 1.36 9.42 1.53 ;
      RECT 9.24 2.85 9.41 3.02 ;
      RECT 8.97 2.11 9.185 2.24 ;
      RECT 8.05 0.165 8.35 0.435 ;
      RECT 8.05 3.945 8.35 4.215 ;
      RECT 7.205 2.15 7.44 2.28 ;
      RECT 7 1.35 7.17 1.52 ;
      RECT 6.975 2.865 7.145 3.035 ;
      RECT 6.965 2.225 7.135 2.395 ;
      RECT 6.825 2.565 6.995 2.735 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 5.735 2.69 5.905 2.86 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 5.475 2.85 5.645 3.02 ;
      RECT 5.45 1.36 5.62 1.53 ;
      RECT 5.19 2.11 5.405 2.24 ;
      RECT 4.27 0.165 4.57 0.435 ;
      RECT 4.27 3.945 4.57 4.215 ;
      RECT 3.425 2.15 3.66 2.28 ;
      RECT 3.22 1.35 3.39 1.52 ;
      RECT 3.195 2.865 3.365 3.035 ;
      RECT 3.185 2.225 3.355 2.395 ;
      RECT 3.045 2.565 3.215 2.735 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 2.34 2.87 2.51 3.04 ;
      RECT 1.95 2.71 2.12 2.88 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.695 1.99 1.865 2.16 ;
      RECT 1.69 1.36 1.86 1.53 ;
      RECT 1.68 2.85 1.85 3.02 ;
      RECT 1.41 2.11 1.625 2.24 ;
      RECT 0.49 0.165 0.79 0.435 ;
      RECT 0.49 3.945 0.79 4.215 ;
    LAYER M10 ;
      RECT 12.48 3.375 15.26 3.58 ;
      RECT 15.05 0.8 15.26 3.58 ;
      RECT 13.97 3.075 15.26 3.58 ;
      RECT 14.75 2.335 15.26 3.58 ;
      RECT 12.48 3.07 13.72 3.58 ;
      RECT 12.48 3.07 13.725 3.22 ;
      RECT 13.875 1.57 14.23 3.125 ;
      RECT 12.48 3.07 14.5 3.125 ;
      RECT 13.97 2.785 14.5 3.58 ;
      RECT 12.48 3.065 13.625 3.58 ;
      RECT 13.525 0.8 13.625 3.58 ;
      RECT 13.24 2.91 13.625 3.58 ;
      RECT 12.48 2.295 12.99 3.58 ;
      RECT 13.24 1.845 13.275 3.58 ;
      RECT 13.875 2.785 15.26 2.825 ;
      RECT 14.745 1.555 14.8 2.825 ;
      RECT 13.525 1.26 13.875 2.82 ;
      RECT 12.48 2.295 13.275 2.815 ;
      RECT 14.59 2.435 15.26 2.825 ;
      RECT 13.525 1.715 14.34 2.82 ;
      RECT 12.48 2.295 14.34 2.66 ;
      RECT 13.39 0.8 13.775 2.66 ;
      RECT 12.48 2.435 15.26 2.535 ;
      RECT 12.935 2.2 14.495 2.535 ;
      RECT 13.39 1.715 14.495 2.535 ;
      RECT 12.48 0.8 12.685 3.58 ;
      RECT 13.235 1.845 14.495 2.535 ;
      RECT 12.935 1.565 12.985 3.58 ;
      RECT 14.48 1.555 14.8 2.185 ;
      RECT 14.76 0.8 15.26 2.085 ;
      RECT 12.48 0.8 12.98 2.045 ;
      RECT 12.48 1.845 15.26 1.95 ;
      RECT 12.48 1.565 13.14 1.95 ;
      RECT 13.23 0.8 13.775 1.595 ;
      RECT 14.125 0.8 14.23 3.58 ;
      RECT 12.48 1.565 13.875 1.595 ;
      RECT 14.48 0.8 14.51 2.185 ;
      RECT 14.125 0.8 14.51 1.465 ;
      RECT 13.23 1.26 14.51 1.32 ;
      RECT 12.48 0.8 13.775 1.315 ;
      RECT 14.025 0.8 15.26 1.305 ;
      RECT 14.015 1.16 15.26 1.305 ;
      RECT 12.48 0.8 15.26 1.01 ;
      RECT 8.7 3.375 11.48 3.58 ;
      RECT 11.27 0.8 11.48 3.58 ;
      RECT 10.19 3.075 11.48 3.58 ;
      RECT 10.97 2.335 11.48 3.58 ;
      RECT 8.7 3.07 9.94 3.58 ;
      RECT 8.7 3.07 9.945 3.22 ;
      RECT 10.095 1.57 10.45 3.125 ;
      RECT 8.7 3.07 10.72 3.125 ;
      RECT 10.19 2.785 10.72 3.58 ;
      RECT 8.7 3.065 9.845 3.58 ;
      RECT 9.745 0.8 9.845 3.58 ;
      RECT 9.46 2.91 9.845 3.58 ;
      RECT 8.7 2.295 9.21 3.58 ;
      RECT 9.46 1.845 9.495 3.58 ;
      RECT 10.095 2.785 11.48 2.825 ;
      RECT 10.965 1.555 11.02 2.825 ;
      RECT 9.745 1.26 10.095 2.82 ;
      RECT 8.7 2.295 9.495 2.815 ;
      RECT 10.81 2.435 11.48 2.825 ;
      RECT 9.745 1.715 10.56 2.82 ;
      RECT 8.7 2.295 10.56 2.66 ;
      RECT 9.61 0.8 9.995 2.66 ;
      RECT 8.7 2.435 11.48 2.535 ;
      RECT 9.155 2.2 10.715 2.535 ;
      RECT 9.61 1.715 10.715 2.535 ;
      RECT 8.7 0.8 8.905 3.58 ;
      RECT 9.455 1.845 10.715 2.535 ;
      RECT 9.155 1.565 9.205 3.58 ;
      RECT 10.7 1.555 11.02 2.185 ;
      RECT 10.98 0.8 11.48 2.085 ;
      RECT 8.7 0.8 9.2 2.045 ;
      RECT 8.7 1.845 11.48 1.95 ;
      RECT 8.7 1.565 9.36 1.95 ;
      RECT 9.45 0.8 9.995 1.595 ;
      RECT 10.345 0.8 10.45 3.58 ;
      RECT 8.7 1.565 10.095 1.595 ;
      RECT 10.7 0.8 10.73 2.185 ;
      RECT 10.345 0.8 10.73 1.465 ;
      RECT 9.45 1.26 10.73 1.32 ;
      RECT 8.7 0.8 9.995 1.315 ;
      RECT 10.245 0.8 11.48 1.305 ;
      RECT 10.235 1.16 11.48 1.305 ;
      RECT 8.7 0.8 11.48 1.01 ;
      RECT 4.92 3.375 7.7 3.58 ;
      RECT 7.49 0.8 7.7 3.58 ;
      RECT 6.41 3.075 7.7 3.58 ;
      RECT 7.19 2.335 7.7 3.58 ;
      RECT 4.92 3.07 6.16 3.58 ;
      RECT 4.92 3.07 6.165 3.22 ;
      RECT 6.315 1.57 6.67 3.125 ;
      RECT 4.92 3.07 6.94 3.125 ;
      RECT 6.41 2.785 6.94 3.58 ;
      RECT 4.92 3.065 6.065 3.58 ;
      RECT 5.965 0.8 6.065 3.58 ;
      RECT 5.68 2.91 6.065 3.58 ;
      RECT 4.92 2.295 5.43 3.58 ;
      RECT 5.68 1.845 5.715 3.58 ;
      RECT 6.315 2.785 7.7 2.825 ;
      RECT 7.185 1.555 7.24 2.825 ;
      RECT 5.965 1.26 6.315 2.82 ;
      RECT 4.92 2.295 5.715 2.815 ;
      RECT 7.03 2.435 7.7 2.825 ;
      RECT 5.965 1.715 6.78 2.82 ;
      RECT 4.92 2.295 6.78 2.66 ;
      RECT 5.83 0.8 6.215 2.66 ;
      RECT 4.92 2.435 7.7 2.535 ;
      RECT 5.375 2.2 6.935 2.535 ;
      RECT 5.83 1.715 6.935 2.535 ;
      RECT 4.92 0.8 5.125 3.58 ;
      RECT 5.675 1.845 6.935 2.535 ;
      RECT 5.375 1.565 5.425 3.58 ;
      RECT 6.92 1.555 7.24 2.185 ;
      RECT 7.2 0.8 7.7 2.085 ;
      RECT 4.92 0.8 5.42 2.045 ;
      RECT 4.92 1.845 7.7 1.95 ;
      RECT 4.92 1.565 5.58 1.95 ;
      RECT 5.67 0.8 6.215 1.595 ;
      RECT 6.565 0.8 6.67 3.58 ;
      RECT 4.92 1.565 6.315 1.595 ;
      RECT 6.92 0.8 6.95 2.185 ;
      RECT 6.565 0.8 6.95 1.465 ;
      RECT 5.67 1.26 6.95 1.32 ;
      RECT 4.92 0.8 6.215 1.315 ;
      RECT 6.465 0.8 7.7 1.305 ;
      RECT 6.455 1.16 7.7 1.305 ;
      RECT 4.92 0.8 7.7 1.01 ;
      RECT 1.14 3.375 3.92 3.58 ;
      RECT 3.71 0.8 3.92 3.58 ;
      RECT 2.63 3.075 3.92 3.58 ;
      RECT 3.41 2.335 3.92 3.58 ;
      RECT 1.14 3.07 2.38 3.58 ;
      RECT 1.14 3.07 2.385 3.22 ;
      RECT 2.535 1.57 2.89 3.125 ;
      RECT 1.14 3.07 3.16 3.125 ;
      RECT 2.63 2.785 3.16 3.58 ;
      RECT 1.14 3.065 2.285 3.58 ;
      RECT 2.185 0.8 2.285 3.58 ;
      RECT 1.9 2.91 2.285 3.58 ;
      RECT 1.14 2.295 1.65 3.58 ;
      RECT 1.9 1.845 1.935 3.58 ;
      RECT 2.535 2.785 3.92 2.825 ;
      RECT 3.405 1.555 3.46 2.825 ;
      RECT 2.185 1.26 2.535 2.82 ;
      RECT 1.14 2.295 1.935 2.815 ;
      RECT 3.25 2.435 3.92 2.825 ;
      RECT 2.185 1.715 3 2.82 ;
      RECT 1.14 2.295 3 2.66 ;
      RECT 2.05 0.8 2.435 2.66 ;
      RECT 1.14 2.435 3.92 2.535 ;
      RECT 1.595 2.2 3.155 2.535 ;
      RECT 2.05 1.715 3.155 2.535 ;
      RECT 1.14 0.8 1.345 3.58 ;
      RECT 1.895 1.845 3.155 2.535 ;
      RECT 1.595 1.565 1.645 3.58 ;
      RECT 3.14 1.555 3.46 2.185 ;
      RECT 3.42 0.8 3.92 2.085 ;
      RECT 1.14 0.8 1.64 2.045 ;
      RECT 1.14 1.845 3.92 1.95 ;
      RECT 1.14 1.565 1.8 1.95 ;
      RECT 1.89 0.8 2.435 1.595 ;
      RECT 2.785 0.8 2.89 3.58 ;
      RECT 1.14 1.565 2.535 1.595 ;
      RECT 3.14 0.8 3.17 2.185 ;
      RECT 2.785 0.8 3.17 1.465 ;
      RECT 1.89 1.26 3.17 1.32 ;
      RECT 1.14 0.8 2.435 1.315 ;
      RECT 2.685 0.8 3.92 1.305 ;
      RECT 2.675 1.16 3.92 1.305 ;
      RECT 1.14 0.8 3.92 1.01 ;
      RECT 15.56 0.1 15.96 0.5 ;
      RECT 15.56 3.88 15.96 4.28 ;
      RECT 14.85 2.135 15 2.285 ;
      RECT 14.56 1.354 14.71 1.504 ;
      RECT 14.551 2.873 14.701 3.023 ;
      RECT 14.545 2.236 14.695 2.386 ;
      RECT 14.392 2.584 14.542 2.734 ;
      RECT 14.278 1.517 14.428 1.667 ;
      RECT 13.926 1.368 14.076 1.518 ;
      RECT 13.824 1.061 13.974 1.211 ;
      RECT 13.771 3.173 13.921 3.323 ;
      RECT 13.675 2.87 13.825 3.02 ;
      RECT 13.324 2.708 13.474 2.858 ;
      RECT 13.19 1.643 13.34 1.793 ;
      RECT 13.038 2.866 13.188 3.016 ;
      RECT 13.037 1.998 13.187 2.148 ;
      RECT 13.03 1.363 13.18 1.513 ;
      RECT 12.733 2.096 12.883 2.246 ;
      RECT 11.78 0.1 12.18 0.5 ;
      RECT 11.78 3.88 12.18 4.28 ;
      RECT 11.07 2.135 11.22 2.285 ;
      RECT 10.78 1.354 10.93 1.504 ;
      RECT 10.771 2.873 10.921 3.023 ;
      RECT 10.765 2.236 10.915 2.386 ;
      RECT 10.612 2.584 10.762 2.734 ;
      RECT 10.498 1.517 10.648 1.667 ;
      RECT 10.146 1.368 10.296 1.518 ;
      RECT 10.044 1.061 10.194 1.211 ;
      RECT 9.991 3.173 10.141 3.323 ;
      RECT 9.895 2.87 10.045 3.02 ;
      RECT 9.544 2.708 9.694 2.858 ;
      RECT 9.41 1.643 9.56 1.793 ;
      RECT 9.258 2.866 9.408 3.016 ;
      RECT 9.257 1.998 9.407 2.148 ;
      RECT 9.25 1.363 9.4 1.513 ;
      RECT 8.953 2.096 9.103 2.246 ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 7.29 2.135 7.44 2.285 ;
      RECT 7 1.354 7.15 1.504 ;
      RECT 6.991 2.873 7.141 3.023 ;
      RECT 6.985 2.236 7.135 2.386 ;
      RECT 6.832 2.584 6.982 2.734 ;
      RECT 6.718 1.517 6.868 1.667 ;
      RECT 6.366 1.368 6.516 1.518 ;
      RECT 6.264 1.061 6.414 1.211 ;
      RECT 6.211 3.173 6.361 3.323 ;
      RECT 6.115 2.87 6.265 3.02 ;
      RECT 5.764 2.708 5.914 2.858 ;
      RECT 5.63 1.643 5.78 1.793 ;
      RECT 5.478 2.866 5.628 3.016 ;
      RECT 5.477 1.998 5.627 2.148 ;
      RECT 5.47 1.363 5.62 1.513 ;
      RECT 5.173 2.096 5.323 2.246 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 3.51 2.135 3.66 2.285 ;
      RECT 3.22 1.354 3.37 1.504 ;
      RECT 3.211 2.873 3.361 3.023 ;
      RECT 3.205 2.236 3.355 2.386 ;
      RECT 3.052 2.584 3.202 2.734 ;
      RECT 2.938 1.517 3.088 1.667 ;
      RECT 2.586 1.368 2.736 1.518 ;
      RECT 2.484 1.061 2.634 1.211 ;
      RECT 2.431 3.173 2.581 3.323 ;
      RECT 2.335 2.87 2.485 3.02 ;
      RECT 1.984 2.708 2.134 2.858 ;
      RECT 1.85 1.643 2 1.793 ;
      RECT 1.698 2.866 1.848 3.016 ;
      RECT 1.697 1.998 1.847 2.148 ;
      RECT 1.69 1.363 1.84 1.513 ;
      RECT 1.393 2.096 1.543 2.246 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
    LAYER NEMANC ;
      RECT 15.56 0.1 15.96 0.5 ;
      RECT 15.56 3.88 15.96 4.28 ;
      RECT 11.78 0.1 12.18 0.5 ;
      RECT 11.78 3.88 12.18 4.28 ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
    LAYER NEMCHAN ;
      RECT 14.635 2.22 14.715 2.37 ;
      RECT 14.635 2.22 14.755 2.355 ;
      RECT 14.635 2.22 14.795 2.34 ;
      RECT 14.635 2.22 14.835 2.325 ;
      RECT 14.875 2.14 14.9 2.305 ;
      RECT 14.595 2.23 14.9 2.3 ;
      RECT 14.715 2.195 14.94 2.29 ;
      RECT 14.595 2.26 14.95 2.285 ;
      RECT 14.675 2.205 14.94 2.29 ;
      RECT 14.755 2.18 14.9 2.305 ;
      RECT 14.835 2.155 14.875 2.315 ;
      RECT 14.795 2.165 14.9 2.305 ;
      RECT 14.56 2.705 14.6 2.975 ;
      RECT 14.52 2.78 14.64 2.95 ;
      RECT 14.52 2.855 14.68 2.93 ;
      RECT 14.52 2.895 14.69 2.915 ;
      RECT 14.48 2.645 14.52 2.88 ;
      RECT 14.44 2.665 14.56 2.805 ;
      RECT 14.4 2.685 14.56 2.735 ;
      RECT 14.48 2.65 14.56 2.88 ;
      RECT 14.395 1.465 14.435 1.64 ;
      RECT 14.355 1.49 14.435 1.625 ;
      RECT 14.355 1.49 14.475 1.62 ;
      RECT 14.355 1.49 14.515 1.595 ;
      RECT 14.315 1.51 14.555 1.565 ;
      RECT 14.555 1.375 14.595 1.55 ;
      RECT 14.555 1.395 14.635 1.525 ;
      RECT 14.395 1.465 14.67 1.51 ;
      RECT 14.435 1.445 14.635 1.525 ;
      RECT 14.515 1.4 14.555 1.57 ;
      RECT 14.475 1.42 14.635 1.525 ;
      RECT 13.95 1.115 13.97 1.46 ;
      RECT 13.95 1.175 14.01 1.445 ;
      RECT 13.91 1.295 14.05 1.435 ;
      RECT 13.91 1.39 14.07 1.425 ;
      RECT 13.87 1.14 13.97 1.345 ;
      RECT 13.83 1.15 13.97 1.22 ;
      RECT 13.91 1.125 13.97 1.435 ;
      RECT 13.8 2.92 13.82 3.26 ;
      RECT 13.8 2.98 13.86 3.25 ;
      RECT 13.76 3.1 13.9 3.24 ;
      RECT 13.76 3.195 13.92 3.23 ;
      RECT 13.72 2.945 13.82 3.16 ;
      RECT 13.68 2.955 13.82 3.035 ;
      RECT 13.76 2.93 13.82 3.24 ;
      RECT 13.155 2.82 13.195 2.99 ;
      RECT 13.115 2.84 13.195 2.975 ;
      RECT 13.115 2.84 13.235 2.97 ;
      RECT 13.115 2.84 13.315 2.93 ;
      RECT 13.075 2.865 13.315 2.915 ;
      RECT 13.075 2.865 13.355 2.905 ;
      RECT 13.355 2.72 13.365 2.895 ;
      RECT 13.275 2.755 13.405 2.88 ;
      RECT 13.155 2.82 13.435 2.86 ;
      RECT 13.195 2.8 13.405 2.88 ;
      RECT 13.235 2.78 13.275 2.95 ;
      RECT 13.315 2.735 13.365 2.895 ;
      RECT 13.2 1.48 13.24 1.745 ;
      RECT 13.16 1.555 13.28 1.72 ;
      RECT 13.16 1.625 13.32 1.7 ;
      RECT 13.16 1.665 13.33 1.685 ;
      RECT 13.12 1.415 13.16 1.65 ;
      RECT 13.08 1.44 13.2 1.58 ;
      RECT 13.04 1.46 13.2 1.51 ;
      RECT 13.12 1.425 13.2 1.65 ;
      RECT 12.825 2.08 12.865 2.23 ;
      RECT 12.825 2.08 12.905 2.225 ;
      RECT 12.825 2.08 12.945 2.21 ;
      RECT 12.825 2.08 12.985 2.2 ;
      RECT 13.065 2 13.09 2.17 ;
      RECT 12.785 2.09 13.09 2.165 ;
      RECT 12.905 2.06 13.13 2.155 ;
      RECT 12.785 2.135 13.135 2.145 ;
      RECT 12.865 2.065 13.13 2.155 ;
      RECT 12.905 2.055 13.09 2.17 ;
      RECT 13.025 2.015 13.065 2.175 ;
      RECT 12.945 2.04 13.09 2.17 ;
      RECT 12.985 2.025 13.025 2.185 ;
      RECT 10.855 2.22 10.935 2.37 ;
      RECT 10.855 2.22 10.975 2.355 ;
      RECT 10.855 2.22 11.015 2.34 ;
      RECT 10.855 2.22 11.055 2.325 ;
      RECT 11.095 2.14 11.12 2.305 ;
      RECT 10.815 2.23 11.12 2.3 ;
      RECT 10.935 2.195 11.16 2.29 ;
      RECT 10.815 2.26 11.17 2.285 ;
      RECT 10.895 2.205 11.16 2.29 ;
      RECT 10.975 2.18 11.12 2.305 ;
      RECT 11.055 2.155 11.095 2.315 ;
      RECT 11.015 2.165 11.12 2.305 ;
      RECT 10.78 2.705 10.82 2.975 ;
      RECT 10.74 2.78 10.86 2.95 ;
      RECT 10.74 2.855 10.9 2.93 ;
      RECT 10.74 2.895 10.91 2.915 ;
      RECT 10.7 2.645 10.74 2.88 ;
      RECT 10.66 2.665 10.78 2.805 ;
      RECT 10.62 2.685 10.78 2.735 ;
      RECT 10.7 2.65 10.78 2.88 ;
      RECT 10.615 1.465 10.655 1.64 ;
      RECT 10.575 1.49 10.655 1.625 ;
      RECT 10.575 1.49 10.695 1.62 ;
      RECT 10.575 1.49 10.735 1.595 ;
      RECT 10.535 1.51 10.775 1.565 ;
      RECT 10.775 1.375 10.815 1.55 ;
      RECT 10.775 1.395 10.855 1.525 ;
      RECT 10.615 1.465 10.89 1.51 ;
      RECT 10.655 1.445 10.855 1.525 ;
      RECT 10.735 1.4 10.775 1.57 ;
      RECT 10.695 1.42 10.855 1.525 ;
      RECT 10.17 1.115 10.19 1.46 ;
      RECT 10.17 1.175 10.23 1.445 ;
      RECT 10.13 1.295 10.27 1.435 ;
      RECT 10.13 1.39 10.29 1.425 ;
      RECT 10.09 1.14 10.19 1.345 ;
      RECT 10.05 1.15 10.19 1.22 ;
      RECT 10.13 1.125 10.19 1.435 ;
      RECT 10.02 2.92 10.04 3.26 ;
      RECT 10.02 2.98 10.08 3.25 ;
      RECT 9.98 3.1 10.12 3.24 ;
      RECT 9.98 3.195 10.14 3.23 ;
      RECT 9.94 2.945 10.04 3.16 ;
      RECT 9.9 2.955 10.04 3.035 ;
      RECT 9.98 2.93 10.04 3.24 ;
      RECT 9.375 2.82 9.415 2.99 ;
      RECT 9.335 2.84 9.415 2.975 ;
      RECT 9.335 2.84 9.455 2.97 ;
      RECT 9.335 2.84 9.535 2.93 ;
      RECT 9.295 2.865 9.535 2.915 ;
      RECT 9.295 2.865 9.575 2.905 ;
      RECT 9.575 2.72 9.585 2.895 ;
      RECT 9.495 2.755 9.625 2.88 ;
      RECT 9.375 2.82 9.655 2.86 ;
      RECT 9.415 2.8 9.625 2.88 ;
      RECT 9.455 2.78 9.495 2.95 ;
      RECT 9.535 2.735 9.585 2.895 ;
      RECT 9.42 1.48 9.46 1.745 ;
      RECT 9.38 1.555 9.5 1.72 ;
      RECT 9.38 1.625 9.54 1.7 ;
      RECT 9.38 1.665 9.55 1.685 ;
      RECT 9.34 1.415 9.38 1.65 ;
      RECT 9.3 1.44 9.42 1.58 ;
      RECT 9.26 1.46 9.42 1.51 ;
      RECT 9.34 1.425 9.42 1.65 ;
      RECT 9.045 2.08 9.085 2.23 ;
      RECT 9.045 2.08 9.125 2.225 ;
      RECT 9.045 2.08 9.165 2.21 ;
      RECT 9.045 2.08 9.205 2.2 ;
      RECT 9.285 2 9.31 2.17 ;
      RECT 9.005 2.09 9.31 2.165 ;
      RECT 9.125 2.06 9.35 2.155 ;
      RECT 9.005 2.135 9.355 2.145 ;
      RECT 9.085 2.065 9.35 2.155 ;
      RECT 9.125 2.055 9.31 2.17 ;
      RECT 9.245 2.015 9.285 2.175 ;
      RECT 9.165 2.04 9.31 2.17 ;
      RECT 9.205 2.025 9.245 2.185 ;
      RECT 7.075 2.22 7.155 2.37 ;
      RECT 7.075 2.22 7.195 2.355 ;
      RECT 7.075 2.22 7.235 2.34 ;
      RECT 7.075 2.22 7.275 2.325 ;
      RECT 7.315 2.14 7.34 2.305 ;
      RECT 7.035 2.23 7.34 2.3 ;
      RECT 7.155 2.195 7.38 2.29 ;
      RECT 7.035 2.26 7.39 2.285 ;
      RECT 7.115 2.205 7.38 2.29 ;
      RECT 7.195 2.18 7.34 2.305 ;
      RECT 7.275 2.155 7.315 2.315 ;
      RECT 7.235 2.165 7.34 2.305 ;
      RECT 7 2.705 7.04 2.975 ;
      RECT 6.96 2.78 7.08 2.95 ;
      RECT 6.96 2.855 7.12 2.93 ;
      RECT 6.96 2.895 7.13 2.915 ;
      RECT 6.92 2.645 6.96 2.88 ;
      RECT 6.88 2.665 7 2.805 ;
      RECT 6.84 2.685 7 2.735 ;
      RECT 6.92 2.65 7 2.88 ;
      RECT 6.835 1.465 6.875 1.64 ;
      RECT 6.795 1.49 6.875 1.625 ;
      RECT 6.795 1.49 6.915 1.62 ;
      RECT 6.795 1.49 6.955 1.595 ;
      RECT 6.755 1.51 6.995 1.565 ;
      RECT 6.995 1.375 7.035 1.55 ;
      RECT 6.995 1.395 7.075 1.525 ;
      RECT 6.835 1.465 7.11 1.51 ;
      RECT 6.875 1.445 7.075 1.525 ;
      RECT 6.955 1.4 6.995 1.57 ;
      RECT 6.915 1.42 7.075 1.525 ;
      RECT 6.39 1.115 6.41 1.46 ;
      RECT 6.39 1.175 6.45 1.445 ;
      RECT 6.35 1.295 6.49 1.435 ;
      RECT 6.35 1.39 6.51 1.425 ;
      RECT 6.31 1.14 6.41 1.345 ;
      RECT 6.27 1.15 6.41 1.22 ;
      RECT 6.35 1.125 6.41 1.435 ;
      RECT 6.24 2.92 6.26 3.26 ;
      RECT 6.24 2.98 6.3 3.25 ;
      RECT 6.2 3.1 6.34 3.24 ;
      RECT 6.2 3.195 6.36 3.23 ;
      RECT 6.16 2.945 6.26 3.16 ;
      RECT 6.12 2.955 6.26 3.035 ;
      RECT 6.2 2.93 6.26 3.24 ;
      RECT 5.595 2.82 5.635 2.99 ;
      RECT 5.555 2.84 5.635 2.975 ;
      RECT 5.555 2.84 5.675 2.97 ;
      RECT 5.555 2.84 5.755 2.93 ;
      RECT 5.515 2.865 5.755 2.915 ;
      RECT 5.515 2.865 5.795 2.905 ;
      RECT 5.795 2.72 5.805 2.895 ;
      RECT 5.715 2.755 5.845 2.88 ;
      RECT 5.595 2.82 5.875 2.86 ;
      RECT 5.635 2.8 5.845 2.88 ;
      RECT 5.675 2.78 5.715 2.95 ;
      RECT 5.755 2.735 5.805 2.895 ;
      RECT 5.64 1.48 5.68 1.745 ;
      RECT 5.6 1.555 5.72 1.72 ;
      RECT 5.6 1.625 5.76 1.7 ;
      RECT 5.6 1.665 5.77 1.685 ;
      RECT 5.56 1.415 5.6 1.65 ;
      RECT 5.52 1.44 5.64 1.58 ;
      RECT 5.48 1.46 5.64 1.51 ;
      RECT 5.56 1.425 5.64 1.65 ;
      RECT 5.265 2.08 5.305 2.23 ;
      RECT 5.265 2.08 5.345 2.225 ;
      RECT 5.265 2.08 5.385 2.21 ;
      RECT 5.265 2.08 5.425 2.2 ;
      RECT 5.505 2 5.53 2.17 ;
      RECT 5.225 2.09 5.53 2.165 ;
      RECT 5.345 2.06 5.57 2.155 ;
      RECT 5.225 2.135 5.575 2.145 ;
      RECT 5.305 2.065 5.57 2.155 ;
      RECT 5.345 2.055 5.53 2.17 ;
      RECT 5.465 2.015 5.505 2.175 ;
      RECT 5.385 2.04 5.53 2.17 ;
      RECT 5.425 2.025 5.465 2.185 ;
      RECT 3.295 2.22 3.375 2.37 ;
      RECT 3.295 2.22 3.415 2.355 ;
      RECT 3.295 2.22 3.455 2.34 ;
      RECT 3.295 2.22 3.495 2.325 ;
      RECT 3.535 2.14 3.56 2.305 ;
      RECT 3.255 2.23 3.56 2.3 ;
      RECT 3.375 2.195 3.6 2.29 ;
      RECT 3.255 2.26 3.61 2.285 ;
      RECT 3.335 2.205 3.6 2.29 ;
      RECT 3.415 2.18 3.56 2.305 ;
      RECT 3.495 2.155 3.535 2.315 ;
      RECT 3.455 2.165 3.56 2.305 ;
      RECT 3.22 2.705 3.26 2.975 ;
      RECT 3.18 2.78 3.3 2.95 ;
      RECT 3.18 2.855 3.34 2.93 ;
      RECT 3.18 2.895 3.35 2.915 ;
      RECT 3.14 2.645 3.18 2.88 ;
      RECT 3.1 2.665 3.22 2.805 ;
      RECT 3.06 2.685 3.22 2.735 ;
      RECT 3.14 2.65 3.22 2.88 ;
      RECT 3.055 1.465 3.095 1.64 ;
      RECT 3.015 1.49 3.095 1.625 ;
      RECT 3.015 1.49 3.135 1.62 ;
      RECT 3.015 1.49 3.175 1.595 ;
      RECT 2.975 1.51 3.215 1.565 ;
      RECT 3.215 1.375 3.255 1.55 ;
      RECT 3.215 1.395 3.295 1.525 ;
      RECT 3.055 1.465 3.33 1.51 ;
      RECT 3.095 1.445 3.295 1.525 ;
      RECT 3.175 1.4 3.215 1.57 ;
      RECT 3.135 1.42 3.295 1.525 ;
      RECT 2.61 1.115 2.63 1.46 ;
      RECT 2.61 1.175 2.67 1.445 ;
      RECT 2.57 1.295 2.71 1.435 ;
      RECT 2.57 1.39 2.73 1.425 ;
      RECT 2.53 1.14 2.63 1.345 ;
      RECT 2.49 1.15 2.63 1.22 ;
      RECT 2.57 1.125 2.63 1.435 ;
      RECT 2.46 2.92 2.48 3.26 ;
      RECT 2.46 2.98 2.52 3.25 ;
      RECT 2.42 3.1 2.56 3.24 ;
      RECT 2.42 3.195 2.58 3.23 ;
      RECT 2.38 2.945 2.48 3.16 ;
      RECT 2.34 2.955 2.48 3.035 ;
      RECT 2.42 2.93 2.48 3.24 ;
      RECT 1.815 2.82 1.855 2.99 ;
      RECT 1.775 2.84 1.855 2.975 ;
      RECT 1.775 2.84 1.895 2.97 ;
      RECT 1.775 2.84 1.975 2.93 ;
      RECT 1.735 2.865 1.975 2.915 ;
      RECT 1.735 2.865 2.015 2.905 ;
      RECT 2.015 2.72 2.025 2.895 ;
      RECT 1.935 2.755 2.065 2.88 ;
      RECT 1.815 2.82 2.095 2.86 ;
      RECT 1.855 2.8 2.065 2.88 ;
      RECT 1.895 2.78 1.935 2.95 ;
      RECT 1.975 2.735 2.025 2.895 ;
      RECT 1.86 1.48 1.9 1.745 ;
      RECT 1.82 1.555 1.94 1.72 ;
      RECT 1.82 1.625 1.98 1.7 ;
      RECT 1.82 1.665 1.99 1.685 ;
      RECT 1.78 1.415 1.82 1.65 ;
      RECT 1.74 1.44 1.86 1.58 ;
      RECT 1.7 1.46 1.86 1.51 ;
      RECT 1.78 1.425 1.86 1.65 ;
      RECT 1.485 2.08 1.525 2.23 ;
      RECT 1.485 2.08 1.565 2.225 ;
      RECT 1.485 2.08 1.605 2.21 ;
      RECT 1.485 2.08 1.645 2.2 ;
      RECT 1.725 2 1.75 2.17 ;
      RECT 1.445 2.09 1.75 2.165 ;
      RECT 1.565 2.06 1.79 2.155 ;
      RECT 1.445 2.135 1.795 2.145 ;
      RECT 1.525 2.065 1.79 2.155 ;
      RECT 1.565 2.055 1.75 2.17 ;
      RECT 1.685 2.015 1.725 2.175 ;
      RECT 1.605 2.04 1.75 2.17 ;
      RECT 1.645 2.025 1.685 2.185 ;
    LAYER NEMBODY ;
      RECT 15.46 3.78 16.06 4.38 ;
      RECT 11.68 3.78 12.28 4.38 ;
      RECT 12.08 0.8 12.28 4.38 ;
      RECT 7.9 3.78 8.5 4.38 ;
      RECT 8.3 0.8 8.5 4.38 ;
      RECT 4.12 3.78 4.72 4.38 ;
      RECT 4.52 0.8 4.72 4.38 ;
      RECT 0.34 3.78 0.94 4.38 ;
      RECT 0.74 0.8 0.94 4.38 ;
      RECT 12.48 3.78 16.06 3.98 ;
      RECT 8.7 3.78 12.28 3.98 ;
      RECT 4.92 3.78 8.5 3.98 ;
      RECT 1.14 3.78 4.72 3.98 ;
      RECT 12.48 0.8 12.68 3.98 ;
      RECT 8.7 0.8 8.9 3.98 ;
      RECT 4.92 0.8 5.12 3.98 ;
      RECT 1.14 0.8 1.34 3.98 ;
      RECT 12.48 3.38 15.66 3.58 ;
      RECT 15.46 0 15.66 3.58 ;
      RECT 8.7 3.38 11.88 3.58 ;
      RECT 11.68 0 11.88 3.58 ;
      RECT 4.92 3.38 8.1 3.58 ;
      RECT 7.9 0 8.1 3.58 ;
      RECT 1.14 3.38 4.32 3.58 ;
      RECT 4.12 0 4.32 3.58 ;
      RECT 12.48 0.8 15.26 3.58 ;
      RECT 15.06 0.4 15.26 3.58 ;
      RECT 8.7 0.8 11.48 3.58 ;
      RECT 11.28 0.4 11.48 3.58 ;
      RECT 4.92 0.8 7.7 3.58 ;
      RECT 7.5 0.4 7.7 3.58 ;
      RECT 1.14 0.8 3.92 3.58 ;
      RECT 3.72 0.4 3.92 3.58 ;
      RECT 12.08 0.8 15.26 1 ;
      RECT 8.3 0.8 11.48 1 ;
      RECT 4.52 0.8 7.7 1 ;
      RECT 0.74 0.8 3.92 1 ;
      RECT 15.46 0 16.06 0.6 ;
      RECT 11.68 0.4 15.26 0.6 ;
      RECT 7.9 0.4 11.48 0.6 ;
      RECT 4.12 0.4 7.7 0.6 ;
      RECT 0.34 0.4 3.92 0.6 ;
      RECT 11.68 0 12.28 0.6 ;
      RECT 7.9 0 8.5 0.6 ;
      RECT 4.12 0 4.72 0.6 ;
      RECT 0.34 0 0.94 0.6 ;
  END
END nem_ohmux_invd0_4i_8b

END LIBRARY
