VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MANUFACTURINGGRID 0.005 ;

MACRO nem_ohmux_invd2_10i_8b
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN nem_ohmux_invd2_10i_8b 0 0 ;
  SIZE 20.18 BY 8.16 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN I0_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.34 6.65 2.51 6.82 ;
    END
  END I0_0
  PIN I0_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.95 6.49 2.12 6.66 ;
    END
  END I0_7
  PIN I0_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.045 6.34 3.215 6.51 ;
    END
  END I0_1
  PIN I0_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.185 6.01 3.355 6.18 ;
    END
  END I0_2
  PIN I0_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.95 5.315 3.12 5.485 ;
    END
  END I0_3
  PIN I0_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.56 5.16 2.73 5.33 ;
    END
  END I0_4
  PIN I0_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.84 5.435 2.01 5.605 ;
    END
  END I0_5
  PIN I0_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.695 5.775 1.865 5.945 ;
    END
  END I0_6
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.28 5.875 2.45 6.045 ;
    END
  END S0
  PIN ZN_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.48 7.565 9.625 7.645 ;
        RECT 9.555 6.815 9.625 7.645 ;
        RECT 9.48 6.815 9.625 6.895 ;
    END
  END ZN_7
  PIN ZN_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.32 7.565 10.465 7.645 ;
        RECT 10.395 6.815 10.465 7.645 ;
        RECT 10.32 6.815 10.465 6.895 ;
    END
  END ZN_2
  PIN ZN_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.9 7.565 10.045 7.645 ;
        RECT 9.975 6.815 10.045 7.645 ;
        RECT 9.9 6.815 10.045 6.895 ;
    END
  END ZN_0
  PIN ZN_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.74 7.565 10.885 7.645 ;
        RECT 10.815 6.815 10.885 7.645 ;
        RECT 10.74 6.815 10.885 6.895 ;
    END
  END ZN_1
  PIN ZN_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.74 5.045 10.885 5.125 ;
        RECT 10.815 4.295 10.885 5.125 ;
        RECT 10.74 4.295 10.885 4.375 ;
    END
  END ZN_3
  PIN ZN_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.275 3.785 9.42 3.865 ;
        RECT 9.275 3.035 9.42 3.115 ;
        RECT 9.275 3.035 9.345 3.865 ;
    END
  END ZN_4
  PIN ZN_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.32 5.045 10.465 5.125 ;
        RECT 10.395 4.295 10.465 5.125 ;
        RECT 10.32 4.295 10.465 4.375 ;
    END
  END ZN_6
  PIN ZN_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.48 5.045 9.625 5.125 ;
        RECT 9.555 4.295 9.625 5.125 ;
        RECT 9.48 4.295 9.625 4.375 ;
    END
  END ZN_5
  PIN I1_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.045 2.56 3.215 2.73 ;
    END
  END I1_3
  PIN I1_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.34 2.87 2.51 3.04 ;
    END
  END I1_4
  PIN I1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.95 1.535 3.12 1.705 ;
    END
  END I1_1
  PIN I1_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.84 1.655 2.01 1.825 ;
    END
  END I1_7
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.365 2.095 2.535 2.265 ;
    END
  END S1
  PIN I1_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.695 1.995 1.865 2.165 ;
    END
  END I1_6
  PIN I1_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.185 2.23 3.355 2.4 ;
    END
  END I1_2
  PIN I1_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.95 2.71 2.12 2.88 ;
    END
  END I1_5
  PIN I1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.56 1.38 2.73 1.55 ;
    END
  END I1_0
  PIN VSNEM
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M8 ;
        RECT 0 0 1.28 8.16 ;
    END
    PORT
      LAYER M8 ;
        RECT 3.78 0 5.06 8.16 ;
    END
    PORT
      LAYER M8 ;
        RECT 7.56 0 8.84 8.16 ;
    END
    PORT
      LAYER M8 ;
        RECT 11.34 0 12.62 8.16 ;
    END
    PORT
      LAYER M8 ;
        RECT 15.12 0 16.4 8.16 ;
    END
    PORT
      LAYER M8 ;
        RECT 18.9 0 20.18 8.16 ;
    END
  END VSNEM
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 9.24 2.705 9.66 2.935 ;
        RECT 9.5 2.705 9.58 3.145 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.24 7.745 10.92 7.975 ;
        RECT 10.58 7.535 10.66 7.975 ;
        RECT 10.16 7.535 10.24 7.975 ;
        RECT 9.74 7.535 9.82 7.975 ;
        RECT 9.32 7.535 9.4 7.975 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.24 5.225 10.92 5.455 ;
        RECT 10.58 5.015 10.66 5.455 ;
        RECT 10.16 5.015 10.24 5.455 ;
        RECT 9.32 5.015 9.4 5.455 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 9.24 6.485 10.92 6.715 ;
        RECT 10.58 6.485 10.66 6.925 ;
        RECT 10.16 6.485 10.24 6.925 ;
        RECT 9.74 6.485 9.82 6.925 ;
        RECT 9.32 6.485 9.4 6.925 ;
    END
    PORT
      LAYER M1 ;
        RECT 9.24 3.965 10.92 4.195 ;
        RECT 10.58 3.965 10.66 4.405 ;
        RECT 10.16 3.965 10.24 4.405 ;
        RECT 9.5 3.755 9.58 4.195 ;
        RECT 9.32 3.965 9.4 4.405 ;
    END
  END VSS
  PIN I2_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.73 6.49 5.9 6.66 ;
    END
  END I2_7
  PIN I2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.12 6.65 6.29 6.82 ;
    END
  END I2_0
  PIN I3_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.12 2.87 6.29 3.04 ;
    END
  END I3_4
  PIN I3_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.475 1.995 5.645 2.165 ;
    END
  END I3_6
  PIN I3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.73 1.535 6.9 1.705 ;
    END
  END I3_1
  PIN I2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.825 6.34 6.995 6.51 ;
    END
  END I2_1
  PIN I2_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.965 6.01 7.135 6.18 ;
    END
  END I2_2
  PIN I2_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.73 5.315 6.9 5.485 ;
    END
  END I2_3
  PIN I2_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.34 5.16 6.51 5.33 ;
    END
  END I2_4
  PIN I3_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.825 2.56 6.995 2.73 ;
    END
  END I3_3
  PIN I2_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.62 5.435 5.79 5.605 ;
    END
  END I2_5
  PIN I3_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.965 2.23 7.135 2.4 ;
    END
  END I3_2
  PIN I3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.34 1.38 6.51 1.55 ;
    END
  END I3_0
  PIN I3_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.73 2.71 5.9 2.88 ;
    END
  END I3_5
  PIN S3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.145 2.095 6.315 2.265 ;
    END
  END S3
  PIN I2_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.475 5.775 5.645 5.945 ;
    END
  END I2_6
  PIN I3_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.62 1.655 5.79 1.825 ;
    END
  END I3_7
  PIN S2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.06 5.875 6.23 6.045 ;
    END
  END S2
  PIN I4_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.245 5.775 9.415 5.945 ;
    END
  END I4_6
  PIN I4_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.4 5.435 9.57 5.605 ;
    END
  END I4_5
  PIN I4_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.455 6.49 9.625 6.66 ;
    END
  END I4_7
  PIN S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.025 5.875 10.195 6.045 ;
    END
  END S4
  PIN I4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.875 6.65 10.045 6.82 ;
    END
  END I4_0
  PIN I4_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.135 5.165 10.305 5.335 ;
    END
  END I4_4
  PIN I4_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.51 5.315 10.68 5.485 ;
    END
  END I4_3
  PIN I4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.605 6.34 10.775 6.51 ;
    END
  END I4_1
  PIN I4_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.755 6.01 10.925 6.18 ;
    END
  END I4_2
  PIN I5_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.24 1.995 9.41 2.165 ;
    END
  END I5_6
  PIN I5_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.39 1.655 9.56 1.825 ;
    END
  END I5_7
  PIN I5_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.505 2.67 9.675 2.84 ;
    END
  END I5_5
  PIN I5_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.875 2.87 10.045 3.04 ;
    END
  END I5_4
  PIN I5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.13 1.38 10.3 1.55 ;
    END
  END I5_0
  PIN I5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.485 1.535 10.655 1.705 ;
    END
  END I5_1
  PIN I5_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.605 2.56 10.775 2.73 ;
    END
  END I5_3
  PIN I5_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 10.755 2.23 10.925 2.4 ;
    END
  END I5_2
  PIN S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 9.925 2.095 10.095 2.265 ;
    END
  END S5
  PIN I6_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.035 5.775 13.205 5.945 ;
    END
  END I6_6
  PIN I6_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.18 5.435 13.35 5.605 ;
    END
  END I6_5
  PIN I6_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.29 6.49 13.46 6.66 ;
    END
  END I6_7
  PIN S6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.62 5.875 13.79 6.045 ;
    END
  END S6
  PIN I6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.68 6.65 13.85 6.82 ;
    END
  END I6_0
  PIN I6_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.9 5.16 14.07 5.33 ;
    END
  END I6_4
  PIN I6_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.29 5.315 14.46 5.485 ;
    END
  END I6_3
  PIN I6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.385 6.34 14.555 6.51 ;
    END
  END I6_1
  PIN I6_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.525 6.01 14.695 6.18 ;
    END
  END I6_2
  PIN I7_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.035 1.995 13.205 2.165 ;
    END
  END I7_6
  PIN I7_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.18 1.655 13.35 1.825 ;
    END
  END I7_7
  PIN I7_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.29 2.71 13.46 2.88 ;
    END
  END I7_5
  PIN I7_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.68 2.87 13.85 3.04 ;
    END
  END I7_4
  PIN S7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.705 2.095 13.875 2.265 ;
    END
  END S7
  PIN I7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 13.9 1.38 14.07 1.55 ;
    END
  END I7_0
  PIN I7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.29 1.535 14.46 1.705 ;
    END
  END I7_1
  PIN I7_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.385 2.56 14.555 2.73 ;
    END
  END I7_3
  PIN I7_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 14.525 2.23 14.695 2.4 ;
    END
  END I7_2
  PIN I9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.07 1.535 18.24 1.705 ;
    END
  END I9_1
  PIN I9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.68 1.38 17.85 1.55 ;
    END
  END I9_0
  PIN S9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.485 2.095 17.655 2.265 ;
    END
  END S9
  PIN I9_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.46 2.87 17.63 3.04 ;
    END
  END I9_4
  PIN I9_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.07 2.71 17.24 2.88 ;
    END
  END I9_5
  PIN I9_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 16.96 1.655 17.13 1.825 ;
    END
  END I9_7
  PIN I9_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 16.815 1.995 16.985 2.165 ;
    END
  END I9_6
  PIN I8_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.305 6.01 18.475 6.18 ;
    END
  END I8_2
  PIN I8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.165 6.34 18.335 6.51 ;
    END
  END I8_1
  PIN I9_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.305 2.23 18.475 2.4 ;
    END
  END I9_2
  PIN I9_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.165 2.56 18.335 2.73 ;
    END
  END I9_3
  PIN I8_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 18.07 5.315 18.24 5.485 ;
    END
  END I8_3
  PIN I8_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.68 5.16 17.85 5.33 ;
    END
  END I8_4
  PIN I8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.46 6.65 17.63 6.82 ;
    END
  END I8_0
  PIN S8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.4 5.875 17.57 6.045 ;
    END
  END S8
  PIN I8_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 17.07 6.49 17.24 6.66 ;
    END
  END I8_7
  PIN I8_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 16.96 5.435 17.13 5.605 ;
    END
  END I8_5
  PIN I8_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 16.815 5.775 16.985 5.945 ;
    END
  END I8_6
  OBS
    LAYER OVERLAP ;
      RECT 0 0 20.18 8.16 ;
    LAYER M1 ;
      RECT 10.535 4.575 10.605 4.845 ;
      RECT 10.535 4.625 10.74 4.695 ;
      RECT 10.535 7.095 10.605 7.365 ;
      RECT 10.535 7.145 10.74 7.215 ;
      RECT 10.115 4.575 10.185 4.845 ;
      RECT 10.115 4.625 10.32 4.695 ;
      RECT 10.115 7.095 10.185 7.365 ;
      RECT 10.115 7.145 10.32 7.215 ;
      RECT 9.695 7.095 9.765 7.365 ;
      RECT 9.695 7.145 9.9 7.215 ;
      RECT 9.555 3.315 9.625 3.585 ;
      RECT 9.42 3.465 9.625 3.535 ;
      RECT 9.275 4.575 9.345 4.845 ;
      RECT 9.275 4.625 9.48 4.695 ;
      RECT 9.275 7.095 9.345 7.365 ;
      RECT 9.275 7.145 9.48 7.215 ;
    LAYER M2 ;
      RECT 10.535 4.455 10.605 4.845 ;
      RECT 10.535 6.975 10.605 7.365 ;
      RECT 10.115 4.455 10.185 4.845 ;
      RECT 10.115 6.975 10.185 7.365 ;
      RECT 9.695 6.975 9.765 7.365 ;
      RECT 9.555 3.195 9.625 3.585 ;
      RECT 9.275 4.455 9.345 4.845 ;
      RECT 9.275 6.975 9.345 7.365 ;
    LAYER M3 ;
      RECT 10.535 4.455 10.605 4.845 ;
      RECT 10.535 6.975 10.605 7.365 ;
      RECT 10.115 4.455 10.185 4.845 ;
      RECT 10.115 6.975 10.185 7.365 ;
      RECT 9.695 6.975 9.765 7.365 ;
      RECT 9.555 3.195 9.625 3.585 ;
      RECT 9.275 4.455 9.345 4.845 ;
      RECT 9.275 6.975 9.345 7.365 ;
    LAYER M4 ;
      RECT 10.535 4.455 10.605 4.845 ;
      RECT 10.535 6.975 10.605 7.365 ;
      RECT 10.115 4.455 10.185 4.845 ;
      RECT 10.115 6.975 10.185 7.365 ;
      RECT 9.695 6.975 9.765 7.365 ;
      RECT 9.555 3.195 9.625 3.585 ;
      RECT 9.275 4.455 9.345 4.845 ;
      RECT 9.275 6.975 9.345 7.365 ;
    LAYER M5 ;
      RECT 10.535 4.455 10.605 4.845 ;
      RECT 10.535 6.975 10.605 7.365 ;
      RECT 10.115 4.455 10.185 4.845 ;
      RECT 10.115 6.975 10.185 7.365 ;
      RECT 9.695 6.975 9.765 7.365 ;
      RECT 9.555 3.195 9.625 3.585 ;
      RECT 9.275 4.455 9.345 4.845 ;
      RECT 9.275 6.975 9.345 7.365 ;
    LAYER M6 ;
      RECT 10.535 4.575 10.605 5.255 ;
      RECT 10.535 6.65 10.605 7.365 ;
      RECT 10.115 4.575 10.185 5.105 ;
      RECT 10.115 6.65 10.185 7.365 ;
      RECT 9.695 6.65 9.765 7.365 ;
      RECT 9.555 2.91 9.625 3.585 ;
      RECT 9.275 4.575 9.345 5.365 ;
      RECT 9.275 6.65 9.345 7.365 ;
    LAYER M7 ;
      RECT 10.505 4.995 10.64 5.235 ;
      RECT 10.53 6.58 10.61 6.92 ;
      RECT 10.02 4.99 10.285 5.095 ;
      RECT 10.115 6.53 10.185 6.92 ;
      RECT 9.695 6.53 9.765 6.92 ;
      RECT 9.535 2.91 9.645 3.17 ;
      RECT 9.27 5.025 9.35 5.365 ;
      RECT 9.275 6.53 9.345 6.92 ;
    LAYER M8 ;
      RECT 18.545 7.115 18.675 7.245 ;
      RECT 18.575 2.15 18.645 7.245 ;
      RECT 18.545 5.93 18.675 6.06 ;
      RECT 18.545 3.335 18.675 3.465 ;
      RECT 18.545 2.15 18.675 2.28 ;
      RECT 18.335 7.515 18.465 7.645 ;
      RECT 18.365 6.665 18.435 7.645 ;
      RECT 18.335 6.665 18.465 6.795 ;
      RECT 17.925 6.695 18.465 6.765 ;
      RECT 17.925 4.28 17.995 6.765 ;
      RECT 17.925 4.28 18.175 4.35 ;
      RECT 18.105 2.905 18.175 4.35 ;
      RECT 17.99 2.905 18.175 2.975 ;
      RECT 17.99 1.81 18.06 2.975 ;
      RECT 17.99 1.81 18.46 1.88 ;
      RECT 18.39 0.505 18.46 1.88 ;
      RECT 18.36 1.37 18.49 1.5 ;
      RECT 18.36 0.505 18.49 0.635 ;
      RECT 18.36 5.15 18.49 5.28 ;
      RECT 18.39 3.735 18.46 5.28 ;
      RECT 18.36 4.285 18.49 4.415 ;
      RECT 18.33 3.735 18.46 3.865 ;
      RECT 18.365 2.885 18.435 3.865 ;
      RECT 18.335 2.885 18.465 3.015 ;
      RECT 17.77 1.735 17.84 4.21 ;
      RECT 17.495 1.735 17.84 1.805 ;
      RECT 17.495 1.105 17.565 1.805 ;
      RECT 17.465 1.105 17.595 1.235 ;
      RECT 17.68 6.915 17.81 7.045 ;
      RECT 17.71 5.73 17.78 7.045 ;
      RECT 17.41 5.73 17.78 5.8 ;
      RECT 17.41 3.94 17.48 5.8 ;
      RECT 17.56 4.885 17.69 5.015 ;
      RECT 17.59 3.135 17.66 5.015 ;
      RECT 17.56 3.135 17.69 3.265 ;
      RECT 16.86 7.315 16.99 7.445 ;
      RECT 16.89 6.04 16.96 7.445 ;
      RECT 16.82 6.65 16.96 6.78 ;
      RECT 16.89 6.04 17.295 6.11 ;
      RECT 17.225 4.88 17.295 6.11 ;
      RECT 17.1 4.88 17.295 4.95 ;
      RECT 17.1 3.06 17.17 4.95 ;
      RECT 17.1 3.06 17.38 3.13 ;
      RECT 17.31 1.44 17.38 3.13 ;
      RECT 16.83 1.44 17.38 1.51 ;
      RECT 16.83 1.38 16.96 1.51 ;
      RECT 16.86 0.705 16.93 1.51 ;
      RECT 16.83 0.705 16.96 0.835 ;
      RECT 16.83 5.16 16.96 5.29 ;
      RECT 16.86 3.535 16.93 5.29 ;
      RECT 16.83 4.485 16.96 4.615 ;
      RECT 16.86 3.535 16.99 3.665 ;
      RECT 16.89 2.87 16.96 3.665 ;
      RECT 16.82 2.87 16.96 3 ;
      RECT 16.615 5.89 16.745 6.02 ;
      RECT 16.645 0.905 16.715 6.02 ;
      RECT 16.615 4.685 16.745 4.815 ;
      RECT 16.615 2.11 16.745 2.24 ;
      RECT 16.615 0.905 16.745 1.035 ;
      RECT 14.765 7.115 14.895 7.245 ;
      RECT 14.795 2.15 14.865 7.245 ;
      RECT 14.765 5.93 14.895 6.06 ;
      RECT 14.765 3.335 14.895 3.465 ;
      RECT 14.765 2.15 14.895 2.28 ;
      RECT 14.555 7.515 14.685 7.645 ;
      RECT 14.585 6.665 14.655 7.645 ;
      RECT 14.555 6.665 14.685 6.795 ;
      RECT 14.145 6.695 14.685 6.765 ;
      RECT 14.145 4.28 14.215 6.765 ;
      RECT 14.145 4.28 14.395 4.35 ;
      RECT 14.325 2.905 14.395 4.35 ;
      RECT 14.21 2.905 14.395 2.975 ;
      RECT 14.21 1.81 14.28 2.975 ;
      RECT 14.21 1.81 14.68 1.88 ;
      RECT 14.61 0.505 14.68 1.88 ;
      RECT 14.58 1.37 14.71 1.5 ;
      RECT 14.58 0.505 14.71 0.635 ;
      RECT 14.58 5.15 14.71 5.28 ;
      RECT 14.61 3.735 14.68 5.28 ;
      RECT 14.58 4.285 14.71 4.415 ;
      RECT 14.55 3.735 14.68 3.865 ;
      RECT 14.585 2.885 14.655 3.865 ;
      RECT 14.555 2.885 14.685 3.015 ;
      RECT 13.99 1.735 14.06 4.21 ;
      RECT 13.715 1.735 14.06 1.805 ;
      RECT 13.715 1.105 13.785 1.805 ;
      RECT 13.685 1.105 13.815 1.235 ;
      RECT 13.9 6.915 14.03 7.045 ;
      RECT 13.93 5.73 14 7.045 ;
      RECT 13.63 5.73 14 5.8 ;
      RECT 13.63 3.94 13.7 5.8 ;
      RECT 13.78 4.885 13.91 5.015 ;
      RECT 13.81 3.135 13.88 5.015 ;
      RECT 13.78 3.135 13.91 3.265 ;
      RECT 13.08 7.315 13.21 7.445 ;
      RECT 13.11 6.04 13.18 7.445 ;
      RECT 13.04 6.65 13.18 6.78 ;
      RECT 13.11 6.04 13.515 6.11 ;
      RECT 13.445 4.88 13.515 6.11 ;
      RECT 13.32 4.88 13.515 4.95 ;
      RECT 13.32 3.06 13.39 4.95 ;
      RECT 13.32 3.06 13.6 3.13 ;
      RECT 13.53 1.44 13.6 3.13 ;
      RECT 13.05 1.44 13.6 1.51 ;
      RECT 13.05 1.38 13.18 1.51 ;
      RECT 13.08 0.705 13.15 1.51 ;
      RECT 13.05 0.705 13.18 0.835 ;
      RECT 13.05 5.16 13.18 5.29 ;
      RECT 13.08 3.535 13.15 5.29 ;
      RECT 13.05 4.485 13.18 4.615 ;
      RECT 13.08 3.535 13.21 3.665 ;
      RECT 13.11 2.87 13.18 3.665 ;
      RECT 13.04 2.87 13.18 3 ;
      RECT 12.835 5.89 12.965 6.02 ;
      RECT 12.865 0.905 12.935 6.02 ;
      RECT 12.835 4.685 12.965 4.815 ;
      RECT 12.835 2.11 12.965 2.24 ;
      RECT 12.835 0.905 12.965 1.035 ;
      RECT 10.985 7.115 11.115 7.245 ;
      RECT 11.015 2.15 11.085 7.245 ;
      RECT 10.985 5.93 11.115 6.06 ;
      RECT 10.985 3.335 11.115 3.465 ;
      RECT 10.985 2.15 11.115 2.28 ;
      RECT 10.365 3.535 10.435 6.785 ;
      RECT 10.365 3.535 10.62 3.605 ;
      RECT 10.55 2.905 10.62 3.605 ;
      RECT 10.435 2.905 10.62 2.975 ;
      RECT 10.435 1.81 10.505 2.975 ;
      RECT 10.435 1.81 10.9 1.88 ;
      RECT 10.83 0.505 10.9 1.88 ;
      RECT 10.8 1.37 10.93 1.5 ;
      RECT 10.8 0.505 10.93 0.635 ;
      RECT 10.8 5.15 10.93 5.28 ;
      RECT 10.83 3.735 10.9 5.28 ;
      RECT 10.8 4.285 10.93 4.415 ;
      RECT 10.77 3.735 10.9 3.865 ;
      RECT 10.805 2.885 10.875 3.865 ;
      RECT 10.775 2.885 10.905 3.015 ;
      RECT 10.775 7.515 10.905 7.645 ;
      RECT 10.805 6.665 10.875 7.645 ;
      RECT 10.775 6.665 10.905 6.795 ;
      RECT 10.535 4.285 10.605 5.245 ;
      RECT 10.505 4.285 10.635 4.415 ;
      RECT 10.505 7.515 10.635 7.645 ;
      RECT 10.535 6.65 10.605 7.645 ;
      RECT 9.665 6.915 9.795 7.045 ;
      RECT 9.695 6.275 9.765 7.045 ;
      RECT 9.695 6.275 9.915 6.345 ;
      RECT 9.845 5.125 9.915 6.345 ;
      RECT 9.915 3.4 9.985 5.195 ;
      RECT 9.915 3.4 10.29 3.47 ;
      RECT 10.22 1.735 10.29 3.47 ;
      RECT 9.94 1.735 10.29 1.805 ;
      RECT 9.94 1.105 10.01 1.805 ;
      RECT 9.91 1.105 10.04 1.235 ;
      RECT 10.115 4.685 10.185 5.095 ;
      RECT 10.085 4.685 10.215 4.815 ;
      RECT 10.085 7.115 10.215 7.245 ;
      RECT 10.115 6.53 10.185 7.245 ;
      RECT 9.245 7.315 9.375 7.445 ;
      RECT 9.275 6.04 9.345 7.445 ;
      RECT 9.26 6.65 9.39 6.78 ;
      RECT 9.275 6.04 9.735 6.11 ;
      RECT 9.665 4.88 9.735 6.11 ;
      RECT 9.665 4.88 9.82 4.95 ;
      RECT 9.75 1.44 9.82 4.95 ;
      RECT 9.27 1.44 9.82 1.51 ;
      RECT 9.27 1.38 9.4 1.51 ;
      RECT 9.3 0.705 9.37 1.51 ;
      RECT 9.27 0.705 9.4 0.835 ;
      RECT 9.455 4.885 9.585 5.015 ;
      RECT 9.455 3.67 9.525 5.015 ;
      RECT 9.455 3.67 9.625 3.74 ;
      RECT 9.555 2.91 9.625 3.74 ;
      RECT 9.525 3.135 9.655 3.265 ;
      RECT 9.245 5.16 9.375 5.29 ;
      RECT 9.275 2.87 9.345 5.29 ;
      RECT 9.24 4.485 9.37 4.615 ;
      RECT 9.24 3.535 9.37 3.665 ;
      RECT 9.275 2.87 9.405 3 ;
      RECT 9.055 5.89 9.185 6.02 ;
      RECT 9.085 0.905 9.155 6.02 ;
      RECT 9.055 4.685 9.185 4.815 ;
      RECT 9.055 2.11 9.185 2.24 ;
      RECT 9.055 0.905 9.185 1.035 ;
      RECT 7.205 7.115 7.335 7.245 ;
      RECT 7.235 2.15 7.305 7.245 ;
      RECT 7.205 5.93 7.335 6.06 ;
      RECT 7.205 3.335 7.335 3.465 ;
      RECT 7.205 2.15 7.335 2.28 ;
      RECT 6.995 7.515 7.125 7.645 ;
      RECT 7.025 6.665 7.095 7.645 ;
      RECT 6.995 6.665 7.125 6.795 ;
      RECT 6.585 6.695 7.125 6.765 ;
      RECT 6.585 4.28 6.655 6.765 ;
      RECT 6.585 4.28 6.835 4.35 ;
      RECT 6.765 2.905 6.835 4.35 ;
      RECT 6.65 2.905 6.835 2.975 ;
      RECT 6.65 1.81 6.72 2.975 ;
      RECT 6.65 1.81 7.12 1.88 ;
      RECT 7.05 0.505 7.12 1.88 ;
      RECT 7.02 1.37 7.15 1.5 ;
      RECT 7.02 0.505 7.15 0.635 ;
      RECT 7.02 5.15 7.15 5.28 ;
      RECT 7.05 3.735 7.12 5.28 ;
      RECT 7.02 4.285 7.15 4.415 ;
      RECT 6.99 3.735 7.12 3.865 ;
      RECT 7.025 2.885 7.095 3.865 ;
      RECT 6.995 2.885 7.125 3.015 ;
      RECT 6.43 1.735 6.5 4.21 ;
      RECT 6.155 1.735 6.5 1.805 ;
      RECT 6.155 1.105 6.225 1.805 ;
      RECT 6.125 1.105 6.255 1.235 ;
      RECT 6.34 6.915 6.47 7.045 ;
      RECT 6.37 5.73 6.44 7.045 ;
      RECT 6.07 5.73 6.44 5.8 ;
      RECT 6.07 3.94 6.14 5.8 ;
      RECT 6.22 4.885 6.35 5.015 ;
      RECT 6.25 3.135 6.32 5.015 ;
      RECT 6.22 3.135 6.35 3.265 ;
      RECT 5.52 7.315 5.65 7.445 ;
      RECT 5.55 6.04 5.62 7.445 ;
      RECT 5.48 6.65 5.62 6.78 ;
      RECT 5.55 6.04 5.955 6.11 ;
      RECT 5.885 4.88 5.955 6.11 ;
      RECT 5.76 4.88 5.955 4.95 ;
      RECT 5.76 3.06 5.83 4.95 ;
      RECT 5.76 3.06 6.04 3.13 ;
      RECT 5.97 1.44 6.04 3.13 ;
      RECT 5.49 1.44 6.04 1.51 ;
      RECT 5.49 1.38 5.62 1.51 ;
      RECT 5.52 0.705 5.59 1.51 ;
      RECT 5.49 0.705 5.62 0.835 ;
      RECT 5.49 5.16 5.62 5.29 ;
      RECT 5.52 3.535 5.59 5.29 ;
      RECT 5.49 4.485 5.62 4.615 ;
      RECT 5.52 3.535 5.65 3.665 ;
      RECT 5.55 2.87 5.62 3.665 ;
      RECT 5.48 2.87 5.62 3 ;
      RECT 5.275 5.89 5.405 6.02 ;
      RECT 5.305 0.905 5.375 6.02 ;
      RECT 5.275 4.685 5.405 4.815 ;
      RECT 5.275 2.11 5.405 2.24 ;
      RECT 5.275 0.905 5.405 1.035 ;
      RECT 3.425 7.115 3.555 7.245 ;
      RECT 3.455 2.15 3.525 7.245 ;
      RECT 3.425 5.93 3.555 6.06 ;
      RECT 3.425 3.335 3.555 3.465 ;
      RECT 3.425 2.15 3.555 2.28 ;
      RECT 3.215 7.515 3.345 7.645 ;
      RECT 3.245 6.665 3.315 7.645 ;
      RECT 3.215 6.665 3.345 6.795 ;
      RECT 2.805 6.695 3.345 6.765 ;
      RECT 2.805 4.28 2.875 6.765 ;
      RECT 2.805 4.28 3.055 4.35 ;
      RECT 2.985 2.905 3.055 4.35 ;
      RECT 2.87 2.905 3.055 2.975 ;
      RECT 2.87 1.81 2.94 2.975 ;
      RECT 2.87 1.81 3.34 1.88 ;
      RECT 3.27 0.505 3.34 1.88 ;
      RECT 3.24 1.37 3.37 1.5 ;
      RECT 3.24 0.505 3.37 0.635 ;
      RECT 3.24 5.15 3.37 5.28 ;
      RECT 3.27 3.735 3.34 5.28 ;
      RECT 3.24 4.285 3.37 4.415 ;
      RECT 3.21 3.735 3.34 3.865 ;
      RECT 3.245 2.885 3.315 3.865 ;
      RECT 3.215 2.885 3.345 3.015 ;
      RECT 2.65 1.735 2.72 4.21 ;
      RECT 2.375 1.735 2.72 1.805 ;
      RECT 2.375 1.105 2.445 1.805 ;
      RECT 2.345 1.105 2.475 1.235 ;
      RECT 2.56 6.915 2.69 7.045 ;
      RECT 2.59 5.73 2.66 7.045 ;
      RECT 2.29 5.73 2.66 5.8 ;
      RECT 2.29 3.94 2.36 5.8 ;
      RECT 2.44 4.885 2.57 5.015 ;
      RECT 2.47 3.135 2.54 5.015 ;
      RECT 2.44 3.135 2.57 3.265 ;
      RECT 1.74 7.315 1.87 7.445 ;
      RECT 1.77 6.04 1.84 7.445 ;
      RECT 1.7 6.65 1.84 6.78 ;
      RECT 1.77 6.04 2.175 6.11 ;
      RECT 2.105 4.88 2.175 6.11 ;
      RECT 1.98 4.88 2.175 4.95 ;
      RECT 1.98 3.06 2.05 4.95 ;
      RECT 1.98 3.06 2.26 3.13 ;
      RECT 2.19 1.44 2.26 3.13 ;
      RECT 1.71 1.44 2.26 1.51 ;
      RECT 1.71 1.38 1.84 1.51 ;
      RECT 1.74 0.705 1.81 1.51 ;
      RECT 1.71 0.705 1.84 0.835 ;
      RECT 1.71 5.16 1.84 5.29 ;
      RECT 1.74 3.535 1.81 5.29 ;
      RECT 1.71 4.485 1.84 4.615 ;
      RECT 1.74 3.535 1.87 3.665 ;
      RECT 1.77 2.87 1.84 3.665 ;
      RECT 1.7 2.87 1.84 3 ;
      RECT 1.495 5.89 1.625 6.02 ;
      RECT 1.525 0.905 1.595 6.02 ;
      RECT 1.495 4.685 1.625 4.815 ;
      RECT 1.495 2.11 1.625 2.24 ;
      RECT 1.495 0.905 1.625 1.035 ;
      RECT 18.305 2.22 18.475 2.39 ;
      RECT 18.305 6.005 18.475 6.175 ;
      RECT 18.165 2.58 18.335 2.75 ;
      RECT 18.165 6.345 18.335 6.515 ;
      RECT 18.07 1.535 18.24 1.705 ;
      RECT 18.07 5.315 18.24 5.485 ;
      RECT 17.68 1.385 17.85 1.555 ;
      RECT 17.68 5.165 17.85 5.335 ;
      RECT 17.485 2.09 17.655 2.26 ;
      RECT 17.46 2.87 17.63 3.04 ;
      RECT 17.46 6.65 17.63 6.82 ;
      RECT 17.4 5.87 17.57 6.04 ;
      RECT 17.07 2.71 17.24 2.88 ;
      RECT 17.07 6.49 17.24 6.66 ;
      RECT 16.96 1.635 17.13 1.805 ;
      RECT 16.96 5.415 17.13 5.585 ;
      RECT 16.815 1.99 16.985 2.16 ;
      RECT 16.815 5.77 16.985 5.94 ;
      RECT 14.525 2.22 14.695 2.39 ;
      RECT 14.525 6.005 14.695 6.175 ;
      RECT 14.385 2.58 14.555 2.75 ;
      RECT 14.385 6.345 14.555 6.515 ;
      RECT 14.29 1.535 14.46 1.705 ;
      RECT 14.29 5.315 14.46 5.485 ;
      RECT 13.9 1.385 14.07 1.555 ;
      RECT 13.9 5.165 14.07 5.335 ;
      RECT 13.705 2.09 13.875 2.26 ;
      RECT 13.68 2.87 13.85 3.04 ;
      RECT 13.68 6.65 13.85 6.82 ;
      RECT 13.62 5.87 13.79 6.04 ;
      RECT 13.29 2.71 13.46 2.88 ;
      RECT 13.29 6.49 13.46 6.66 ;
      RECT 13.18 1.635 13.35 1.805 ;
      RECT 13.18 5.415 13.35 5.585 ;
      RECT 13.035 1.99 13.205 2.16 ;
      RECT 13.035 5.77 13.205 5.94 ;
      RECT 10.745 2.225 10.915 2.395 ;
      RECT 10.745 6.005 10.915 6.175 ;
      RECT 10.605 2.565 10.775 2.735 ;
      RECT 10.605 6.345 10.775 6.515 ;
      RECT 10.51 1.535 10.68 1.705 ;
      RECT 10.51 5.315 10.68 5.485 ;
      RECT 10.12 1.385 10.29 1.555 ;
      RECT 10.12 5.165 10.29 5.335 ;
      RECT 10.025 5.87 10.195 6.04 ;
      RECT 9.925 2.09 10.095 2.26 ;
      RECT 9.9 2.87 10.07 3.04 ;
      RECT 9.875 6.65 10.045 6.82 ;
      RECT 9.51 2.67 9.68 2.84 ;
      RECT 9.465 6.49 9.625 6.675 ;
      RECT 9.4 1.635 9.57 1.805 ;
      RECT 9.39 5.415 9.56 5.585 ;
      RECT 9.255 1.99 9.425 2.16 ;
      RECT 9.255 5.77 9.425 5.94 ;
      RECT 6.965 2.22 7.135 2.39 ;
      RECT 6.965 6.005 7.135 6.175 ;
      RECT 6.825 2.58 6.995 2.75 ;
      RECT 6.825 6.345 6.995 6.515 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.73 5.315 6.9 5.485 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.34 5.165 6.51 5.335 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 6.12 2.87 6.29 3.04 ;
      RECT 6.12 6.65 6.29 6.82 ;
      RECT 6.06 5.87 6.23 6.04 ;
      RECT 5.73 2.71 5.9 2.88 ;
      RECT 5.73 6.49 5.9 6.66 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.62 5.415 5.79 5.585 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 5.475 5.77 5.645 5.94 ;
      RECT 3.185 2.22 3.355 2.39 ;
      RECT 3.185 6.005 3.355 6.175 ;
      RECT 3.045 2.58 3.215 2.75 ;
      RECT 3.045 6.345 3.215 6.515 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.95 5.315 3.12 5.485 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.56 5.165 2.73 5.335 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 2.34 2.87 2.51 3.04 ;
      RECT 2.34 6.65 2.51 6.82 ;
      RECT 2.28 5.87 2.45 6.04 ;
      RECT 1.95 2.71 2.12 2.88 ;
      RECT 1.95 6.49 2.12 6.66 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.84 5.415 2.01 5.585 ;
      RECT 1.695 1.99 1.865 2.16 ;
      RECT 1.695 5.77 1.865 5.94 ;
    LAYER M9 ;
      RECT 17.75 3.96 17.86 4.19 ;
      RECT 17.39 3.96 17.5 4.19 ;
      RECT 17.39 4.04 17.86 4.11 ;
      RECT 13.97 3.96 14.08 4.19 ;
      RECT 13.61 3.96 13.72 4.19 ;
      RECT 13.61 4.04 14.08 4.11 ;
      RECT 10.755 6.645 10.925 6.815 ;
      RECT 10.345 6.695 10.925 6.765 ;
      RECT 10.345 6.535 10.455 6.765 ;
      RECT 6.41 3.96 6.52 4.19 ;
      RECT 6.05 3.96 6.16 4.19 ;
      RECT 6.05 4.04 6.52 4.11 ;
      RECT 2.63 3.96 2.74 4.19 ;
      RECT 2.27 3.96 2.38 4.19 ;
      RECT 2.27 4.04 2.74 4.11 ;
      RECT 19.39 0.165 19.69 0.435 ;
      RECT 19.39 3.945 19.69 4.215 ;
      RECT 19.39 7.725 19.69 7.995 ;
      RECT 18.545 2.15 18.78 2.28 ;
      RECT 18.545 5.93 18.78 6.06 ;
      RECT 1.495 0.505 18.675 0.635 ;
      RECT 1.495 0.705 18.675 0.835 ;
      RECT 1.495 0.905 18.675 1.035 ;
      RECT 1.495 1.105 18.675 1.235 ;
      RECT 1.495 3.135 18.675 3.265 ;
      RECT 1.495 3.335 18.675 3.465 ;
      RECT 1.495 3.535 18.675 3.665 ;
      RECT 1.495 3.735 18.675 3.865 ;
      RECT 1.495 4.285 18.675 4.415 ;
      RECT 1.495 4.485 18.675 4.615 ;
      RECT 1.495 4.685 18.675 4.815 ;
      RECT 1.495 4.885 18.675 5.015 ;
      RECT 1.495 6.915 18.675 7.045 ;
      RECT 1.495 7.115 18.675 7.245 ;
      RECT 1.495 7.315 18.675 7.445 ;
      RECT 1.495 7.515 18.675 7.645 ;
      RECT 18.34 1.35 18.51 1.52 ;
      RECT 18.34 5.13 18.51 5.3 ;
      RECT 18.315 2.865 18.485 3.035 ;
      RECT 18.315 6.645 18.485 6.815 ;
      RECT 18.305 2.22 18.475 2.39 ;
      RECT 18.305 6.005 18.475 6.175 ;
      RECT 18.165 2.58 18.335 2.75 ;
      RECT 18.165 6.345 18.335 6.515 ;
      RECT 18.07 1.535 18.24 1.705 ;
      RECT 18.07 5.315 18.24 5.485 ;
      RECT 17.68 1.385 17.85 1.555 ;
      RECT 17.68 5.165 17.85 5.335 ;
      RECT 17.485 2.09 17.655 2.26 ;
      RECT 17.46 2.87 17.63 3.04 ;
      RECT 17.46 6.65 17.63 6.82 ;
      RECT 17.4 5.87 17.57 6.04 ;
      RECT 17.07 2.71 17.24 2.88 ;
      RECT 17.07 6.49 17.24 6.66 ;
      RECT 16.96 1.635 17.13 1.805 ;
      RECT 16.96 5.415 17.13 5.585 ;
      RECT 16.815 1.99 16.985 2.16 ;
      RECT 16.815 5.77 16.985 5.94 ;
      RECT 16.81 1.36 16.98 1.53 ;
      RECT 16.81 5.14 16.98 5.31 ;
      RECT 16.8 2.85 16.97 3.02 ;
      RECT 16.8 6.63 16.97 6.8 ;
      RECT 16.53 2.11 16.745 2.24 ;
      RECT 16.53 5.89 16.745 6.02 ;
      RECT 15.61 0.165 15.91 0.435 ;
      RECT 15.61 3.945 15.91 4.215 ;
      RECT 15.61 7.725 15.91 7.995 ;
      RECT 14.765 2.15 15 2.28 ;
      RECT 14.765 5.93 15 6.06 ;
      RECT 14.56 1.35 14.73 1.52 ;
      RECT 14.56 5.13 14.73 5.3 ;
      RECT 14.535 2.865 14.705 3.035 ;
      RECT 14.535 6.645 14.705 6.815 ;
      RECT 14.525 2.22 14.695 2.39 ;
      RECT 14.525 6.005 14.695 6.175 ;
      RECT 14.385 2.58 14.555 2.75 ;
      RECT 14.385 6.345 14.555 6.515 ;
      RECT 14.29 1.535 14.46 1.705 ;
      RECT 14.29 5.315 14.46 5.485 ;
      RECT 13.9 1.385 14.07 1.555 ;
      RECT 13.9 5.165 14.07 5.335 ;
      RECT 13.705 2.09 13.875 2.26 ;
      RECT 13.68 2.87 13.85 3.04 ;
      RECT 13.68 6.65 13.85 6.82 ;
      RECT 13.62 5.87 13.79 6.04 ;
      RECT 13.29 2.71 13.46 2.88 ;
      RECT 13.29 6.49 13.46 6.66 ;
      RECT 13.18 1.635 13.35 1.805 ;
      RECT 13.18 5.415 13.35 5.585 ;
      RECT 13.035 1.99 13.205 2.16 ;
      RECT 13.035 5.77 13.205 5.94 ;
      RECT 13.03 1.36 13.2 1.53 ;
      RECT 13.03 5.14 13.2 5.31 ;
      RECT 13.02 2.85 13.19 3.02 ;
      RECT 13.02 6.63 13.19 6.8 ;
      RECT 12.75 2.11 12.965 2.24 ;
      RECT 12.75 5.89 12.965 6.02 ;
      RECT 11.83 0.165 12.13 0.435 ;
      RECT 11.83 3.945 12.13 4.215 ;
      RECT 11.83 7.725 12.13 7.995 ;
      RECT 10.985 2.15 11.22 2.28 ;
      RECT 10.985 5.93 11.22 6.06 ;
      RECT 10.78 1.35 10.95 1.52 ;
      RECT 10.78 5.13 10.95 5.3 ;
      RECT 10.755 2.865 10.925 3.035 ;
      RECT 10.745 2.225 10.915 2.395 ;
      RECT 10.745 6.005 10.915 6.175 ;
      RECT 10.605 2.565 10.775 2.735 ;
      RECT 10.605 6.345 10.775 6.515 ;
      RECT 10.51 1.535 10.68 1.705 ;
      RECT 10.51 5.315 10.68 5.485 ;
      RECT 10.12 1.385 10.29 1.555 ;
      RECT 10.12 5.165 10.29 5.335 ;
      RECT 10.025 5.87 10.195 6.04 ;
      RECT 9.925 2.09 10.095 2.26 ;
      RECT 9.9 2.87 10.07 3.04 ;
      RECT 9.875 6.65 10.045 6.82 ;
      RECT 9.51 2.71 9.68 2.88 ;
      RECT 9.51 6.49 9.68 6.66 ;
      RECT 9.4 1.635 9.57 1.805 ;
      RECT 9.39 5.415 9.56 5.585 ;
      RECT 9.255 1.99 9.425 2.16 ;
      RECT 9.255 2.85 9.425 3.02 ;
      RECT 9.255 5.77 9.425 5.94 ;
      RECT 9.25 1.36 9.42 1.53 ;
      RECT 9.24 6.63 9.41 6.8 ;
      RECT 9.225 5.14 9.395 5.31 ;
      RECT 8.97 2.11 9.185 2.24 ;
      RECT 8.97 5.89 9.185 6.02 ;
      RECT 8.05 0.165 8.35 0.435 ;
      RECT 8.05 3.945 8.35 4.215 ;
      RECT 8.05 7.725 8.35 7.995 ;
      RECT 7.205 2.15 7.44 2.28 ;
      RECT 7.205 5.93 7.44 6.06 ;
      RECT 7 1.35 7.17 1.52 ;
      RECT 7 5.13 7.17 5.3 ;
      RECT 6.975 2.865 7.145 3.035 ;
      RECT 6.975 6.645 7.145 6.815 ;
      RECT 6.965 2.22 7.135 2.39 ;
      RECT 6.965 6.005 7.135 6.175 ;
      RECT 6.825 2.58 6.995 2.75 ;
      RECT 6.825 6.345 6.995 6.515 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.73 5.315 6.9 5.485 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.34 5.165 6.51 5.335 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 6.12 2.87 6.29 3.04 ;
      RECT 6.12 6.65 6.29 6.82 ;
      RECT 6.06 5.87 6.23 6.04 ;
      RECT 5.73 2.71 5.9 2.88 ;
      RECT 5.73 6.49 5.9 6.66 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.62 5.415 5.79 5.585 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 5.475 5.77 5.645 5.94 ;
      RECT 5.47 1.36 5.64 1.53 ;
      RECT 5.47 5.14 5.64 5.31 ;
      RECT 5.46 2.85 5.63 3.02 ;
      RECT 5.46 6.63 5.63 6.8 ;
      RECT 5.19 2.11 5.405 2.24 ;
      RECT 5.19 5.89 5.405 6.02 ;
      RECT 4.27 0.165 4.57 0.435 ;
      RECT 4.27 3.945 4.57 4.215 ;
      RECT 4.27 7.725 4.57 7.995 ;
      RECT 3.425 2.15 3.66 2.28 ;
      RECT 3.425 5.93 3.66 6.06 ;
      RECT 3.22 1.35 3.39 1.52 ;
      RECT 3.22 5.13 3.39 5.3 ;
      RECT 3.195 2.865 3.365 3.035 ;
      RECT 3.195 6.645 3.365 6.815 ;
      RECT 3.185 2.22 3.355 2.39 ;
      RECT 3.185 6.005 3.355 6.175 ;
      RECT 3.045 2.58 3.215 2.75 ;
      RECT 3.045 6.345 3.215 6.515 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.95 5.315 3.12 5.485 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.56 5.165 2.73 5.335 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 2.34 2.87 2.51 3.04 ;
      RECT 2.34 6.65 2.51 6.82 ;
      RECT 2.28 5.87 2.45 6.04 ;
      RECT 1.95 2.71 2.12 2.88 ;
      RECT 1.95 6.49 2.12 6.66 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.84 5.415 2.01 5.585 ;
      RECT 1.695 1.99 1.865 2.16 ;
      RECT 1.695 5.77 1.865 5.94 ;
      RECT 1.69 1.36 1.86 1.53 ;
      RECT 1.69 5.14 1.86 5.31 ;
      RECT 1.68 2.85 1.85 3.02 ;
      RECT 1.68 6.63 1.85 6.8 ;
      RECT 1.41 2.11 1.625 2.24 ;
      RECT 1.41 5.89 1.625 6.02 ;
      RECT 0.49 0.165 0.79 0.435 ;
      RECT 0.49 3.945 0.79 4.215 ;
      RECT 0.49 7.725 0.79 7.995 ;
    LAYER M10 ;
      RECT 16.26 3.375 19.04 3.58 ;
      RECT 18.83 0.8 19.04 3.58 ;
      RECT 17.75 3.075 19.04 3.58 ;
      RECT 18.53 2.335 19.04 3.58 ;
      RECT 16.26 3.07 17.5 3.58 ;
      RECT 16.26 3.07 17.505 3.22 ;
      RECT 17.655 1.57 18.01 3.125 ;
      RECT 16.26 3.07 18.28 3.125 ;
      RECT 17.75 2.785 18.28 3.58 ;
      RECT 16.26 3.065 17.405 3.58 ;
      RECT 17.305 0.8 17.405 3.58 ;
      RECT 17.02 2.91 17.405 3.58 ;
      RECT 16.26 2.295 16.77 3.58 ;
      RECT 17.02 1.845 17.055 3.58 ;
      RECT 17.655 2.785 19.04 2.825 ;
      RECT 18.525 1.555 18.58 2.825 ;
      RECT 17.305 1.26 17.655 2.82 ;
      RECT 16.26 2.295 17.055 2.815 ;
      RECT 18.37 2.435 19.04 2.825 ;
      RECT 17.305 1.715 18.12 2.82 ;
      RECT 16.26 2.295 18.12 2.66 ;
      RECT 17.17 0.8 17.555 2.66 ;
      RECT 16.26 2.435 19.04 2.535 ;
      RECT 16.715 2.2 18.275 2.535 ;
      RECT 17.17 1.715 18.275 2.535 ;
      RECT 16.26 0.8 16.465 3.58 ;
      RECT 17.015 1.845 18.275 2.535 ;
      RECT 16.715 1.565 16.765 3.58 ;
      RECT 18.26 1.555 18.58 2.185 ;
      RECT 18.54 0.8 19.04 2.085 ;
      RECT 16.26 0.8 16.76 2.045 ;
      RECT 16.26 1.845 19.04 1.95 ;
      RECT 16.26 1.565 16.92 1.95 ;
      RECT 17.01 0.8 17.555 1.595 ;
      RECT 17.905 0.8 18.01 3.58 ;
      RECT 16.26 1.565 17.655 1.595 ;
      RECT 18.26 0.8 18.29 2.185 ;
      RECT 17.905 0.8 18.29 1.465 ;
      RECT 17.01 1.26 18.29 1.32 ;
      RECT 16.26 0.8 17.555 1.315 ;
      RECT 17.805 0.8 19.04 1.305 ;
      RECT 17.795 1.16 19.04 1.305 ;
      RECT 16.26 0.8 19.04 1.01 ;
      RECT 16.26 7.155 19.04 7.36 ;
      RECT 18.83 4.58 19.04 7.36 ;
      RECT 17.75 6.855 19.04 7.36 ;
      RECT 18.53 6.115 19.04 7.36 ;
      RECT 16.26 6.85 17.5 7.36 ;
      RECT 16.26 6.85 17.505 7 ;
      RECT 17.655 5.35 18.01 6.905 ;
      RECT 16.26 6.85 18.28 6.905 ;
      RECT 17.75 6.565 18.28 7.36 ;
      RECT 16.26 6.845 17.405 7.36 ;
      RECT 17.305 4.58 17.405 7.36 ;
      RECT 17.02 6.69 17.405 7.36 ;
      RECT 16.26 6.075 16.77 7.36 ;
      RECT 17.02 5.625 17.055 7.36 ;
      RECT 17.655 6.565 19.04 6.605 ;
      RECT 18.525 5.335 18.58 6.605 ;
      RECT 17.305 5.04 17.655 6.6 ;
      RECT 16.26 6.075 17.055 6.595 ;
      RECT 18.37 6.215 19.04 6.605 ;
      RECT 17.305 5.495 18.12 6.6 ;
      RECT 16.26 6.075 18.12 6.44 ;
      RECT 17.17 4.58 17.555 6.44 ;
      RECT 16.26 6.215 19.04 6.315 ;
      RECT 16.715 5.98 18.275 6.315 ;
      RECT 17.17 5.495 18.275 6.315 ;
      RECT 16.26 4.58 16.465 7.36 ;
      RECT 17.015 5.625 18.275 6.315 ;
      RECT 16.715 5.345 16.765 7.36 ;
      RECT 18.26 5.335 18.58 5.965 ;
      RECT 18.54 4.58 19.04 5.865 ;
      RECT 16.26 4.58 16.76 5.825 ;
      RECT 16.26 5.625 19.04 5.73 ;
      RECT 16.26 5.345 16.92 5.73 ;
      RECT 17.01 4.58 17.555 5.375 ;
      RECT 17.905 4.58 18.01 7.36 ;
      RECT 16.26 5.345 17.655 5.375 ;
      RECT 18.26 4.58 18.29 5.965 ;
      RECT 17.905 4.58 18.29 5.245 ;
      RECT 17.01 5.04 18.29 5.1 ;
      RECT 16.26 4.58 17.555 5.095 ;
      RECT 17.805 4.58 19.04 5.085 ;
      RECT 17.795 4.94 19.04 5.085 ;
      RECT 16.26 4.58 19.04 4.79 ;
      RECT 12.48 3.375 15.26 3.58 ;
      RECT 15.05 0.8 15.26 3.58 ;
      RECT 13.97 3.075 15.26 3.58 ;
      RECT 14.75 2.335 15.26 3.58 ;
      RECT 12.48 3.07 13.72 3.58 ;
      RECT 12.48 3.07 13.725 3.22 ;
      RECT 13.875 1.57 14.23 3.125 ;
      RECT 12.48 3.07 14.5 3.125 ;
      RECT 13.97 2.785 14.5 3.58 ;
      RECT 12.48 3.065 13.625 3.58 ;
      RECT 13.525 0.8 13.625 3.58 ;
      RECT 13.24 2.91 13.625 3.58 ;
      RECT 12.48 2.295 12.99 3.58 ;
      RECT 13.24 1.845 13.275 3.58 ;
      RECT 13.875 2.785 15.26 2.825 ;
      RECT 14.745 1.555 14.8 2.825 ;
      RECT 13.525 1.26 13.875 2.82 ;
      RECT 12.48 2.295 13.275 2.815 ;
      RECT 14.59 2.435 15.26 2.825 ;
      RECT 13.525 1.715 14.34 2.82 ;
      RECT 12.48 2.295 14.34 2.66 ;
      RECT 13.39 0.8 13.775 2.66 ;
      RECT 12.48 2.435 15.26 2.535 ;
      RECT 12.935 2.2 14.495 2.535 ;
      RECT 13.39 1.715 14.495 2.535 ;
      RECT 12.48 0.8 12.685 3.58 ;
      RECT 13.235 1.845 14.495 2.535 ;
      RECT 12.935 1.565 12.985 3.58 ;
      RECT 14.48 1.555 14.8 2.185 ;
      RECT 14.76 0.8 15.26 2.085 ;
      RECT 12.48 0.8 12.98 2.045 ;
      RECT 12.48 1.845 15.26 1.95 ;
      RECT 12.48 1.565 13.14 1.95 ;
      RECT 13.23 0.8 13.775 1.595 ;
      RECT 14.125 0.8 14.23 3.58 ;
      RECT 12.48 1.565 13.875 1.595 ;
      RECT 14.48 0.8 14.51 2.185 ;
      RECT 14.125 0.8 14.51 1.465 ;
      RECT 13.23 1.26 14.51 1.32 ;
      RECT 12.48 0.8 13.775 1.315 ;
      RECT 14.025 0.8 15.26 1.305 ;
      RECT 14.015 1.16 15.26 1.305 ;
      RECT 12.48 0.8 15.26 1.01 ;
      RECT 12.48 7.155 15.26 7.36 ;
      RECT 15.05 4.58 15.26 7.36 ;
      RECT 13.97 6.855 15.26 7.36 ;
      RECT 14.75 6.115 15.26 7.36 ;
      RECT 12.48 6.85 13.72 7.36 ;
      RECT 12.48 6.85 13.725 7 ;
      RECT 13.875 5.35 14.23 6.905 ;
      RECT 12.48 6.85 14.5 6.905 ;
      RECT 13.97 6.565 14.5 7.36 ;
      RECT 12.48 6.845 13.625 7.36 ;
      RECT 13.525 4.58 13.625 7.36 ;
      RECT 13.24 6.69 13.625 7.36 ;
      RECT 12.48 6.075 12.99 7.36 ;
      RECT 13.24 5.625 13.275 7.36 ;
      RECT 13.875 6.565 15.26 6.605 ;
      RECT 14.745 5.335 14.8 6.605 ;
      RECT 13.525 5.04 13.875 6.6 ;
      RECT 12.48 6.075 13.275 6.595 ;
      RECT 14.59 6.215 15.26 6.605 ;
      RECT 13.525 5.495 14.34 6.6 ;
      RECT 12.48 6.075 14.34 6.44 ;
      RECT 13.39 4.58 13.775 6.44 ;
      RECT 12.48 6.215 15.26 6.315 ;
      RECT 12.935 5.98 14.495 6.315 ;
      RECT 13.39 5.495 14.495 6.315 ;
      RECT 12.48 4.58 12.685 7.36 ;
      RECT 13.235 5.625 14.495 6.315 ;
      RECT 12.935 5.345 12.985 7.36 ;
      RECT 14.48 5.335 14.8 5.965 ;
      RECT 14.76 4.58 15.26 5.865 ;
      RECT 12.48 4.58 12.98 5.825 ;
      RECT 12.48 5.625 15.26 5.73 ;
      RECT 12.48 5.345 13.14 5.73 ;
      RECT 13.23 4.58 13.775 5.375 ;
      RECT 14.125 4.58 14.23 7.36 ;
      RECT 12.48 5.345 13.875 5.375 ;
      RECT 14.48 4.58 14.51 5.965 ;
      RECT 14.125 4.58 14.51 5.245 ;
      RECT 13.23 5.04 14.51 5.1 ;
      RECT 12.48 4.58 13.775 5.095 ;
      RECT 14.025 4.58 15.26 5.085 ;
      RECT 14.015 4.94 15.26 5.085 ;
      RECT 12.48 4.58 15.26 4.79 ;
      RECT 8.7 3.375 11.48 3.58 ;
      RECT 11.27 0.8 11.48 3.58 ;
      RECT 10.19 3.075 11.48 3.58 ;
      RECT 10.97 2.335 11.48 3.58 ;
      RECT 8.7 3.07 9.94 3.58 ;
      RECT 8.7 3.07 9.945 3.22 ;
      RECT 10.095 1.57 10.45 3.125 ;
      RECT 8.7 3.07 10.72 3.125 ;
      RECT 10.19 2.785 10.72 3.58 ;
      RECT 8.7 3.065 9.845 3.58 ;
      RECT 9.745 0.8 9.845 3.58 ;
      RECT 9.46 2.91 9.845 3.58 ;
      RECT 8.7 2.295 9.21 3.58 ;
      RECT 9.46 1.845 9.495 3.58 ;
      RECT 10.095 2.785 11.48 2.825 ;
      RECT 10.965 1.555 11.02 2.825 ;
      RECT 9.745 1.26 10.095 2.82 ;
      RECT 8.7 2.295 9.495 2.815 ;
      RECT 10.81 2.435 11.48 2.825 ;
      RECT 9.745 1.715 10.56 2.82 ;
      RECT 8.7 2.295 10.56 2.66 ;
      RECT 9.61 0.8 9.995 2.66 ;
      RECT 8.7 2.435 11.48 2.535 ;
      RECT 9.155 2.2 10.715 2.535 ;
      RECT 9.61 1.715 10.715 2.535 ;
      RECT 8.7 0.8 8.905 3.58 ;
      RECT 9.455 1.845 10.715 2.535 ;
      RECT 9.155 1.565 9.205 3.58 ;
      RECT 10.7 1.555 11.02 2.185 ;
      RECT 10.98 0.8 11.48 2.085 ;
      RECT 8.7 0.8 9.2 2.045 ;
      RECT 8.7 1.845 11.48 1.95 ;
      RECT 8.7 1.565 9.36 1.95 ;
      RECT 9.45 0.8 9.995 1.595 ;
      RECT 10.345 0.8 10.45 3.58 ;
      RECT 8.7 1.565 10.095 1.595 ;
      RECT 10.7 0.8 10.73 2.185 ;
      RECT 10.345 0.8 10.73 1.465 ;
      RECT 9.45 1.26 10.73 1.32 ;
      RECT 8.7 0.8 9.995 1.315 ;
      RECT 10.245 0.8 11.48 1.305 ;
      RECT 10.235 1.16 11.48 1.305 ;
      RECT 8.7 0.8 11.48 1.01 ;
      RECT 8.7 7.155 11.48 7.36 ;
      RECT 11.27 4.58 11.48 7.36 ;
      RECT 10.19 6.855 11.48 7.36 ;
      RECT 10.97 6.115 11.48 7.36 ;
      RECT 8.7 6.85 9.94 7.36 ;
      RECT 8.7 6.85 9.945 7 ;
      RECT 10.095 5.35 10.45 6.905 ;
      RECT 8.7 6.85 10.72 6.905 ;
      RECT 10.19 6.565 10.72 7.36 ;
      RECT 8.7 6.845 9.845 7.36 ;
      RECT 9.745 4.58 9.845 7.36 ;
      RECT 9.46 6.69 9.845 7.36 ;
      RECT 8.7 6.075 9.21 7.36 ;
      RECT 9.46 5.625 9.495 7.36 ;
      RECT 10.095 6.565 11.48 6.605 ;
      RECT 10.965 5.335 11.02 6.605 ;
      RECT 9.745 5.04 10.095 6.6 ;
      RECT 8.7 6.075 9.495 6.595 ;
      RECT 10.81 6.215 11.48 6.605 ;
      RECT 9.745 5.495 10.56 6.6 ;
      RECT 8.7 6.075 10.56 6.44 ;
      RECT 9.61 4.58 9.995 6.44 ;
      RECT 8.7 6.215 11.48 6.315 ;
      RECT 9.155 5.98 10.715 6.315 ;
      RECT 9.61 5.495 10.715 6.315 ;
      RECT 8.7 4.58 8.905 7.36 ;
      RECT 9.455 5.625 10.715 6.315 ;
      RECT 9.155 5.345 9.205 7.36 ;
      RECT 10.7 5.335 11.02 5.965 ;
      RECT 10.98 4.58 11.48 5.865 ;
      RECT 8.7 4.58 9.2 5.825 ;
      RECT 8.7 5.625 11.48 5.73 ;
      RECT 8.7 5.345 9.36 5.73 ;
      RECT 9.45 4.58 9.995 5.375 ;
      RECT 10.345 4.58 10.45 7.36 ;
      RECT 8.7 5.345 10.095 5.375 ;
      RECT 10.7 4.58 10.73 5.965 ;
      RECT 10.345 4.58 10.73 5.245 ;
      RECT 9.45 5.04 10.73 5.1 ;
      RECT 8.7 4.58 9.995 5.095 ;
      RECT 10.245 4.58 11.48 5.085 ;
      RECT 10.235 4.94 11.48 5.085 ;
      RECT 8.7 4.58 11.48 4.79 ;
      RECT 9.25 5.145 9.4 5.295 ;
      RECT 9.245 5.16 9.4 5.29 ;
      RECT 4.92 3.375 7.7 3.58 ;
      RECT 7.49 0.8 7.7 3.58 ;
      RECT 6.41 3.075 7.7 3.58 ;
      RECT 7.19 2.335 7.7 3.58 ;
      RECT 4.92 3.07 6.16 3.58 ;
      RECT 4.92 3.07 6.165 3.22 ;
      RECT 6.315 1.57 6.67 3.125 ;
      RECT 4.92 3.07 6.94 3.125 ;
      RECT 6.41 2.785 6.94 3.58 ;
      RECT 4.92 3.065 6.065 3.58 ;
      RECT 5.965 0.8 6.065 3.58 ;
      RECT 5.68 2.91 6.065 3.58 ;
      RECT 4.92 2.295 5.43 3.58 ;
      RECT 5.68 1.845 5.715 3.58 ;
      RECT 6.315 2.785 7.7 2.825 ;
      RECT 7.185 1.555 7.24 2.825 ;
      RECT 5.965 1.26 6.315 2.82 ;
      RECT 4.92 2.295 5.715 2.815 ;
      RECT 7.03 2.435 7.7 2.825 ;
      RECT 5.965 1.715 6.78 2.82 ;
      RECT 4.92 2.295 6.78 2.66 ;
      RECT 5.83 0.8 6.215 2.66 ;
      RECT 4.92 2.435 7.7 2.535 ;
      RECT 5.375 2.2 6.935 2.535 ;
      RECT 5.83 1.715 6.935 2.535 ;
      RECT 4.92 0.8 5.125 3.58 ;
      RECT 5.675 1.845 6.935 2.535 ;
      RECT 5.375 1.565 5.425 3.58 ;
      RECT 6.92 1.555 7.24 2.185 ;
      RECT 7.2 0.8 7.7 2.085 ;
      RECT 4.92 0.8 5.42 2.045 ;
      RECT 4.92 1.845 7.7 1.95 ;
      RECT 4.92 1.565 5.58 1.95 ;
      RECT 5.67 0.8 6.215 1.595 ;
      RECT 6.565 0.8 6.67 3.58 ;
      RECT 4.92 1.565 6.315 1.595 ;
      RECT 6.92 0.8 6.95 2.185 ;
      RECT 6.565 0.8 6.95 1.465 ;
      RECT 5.67 1.26 6.95 1.32 ;
      RECT 4.92 0.8 6.215 1.315 ;
      RECT 6.465 0.8 7.7 1.305 ;
      RECT 6.455 1.16 7.7 1.305 ;
      RECT 4.92 0.8 7.7 1.01 ;
      RECT 4.92 7.155 7.7 7.36 ;
      RECT 7.49 4.58 7.7 7.36 ;
      RECT 6.41 6.855 7.7 7.36 ;
      RECT 7.19 6.115 7.7 7.36 ;
      RECT 4.92 6.85 6.16 7.36 ;
      RECT 4.92 6.85 6.165 7 ;
      RECT 6.315 5.35 6.67 6.905 ;
      RECT 4.92 6.85 6.94 6.905 ;
      RECT 6.41 6.565 6.94 7.36 ;
      RECT 4.92 6.845 6.065 7.36 ;
      RECT 5.965 4.58 6.065 7.36 ;
      RECT 5.68 6.69 6.065 7.36 ;
      RECT 4.92 6.075 5.43 7.36 ;
      RECT 5.68 5.625 5.715 7.36 ;
      RECT 6.315 6.565 7.7 6.605 ;
      RECT 7.185 5.335 7.24 6.605 ;
      RECT 5.965 5.04 6.315 6.6 ;
      RECT 4.92 6.075 5.715 6.595 ;
      RECT 7.03 6.215 7.7 6.605 ;
      RECT 5.965 5.495 6.78 6.6 ;
      RECT 4.92 6.075 6.78 6.44 ;
      RECT 5.83 4.58 6.215 6.44 ;
      RECT 4.92 6.215 7.7 6.315 ;
      RECT 5.375 5.98 6.935 6.315 ;
      RECT 5.83 5.495 6.935 6.315 ;
      RECT 4.92 4.58 5.125 7.36 ;
      RECT 5.675 5.625 6.935 6.315 ;
      RECT 5.375 5.345 5.425 7.36 ;
      RECT 6.92 5.335 7.24 5.965 ;
      RECT 7.2 4.58 7.7 5.865 ;
      RECT 4.92 4.58 5.42 5.825 ;
      RECT 4.92 5.625 7.7 5.73 ;
      RECT 4.92 5.345 5.58 5.73 ;
      RECT 5.67 4.58 6.215 5.375 ;
      RECT 6.565 4.58 6.67 7.36 ;
      RECT 4.92 5.345 6.315 5.375 ;
      RECT 6.92 4.58 6.95 5.965 ;
      RECT 6.565 4.58 6.95 5.245 ;
      RECT 5.67 5.04 6.95 5.1 ;
      RECT 4.92 4.58 6.215 5.095 ;
      RECT 6.465 4.58 7.7 5.085 ;
      RECT 6.455 4.94 7.7 5.085 ;
      RECT 4.92 4.58 7.7 4.79 ;
      RECT 1.14 3.375 3.92 3.58 ;
      RECT 3.71 0.8 3.92 3.58 ;
      RECT 2.63 3.075 3.92 3.58 ;
      RECT 3.41 2.335 3.92 3.58 ;
      RECT 1.14 3.07 2.38 3.58 ;
      RECT 1.14 3.07 2.385 3.22 ;
      RECT 2.535 1.57 2.89 3.125 ;
      RECT 1.14 3.07 3.16 3.125 ;
      RECT 2.63 2.785 3.16 3.58 ;
      RECT 1.14 3.065 2.285 3.58 ;
      RECT 2.185 0.8 2.285 3.58 ;
      RECT 1.9 2.91 2.285 3.58 ;
      RECT 1.14 2.295 1.65 3.58 ;
      RECT 1.9 1.845 1.935 3.58 ;
      RECT 2.535 2.785 3.92 2.825 ;
      RECT 3.405 1.555 3.46 2.825 ;
      RECT 2.185 1.26 2.535 2.82 ;
      RECT 1.14 2.295 1.935 2.815 ;
      RECT 3.25 2.435 3.92 2.825 ;
      RECT 2.185 1.715 3 2.82 ;
      RECT 1.14 2.295 3 2.66 ;
      RECT 2.05 0.8 2.435 2.66 ;
      RECT 1.14 2.435 3.92 2.535 ;
      RECT 1.595 2.2 3.155 2.535 ;
      RECT 2.05 1.715 3.155 2.535 ;
      RECT 1.14 0.8 1.345 3.58 ;
      RECT 1.895 1.845 3.155 2.535 ;
      RECT 1.595 1.565 1.645 3.58 ;
      RECT 3.14 1.555 3.46 2.185 ;
      RECT 3.42 0.8 3.92 2.085 ;
      RECT 1.14 0.8 1.64 2.045 ;
      RECT 1.14 1.845 3.92 1.95 ;
      RECT 1.14 1.565 1.8 1.95 ;
      RECT 1.89 0.8 2.435 1.595 ;
      RECT 2.785 0.8 2.89 3.58 ;
      RECT 1.14 1.565 2.535 1.595 ;
      RECT 3.14 0.8 3.17 2.185 ;
      RECT 2.785 0.8 3.17 1.465 ;
      RECT 1.89 1.26 3.17 1.32 ;
      RECT 1.14 0.8 2.435 1.315 ;
      RECT 2.685 0.8 3.92 1.305 ;
      RECT 2.675 1.16 3.92 1.305 ;
      RECT 1.14 0.8 3.92 1.01 ;
      RECT 1.14 7.155 3.92 7.36 ;
      RECT 3.71 4.58 3.92 7.36 ;
      RECT 2.63 6.855 3.92 7.36 ;
      RECT 3.41 6.115 3.92 7.36 ;
      RECT 1.14 6.85 2.38 7.36 ;
      RECT 1.14 6.85 2.385 7 ;
      RECT 2.535 5.35 2.89 6.905 ;
      RECT 1.14 6.85 3.16 6.905 ;
      RECT 2.63 6.565 3.16 7.36 ;
      RECT 1.14 6.845 2.285 7.36 ;
      RECT 2.185 4.58 2.285 7.36 ;
      RECT 1.9 6.69 2.285 7.36 ;
      RECT 1.14 6.075 1.65 7.36 ;
      RECT 1.9 5.625 1.935 7.36 ;
      RECT 2.535 6.565 3.92 6.605 ;
      RECT 3.405 5.335 3.46 6.605 ;
      RECT 2.185 5.04 2.535 6.6 ;
      RECT 1.14 6.075 1.935 6.595 ;
      RECT 3.25 6.215 3.92 6.605 ;
      RECT 2.185 5.495 3 6.6 ;
      RECT 1.14 6.075 3 6.44 ;
      RECT 2.05 4.58 2.435 6.44 ;
      RECT 1.14 6.215 3.92 6.315 ;
      RECT 1.595 5.98 3.155 6.315 ;
      RECT 2.05 5.495 3.155 6.315 ;
      RECT 1.14 4.58 1.345 7.36 ;
      RECT 1.895 5.625 3.155 6.315 ;
      RECT 1.595 5.345 1.645 7.36 ;
      RECT 3.14 5.335 3.46 5.965 ;
      RECT 3.42 4.58 3.92 5.865 ;
      RECT 1.14 4.58 1.64 5.825 ;
      RECT 1.14 5.625 3.92 5.73 ;
      RECT 1.14 5.345 1.8 5.73 ;
      RECT 1.89 4.58 2.435 5.375 ;
      RECT 2.785 4.58 2.89 7.36 ;
      RECT 1.14 5.345 2.535 5.375 ;
      RECT 3.14 4.58 3.17 5.965 ;
      RECT 2.785 4.58 3.17 5.245 ;
      RECT 1.89 5.04 3.17 5.1 ;
      RECT 1.14 4.58 2.435 5.095 ;
      RECT 2.685 4.58 3.92 5.085 ;
      RECT 2.675 4.94 3.92 5.085 ;
      RECT 1.14 4.58 3.92 4.79 ;
      RECT 19.34 0.1 19.74 0.5 ;
      RECT 19.34 3.88 19.74 4.28 ;
      RECT 19.34 7.66 19.74 8.06 ;
      RECT 18.63 2.135 18.78 2.285 ;
      RECT 18.63 5.915 18.78 6.065 ;
      RECT 18.34 1.354 18.49 1.504 ;
      RECT 18.34 5.134 18.49 5.284 ;
      RECT 18.331 2.873 18.481 3.023 ;
      RECT 18.331 6.653 18.481 6.803 ;
      RECT 18.325 2.236 18.475 2.386 ;
      RECT 18.325 6.016 18.475 6.166 ;
      RECT 18.172 2.584 18.322 2.734 ;
      RECT 18.172 6.364 18.322 6.514 ;
      RECT 18.058 1.517 18.208 1.667 ;
      RECT 18.058 5.297 18.208 5.447 ;
      RECT 17.706 1.368 17.856 1.518 ;
      RECT 17.706 5.148 17.856 5.298 ;
      RECT 17.604 1.061 17.754 1.211 ;
      RECT 17.604 4.841 17.754 4.991 ;
      RECT 17.551 3.173 17.701 3.323 ;
      RECT 17.551 6.953 17.701 7.103 ;
      RECT 17.455 2.87 17.605 3.02 ;
      RECT 17.455 6.65 17.605 6.8 ;
      RECT 17.104 2.708 17.254 2.858 ;
      RECT 17.104 6.488 17.254 6.638 ;
      RECT 16.97 1.643 17.12 1.793 ;
      RECT 16.97 5.423 17.12 5.573 ;
      RECT 16.818 2.866 16.968 3.016 ;
      RECT 16.818 6.646 16.968 6.796 ;
      RECT 16.817 1.998 16.967 2.148 ;
      RECT 16.817 5.778 16.967 5.928 ;
      RECT 16.81 1.363 16.96 1.513 ;
      RECT 16.81 5.143 16.96 5.293 ;
      RECT 16.513 2.096 16.663 2.246 ;
      RECT 16.513 5.876 16.663 6.026 ;
      RECT 15.56 0.1 15.96 0.5 ;
      RECT 15.56 3.88 15.96 4.28 ;
      RECT 15.56 7.66 15.96 8.06 ;
      RECT 14.85 2.135 15 2.285 ;
      RECT 14.85 5.915 15 6.065 ;
      RECT 14.56 1.354 14.71 1.504 ;
      RECT 14.56 5.134 14.71 5.284 ;
      RECT 14.551 2.873 14.701 3.023 ;
      RECT 14.551 6.653 14.701 6.803 ;
      RECT 14.545 2.236 14.695 2.386 ;
      RECT 14.545 6.016 14.695 6.166 ;
      RECT 14.392 2.584 14.542 2.734 ;
      RECT 14.392 6.364 14.542 6.514 ;
      RECT 14.278 1.517 14.428 1.667 ;
      RECT 14.278 5.297 14.428 5.447 ;
      RECT 13.926 1.368 14.076 1.518 ;
      RECT 13.926 5.148 14.076 5.298 ;
      RECT 13.824 1.061 13.974 1.211 ;
      RECT 13.824 4.841 13.974 4.991 ;
      RECT 13.771 3.173 13.921 3.323 ;
      RECT 13.771 6.953 13.921 7.103 ;
      RECT 13.675 2.87 13.825 3.02 ;
      RECT 13.675 6.65 13.825 6.8 ;
      RECT 13.324 2.708 13.474 2.858 ;
      RECT 13.324 6.488 13.474 6.638 ;
      RECT 13.19 1.643 13.34 1.793 ;
      RECT 13.19 5.423 13.34 5.573 ;
      RECT 13.038 2.866 13.188 3.016 ;
      RECT 13.038 6.646 13.188 6.796 ;
      RECT 13.037 1.998 13.187 2.148 ;
      RECT 13.037 5.778 13.187 5.928 ;
      RECT 13.03 1.363 13.18 1.513 ;
      RECT 13.03 5.143 13.18 5.293 ;
      RECT 12.733 2.096 12.883 2.246 ;
      RECT 12.733 5.876 12.883 6.026 ;
      RECT 11.78 0.1 12.18 0.5 ;
      RECT 11.78 3.88 12.18 4.28 ;
      RECT 11.78 7.66 12.18 8.06 ;
      RECT 11.07 2.135 11.22 2.285 ;
      RECT 11.07 5.915 11.22 6.065 ;
      RECT 10.78 1.354 10.93 1.504 ;
      RECT 10.78 5.134 10.93 5.284 ;
      RECT 10.771 2.873 10.921 3.023 ;
      RECT 10.771 6.653 10.921 6.803 ;
      RECT 10.765 2.236 10.915 2.386 ;
      RECT 10.765 6.016 10.915 6.166 ;
      RECT 10.612 2.584 10.762 2.734 ;
      RECT 10.612 6.364 10.762 6.514 ;
      RECT 10.498 1.517 10.648 1.667 ;
      RECT 10.498 5.297 10.648 5.447 ;
      RECT 10.146 1.368 10.296 1.518 ;
      RECT 10.146 5.148 10.296 5.298 ;
      RECT 10.044 1.061 10.194 1.211 ;
      RECT 10.044 4.841 10.194 4.991 ;
      RECT 9.991 3.173 10.141 3.323 ;
      RECT 9.991 6.953 10.141 7.103 ;
      RECT 9.895 2.87 10.045 3.02 ;
      RECT 9.895 6.65 10.045 6.8 ;
      RECT 9.544 2.708 9.694 2.858 ;
      RECT 9.544 6.488 9.694 6.638 ;
      RECT 9.41 1.643 9.56 1.793 ;
      RECT 9.41 5.423 9.56 5.573 ;
      RECT 9.258 2.866 9.408 3.016 ;
      RECT 9.258 6.646 9.408 6.796 ;
      RECT 9.257 1.998 9.407 2.148 ;
      RECT 9.257 5.778 9.407 5.928 ;
      RECT 9.25 1.363 9.4 1.513 ;
      RECT 8.953 2.096 9.103 2.246 ;
      RECT 8.953 5.876 9.103 6.026 ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 8 7.66 8.4 8.06 ;
      RECT 7.29 2.135 7.44 2.285 ;
      RECT 7.29 5.915 7.44 6.065 ;
      RECT 7 1.354 7.15 1.504 ;
      RECT 7 5.134 7.15 5.284 ;
      RECT 6.991 2.873 7.141 3.023 ;
      RECT 6.991 6.653 7.141 6.803 ;
      RECT 6.985 2.236 7.135 2.386 ;
      RECT 6.985 6.016 7.135 6.166 ;
      RECT 6.832 2.584 6.982 2.734 ;
      RECT 6.832 6.364 6.982 6.514 ;
      RECT 6.718 1.517 6.868 1.667 ;
      RECT 6.718 5.297 6.868 5.447 ;
      RECT 6.366 1.368 6.516 1.518 ;
      RECT 6.366 5.148 6.516 5.298 ;
      RECT 6.264 1.061 6.414 1.211 ;
      RECT 6.264 4.841 6.414 4.991 ;
      RECT 6.211 3.173 6.361 3.323 ;
      RECT 6.211 6.953 6.361 7.103 ;
      RECT 6.115 2.87 6.265 3.02 ;
      RECT 6.115 6.65 6.265 6.8 ;
      RECT 5.764 2.708 5.914 2.858 ;
      RECT 5.764 6.488 5.914 6.638 ;
      RECT 5.63 1.643 5.78 1.793 ;
      RECT 5.63 5.423 5.78 5.573 ;
      RECT 5.478 2.866 5.628 3.016 ;
      RECT 5.478 6.646 5.628 6.796 ;
      RECT 5.477 1.998 5.627 2.148 ;
      RECT 5.477 5.778 5.627 5.928 ;
      RECT 5.47 1.363 5.62 1.513 ;
      RECT 5.47 5.143 5.62 5.293 ;
      RECT 5.173 2.096 5.323 2.246 ;
      RECT 5.173 5.876 5.323 6.026 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 4.22 7.66 4.62 8.06 ;
      RECT 3.51 2.135 3.66 2.285 ;
      RECT 3.51 5.915 3.66 6.065 ;
      RECT 3.22 1.354 3.37 1.504 ;
      RECT 3.22 5.134 3.37 5.284 ;
      RECT 3.211 2.873 3.361 3.023 ;
      RECT 3.211 6.653 3.361 6.803 ;
      RECT 3.205 2.236 3.355 2.386 ;
      RECT 3.205 6.016 3.355 6.166 ;
      RECT 3.052 2.584 3.202 2.734 ;
      RECT 3.052 6.364 3.202 6.514 ;
      RECT 2.938 1.517 3.088 1.667 ;
      RECT 2.938 5.297 3.088 5.447 ;
      RECT 2.586 1.368 2.736 1.518 ;
      RECT 2.586 5.148 2.736 5.298 ;
      RECT 2.484 1.061 2.634 1.211 ;
      RECT 2.484 4.841 2.634 4.991 ;
      RECT 2.431 3.173 2.581 3.323 ;
      RECT 2.431 6.953 2.581 7.103 ;
      RECT 2.335 2.87 2.485 3.02 ;
      RECT 2.335 6.65 2.485 6.8 ;
      RECT 1.984 2.708 2.134 2.858 ;
      RECT 1.984 6.488 2.134 6.638 ;
      RECT 1.85 1.643 2 1.793 ;
      RECT 1.85 5.423 2 5.573 ;
      RECT 1.698 2.866 1.848 3.016 ;
      RECT 1.698 6.646 1.848 6.796 ;
      RECT 1.697 1.998 1.847 2.148 ;
      RECT 1.697 5.778 1.847 5.928 ;
      RECT 1.69 1.363 1.84 1.513 ;
      RECT 1.69 5.143 1.84 5.293 ;
      RECT 1.393 2.096 1.543 2.246 ;
      RECT 1.393 5.876 1.543 6.026 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
      RECT 0.44 7.66 0.84 8.06 ;
    LAYER NEMANC ;
      RECT 19.34 0.1 19.74 0.5 ;
      RECT 19.34 3.88 19.74 4.28 ;
      RECT 19.34 7.66 19.74 8.06 ;
      RECT 15.56 0.1 15.96 0.5 ;
      RECT 15.56 3.88 15.96 4.28 ;
      RECT 15.56 7.66 15.96 8.06 ;
      RECT 11.78 0.1 12.18 0.5 ;
      RECT 11.78 3.88 12.18 4.28 ;
      RECT 11.78 7.66 12.18 8.06 ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 8 7.66 8.4 8.06 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 4.22 7.66 4.62 8.06 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
      RECT 0.44 7.66 0.84 8.06 ;
    LAYER NEMCHAN ;
      RECT 18.415 2.22 18.495 2.37 ;
      RECT 18.415 2.22 18.535 2.355 ;
      RECT 18.415 2.22 18.575 2.34 ;
      RECT 18.415 2.22 18.615 2.325 ;
      RECT 18.655 2.14 18.68 2.305 ;
      RECT 18.375 2.23 18.68 2.3 ;
      RECT 18.495 2.195 18.72 2.29 ;
      RECT 18.375 2.26 18.73 2.285 ;
      RECT 18.455 2.205 18.72 2.29 ;
      RECT 18.535 2.18 18.68 2.305 ;
      RECT 18.615 2.155 18.655 2.315 ;
      RECT 18.575 2.165 18.68 2.305 ;
      RECT 18.415 6 18.495 6.15 ;
      RECT 18.415 6 18.535 6.135 ;
      RECT 18.415 6 18.575 6.12 ;
      RECT 18.415 6 18.615 6.105 ;
      RECT 18.655 5.92 18.68 6.085 ;
      RECT 18.375 6.01 18.68 6.08 ;
      RECT 18.495 5.975 18.72 6.07 ;
      RECT 18.375 6.04 18.73 6.065 ;
      RECT 18.455 5.985 18.72 6.07 ;
      RECT 18.535 5.96 18.68 6.085 ;
      RECT 18.615 5.935 18.655 6.095 ;
      RECT 18.575 5.945 18.68 6.085 ;
      RECT 18.34 2.705 18.38 2.975 ;
      RECT 18.3 2.78 18.42 2.95 ;
      RECT 18.3 2.855 18.46 2.93 ;
      RECT 18.3 2.895 18.47 2.915 ;
      RECT 18.26 2.645 18.3 2.88 ;
      RECT 18.22 2.665 18.34 2.805 ;
      RECT 18.18 2.685 18.34 2.735 ;
      RECT 18.26 2.65 18.34 2.88 ;
      RECT 18.34 6.485 18.38 6.755 ;
      RECT 18.3 6.56 18.42 6.73 ;
      RECT 18.3 6.635 18.46 6.71 ;
      RECT 18.3 6.675 18.47 6.695 ;
      RECT 18.26 6.425 18.3 6.66 ;
      RECT 18.22 6.445 18.34 6.585 ;
      RECT 18.18 6.465 18.34 6.515 ;
      RECT 18.26 6.43 18.34 6.66 ;
      RECT 18.175 1.465 18.215 1.64 ;
      RECT 18.135 1.49 18.215 1.625 ;
      RECT 18.135 1.49 18.255 1.62 ;
      RECT 18.135 1.49 18.295 1.595 ;
      RECT 18.095 1.51 18.335 1.565 ;
      RECT 18.335 1.375 18.375 1.55 ;
      RECT 18.335 1.395 18.415 1.525 ;
      RECT 18.175 1.465 18.45 1.51 ;
      RECT 18.215 1.445 18.415 1.525 ;
      RECT 18.295 1.4 18.335 1.57 ;
      RECT 18.255 1.42 18.415 1.525 ;
      RECT 18.175 5.245 18.215 5.42 ;
      RECT 18.135 5.27 18.215 5.405 ;
      RECT 18.135 5.27 18.255 5.4 ;
      RECT 18.135 5.27 18.295 5.375 ;
      RECT 18.095 5.29 18.335 5.345 ;
      RECT 18.335 5.155 18.375 5.33 ;
      RECT 18.335 5.175 18.415 5.305 ;
      RECT 18.175 5.245 18.45 5.29 ;
      RECT 18.215 5.225 18.415 5.305 ;
      RECT 18.295 5.18 18.335 5.35 ;
      RECT 18.255 5.2 18.415 5.305 ;
      RECT 17.73 1.115 17.75 1.46 ;
      RECT 17.73 1.175 17.79 1.445 ;
      RECT 17.69 1.295 17.83 1.435 ;
      RECT 17.69 1.39 17.85 1.425 ;
      RECT 17.65 1.14 17.75 1.345 ;
      RECT 17.61 1.15 17.75 1.22 ;
      RECT 17.69 1.125 17.75 1.435 ;
      RECT 17.73 4.895 17.75 5.24 ;
      RECT 17.73 4.955 17.79 5.225 ;
      RECT 17.69 5.075 17.83 5.215 ;
      RECT 17.69 5.17 17.85 5.205 ;
      RECT 17.65 4.92 17.75 5.125 ;
      RECT 17.61 4.93 17.75 5 ;
      RECT 17.69 4.905 17.75 5.215 ;
      RECT 17.58 2.92 17.6 3.26 ;
      RECT 17.58 2.98 17.64 3.25 ;
      RECT 17.54 3.1 17.68 3.24 ;
      RECT 17.54 3.195 17.7 3.23 ;
      RECT 17.5 2.945 17.6 3.16 ;
      RECT 17.46 2.955 17.6 3.035 ;
      RECT 17.54 2.93 17.6 3.24 ;
      RECT 17.58 6.7 17.6 7.04 ;
      RECT 17.58 6.76 17.64 7.03 ;
      RECT 17.54 6.88 17.68 7.02 ;
      RECT 17.54 6.975 17.7 7.01 ;
      RECT 17.5 6.725 17.6 6.94 ;
      RECT 17.46 6.735 17.6 6.815 ;
      RECT 17.54 6.71 17.6 7.02 ;
      RECT 16.935 2.82 16.975 2.99 ;
      RECT 16.895 2.84 16.975 2.975 ;
      RECT 16.895 2.84 17.015 2.97 ;
      RECT 16.895 2.84 17.095 2.93 ;
      RECT 16.855 2.865 17.095 2.915 ;
      RECT 16.855 2.865 17.135 2.905 ;
      RECT 17.135 2.72 17.145 2.895 ;
      RECT 17.055 2.755 17.185 2.88 ;
      RECT 16.935 2.82 17.215 2.86 ;
      RECT 16.975 2.8 17.185 2.88 ;
      RECT 17.015 2.78 17.055 2.95 ;
      RECT 17.095 2.735 17.145 2.895 ;
      RECT 16.935 6.6 16.975 6.77 ;
      RECT 16.895 6.62 16.975 6.755 ;
      RECT 16.895 6.62 17.015 6.75 ;
      RECT 16.895 6.62 17.095 6.71 ;
      RECT 16.855 6.645 17.095 6.695 ;
      RECT 16.855 6.645 17.135 6.685 ;
      RECT 17.135 6.5 17.145 6.675 ;
      RECT 17.055 6.535 17.185 6.66 ;
      RECT 16.935 6.6 17.215 6.64 ;
      RECT 16.975 6.58 17.185 6.66 ;
      RECT 17.015 6.56 17.055 6.73 ;
      RECT 17.095 6.515 17.145 6.675 ;
      RECT 16.98 1.48 17.02 1.745 ;
      RECT 16.94 1.555 17.06 1.72 ;
      RECT 16.94 1.625 17.1 1.7 ;
      RECT 16.94 1.665 17.11 1.685 ;
      RECT 16.9 1.415 16.94 1.65 ;
      RECT 16.86 1.44 16.98 1.58 ;
      RECT 16.82 1.46 16.98 1.51 ;
      RECT 16.9 1.425 16.98 1.65 ;
      RECT 16.98 5.26 17.02 5.525 ;
      RECT 16.94 5.335 17.06 5.5 ;
      RECT 16.94 5.405 17.1 5.48 ;
      RECT 16.94 5.445 17.11 5.465 ;
      RECT 16.9 5.195 16.94 5.43 ;
      RECT 16.86 5.22 16.98 5.36 ;
      RECT 16.82 5.24 16.98 5.29 ;
      RECT 16.9 5.205 16.98 5.43 ;
      RECT 16.605 2.08 16.645 2.23 ;
      RECT 16.605 2.08 16.685 2.225 ;
      RECT 16.605 2.08 16.725 2.21 ;
      RECT 16.605 2.08 16.765 2.2 ;
      RECT 16.845 2 16.87 2.17 ;
      RECT 16.565 2.09 16.87 2.165 ;
      RECT 16.685 2.06 16.91 2.155 ;
      RECT 16.565 2.135 16.915 2.145 ;
      RECT 16.645 2.065 16.91 2.155 ;
      RECT 16.685 2.055 16.87 2.17 ;
      RECT 16.805 2.015 16.845 2.175 ;
      RECT 16.725 2.04 16.87 2.17 ;
      RECT 16.765 2.025 16.805 2.185 ;
      RECT 16.605 5.86 16.645 6.01 ;
      RECT 16.605 5.86 16.685 6.005 ;
      RECT 16.605 5.86 16.725 5.99 ;
      RECT 16.605 5.86 16.765 5.98 ;
      RECT 16.845 5.78 16.87 5.95 ;
      RECT 16.565 5.87 16.87 5.945 ;
      RECT 16.685 5.84 16.91 5.935 ;
      RECT 16.565 5.915 16.915 5.925 ;
      RECT 16.645 5.845 16.91 5.935 ;
      RECT 16.685 5.835 16.87 5.95 ;
      RECT 16.805 5.795 16.845 5.955 ;
      RECT 16.725 5.82 16.87 5.95 ;
      RECT 16.765 5.805 16.805 5.965 ;
      RECT 14.635 2.22 14.715 2.37 ;
      RECT 14.635 2.22 14.755 2.355 ;
      RECT 14.635 2.22 14.795 2.34 ;
      RECT 14.635 2.22 14.835 2.325 ;
      RECT 14.875 2.14 14.9 2.305 ;
      RECT 14.595 2.23 14.9 2.3 ;
      RECT 14.715 2.195 14.94 2.29 ;
      RECT 14.595 2.26 14.95 2.285 ;
      RECT 14.675 2.205 14.94 2.29 ;
      RECT 14.755 2.18 14.9 2.305 ;
      RECT 14.835 2.155 14.875 2.315 ;
      RECT 14.795 2.165 14.9 2.305 ;
      RECT 14.635 6 14.715 6.15 ;
      RECT 14.635 6 14.755 6.135 ;
      RECT 14.635 6 14.795 6.12 ;
      RECT 14.635 6 14.835 6.105 ;
      RECT 14.875 5.92 14.9 6.085 ;
      RECT 14.595 6.01 14.9 6.08 ;
      RECT 14.715 5.975 14.94 6.07 ;
      RECT 14.595 6.04 14.95 6.065 ;
      RECT 14.675 5.985 14.94 6.07 ;
      RECT 14.755 5.96 14.9 6.085 ;
      RECT 14.835 5.935 14.875 6.095 ;
      RECT 14.795 5.945 14.9 6.085 ;
      RECT 14.56 2.705 14.6 2.975 ;
      RECT 14.52 2.78 14.64 2.95 ;
      RECT 14.52 2.855 14.68 2.93 ;
      RECT 14.52 2.895 14.69 2.915 ;
      RECT 14.48 2.645 14.52 2.88 ;
      RECT 14.44 2.665 14.56 2.805 ;
      RECT 14.4 2.685 14.56 2.735 ;
      RECT 14.48 2.65 14.56 2.88 ;
      RECT 14.56 6.485 14.6 6.755 ;
      RECT 14.52 6.56 14.64 6.73 ;
      RECT 14.52 6.635 14.68 6.71 ;
      RECT 14.52 6.675 14.69 6.695 ;
      RECT 14.48 6.425 14.52 6.66 ;
      RECT 14.44 6.445 14.56 6.585 ;
      RECT 14.4 6.465 14.56 6.515 ;
      RECT 14.48 6.43 14.56 6.66 ;
      RECT 14.395 1.465 14.435 1.64 ;
      RECT 14.355 1.49 14.435 1.625 ;
      RECT 14.355 1.49 14.475 1.62 ;
      RECT 14.355 1.49 14.515 1.595 ;
      RECT 14.315 1.51 14.555 1.565 ;
      RECT 14.555 1.375 14.595 1.55 ;
      RECT 14.555 1.395 14.635 1.525 ;
      RECT 14.395 1.465 14.67 1.51 ;
      RECT 14.435 1.445 14.635 1.525 ;
      RECT 14.515 1.4 14.555 1.57 ;
      RECT 14.475 1.42 14.635 1.525 ;
      RECT 14.395 5.245 14.435 5.42 ;
      RECT 14.355 5.27 14.435 5.405 ;
      RECT 14.355 5.27 14.475 5.4 ;
      RECT 14.355 5.27 14.515 5.375 ;
      RECT 14.315 5.29 14.555 5.345 ;
      RECT 14.555 5.155 14.595 5.33 ;
      RECT 14.555 5.175 14.635 5.305 ;
      RECT 14.395 5.245 14.67 5.29 ;
      RECT 14.435 5.225 14.635 5.305 ;
      RECT 14.515 5.18 14.555 5.35 ;
      RECT 14.475 5.2 14.635 5.305 ;
      RECT 13.95 1.115 13.97 1.46 ;
      RECT 13.95 1.175 14.01 1.445 ;
      RECT 13.91 1.295 14.05 1.435 ;
      RECT 13.91 1.39 14.07 1.425 ;
      RECT 13.87 1.14 13.97 1.345 ;
      RECT 13.83 1.15 13.97 1.22 ;
      RECT 13.91 1.125 13.97 1.435 ;
      RECT 13.95 4.895 13.97 5.24 ;
      RECT 13.95 4.955 14.01 5.225 ;
      RECT 13.91 5.075 14.05 5.215 ;
      RECT 13.91 5.17 14.07 5.205 ;
      RECT 13.87 4.92 13.97 5.125 ;
      RECT 13.83 4.93 13.97 5 ;
      RECT 13.91 4.905 13.97 5.215 ;
      RECT 13.8 2.92 13.82 3.26 ;
      RECT 13.8 2.98 13.86 3.25 ;
      RECT 13.76 3.1 13.9 3.24 ;
      RECT 13.76 3.195 13.92 3.23 ;
      RECT 13.72 2.945 13.82 3.16 ;
      RECT 13.68 2.955 13.82 3.035 ;
      RECT 13.76 2.93 13.82 3.24 ;
      RECT 13.8 6.7 13.82 7.04 ;
      RECT 13.8 6.76 13.86 7.03 ;
      RECT 13.76 6.88 13.9 7.02 ;
      RECT 13.76 6.975 13.92 7.01 ;
      RECT 13.72 6.725 13.82 6.94 ;
      RECT 13.68 6.735 13.82 6.815 ;
      RECT 13.76 6.71 13.82 7.02 ;
      RECT 13.155 2.82 13.195 2.99 ;
      RECT 13.115 2.84 13.195 2.975 ;
      RECT 13.115 2.84 13.235 2.97 ;
      RECT 13.115 2.84 13.315 2.93 ;
      RECT 13.075 2.865 13.315 2.915 ;
      RECT 13.075 2.865 13.355 2.905 ;
      RECT 13.355 2.72 13.365 2.895 ;
      RECT 13.275 2.755 13.405 2.88 ;
      RECT 13.155 2.82 13.435 2.86 ;
      RECT 13.195 2.8 13.405 2.88 ;
      RECT 13.235 2.78 13.275 2.95 ;
      RECT 13.315 2.735 13.365 2.895 ;
      RECT 13.155 6.6 13.195 6.77 ;
      RECT 13.115 6.62 13.195 6.755 ;
      RECT 13.115 6.62 13.235 6.75 ;
      RECT 13.115 6.62 13.315 6.71 ;
      RECT 13.075 6.645 13.315 6.695 ;
      RECT 13.075 6.645 13.355 6.685 ;
      RECT 13.355 6.5 13.365 6.675 ;
      RECT 13.275 6.535 13.405 6.66 ;
      RECT 13.155 6.6 13.435 6.64 ;
      RECT 13.195 6.58 13.405 6.66 ;
      RECT 13.235 6.56 13.275 6.73 ;
      RECT 13.315 6.515 13.365 6.675 ;
      RECT 13.2 1.48 13.24 1.745 ;
      RECT 13.16 1.555 13.28 1.72 ;
      RECT 13.16 1.625 13.32 1.7 ;
      RECT 13.16 1.665 13.33 1.685 ;
      RECT 13.12 1.415 13.16 1.65 ;
      RECT 13.08 1.44 13.2 1.58 ;
      RECT 13.04 1.46 13.2 1.51 ;
      RECT 13.12 1.425 13.2 1.65 ;
      RECT 13.2 5.26 13.24 5.525 ;
      RECT 13.16 5.335 13.28 5.5 ;
      RECT 13.16 5.405 13.32 5.48 ;
      RECT 13.16 5.445 13.33 5.465 ;
      RECT 13.12 5.195 13.16 5.43 ;
      RECT 13.08 5.22 13.2 5.36 ;
      RECT 13.04 5.24 13.2 5.29 ;
      RECT 13.12 5.205 13.2 5.43 ;
      RECT 12.825 2.08 12.865 2.23 ;
      RECT 12.825 2.08 12.905 2.225 ;
      RECT 12.825 2.08 12.945 2.21 ;
      RECT 12.825 2.08 12.985 2.2 ;
      RECT 13.065 2 13.09 2.17 ;
      RECT 12.785 2.09 13.09 2.165 ;
      RECT 12.905 2.06 13.13 2.155 ;
      RECT 12.785 2.135 13.135 2.145 ;
      RECT 12.865 2.065 13.13 2.155 ;
      RECT 12.905 2.055 13.09 2.17 ;
      RECT 13.025 2.015 13.065 2.175 ;
      RECT 12.945 2.04 13.09 2.17 ;
      RECT 12.985 2.025 13.025 2.185 ;
      RECT 12.825 5.86 12.865 6.01 ;
      RECT 12.825 5.86 12.905 6.005 ;
      RECT 12.825 5.86 12.945 5.99 ;
      RECT 12.825 5.86 12.985 5.98 ;
      RECT 13.065 5.78 13.09 5.95 ;
      RECT 12.785 5.87 13.09 5.945 ;
      RECT 12.905 5.84 13.13 5.935 ;
      RECT 12.785 5.915 13.135 5.925 ;
      RECT 12.865 5.845 13.13 5.935 ;
      RECT 12.905 5.835 13.09 5.95 ;
      RECT 13.025 5.795 13.065 5.955 ;
      RECT 12.945 5.82 13.09 5.95 ;
      RECT 12.985 5.805 13.025 5.965 ;
      RECT 10.855 2.22 10.935 2.37 ;
      RECT 10.855 2.22 10.975 2.355 ;
      RECT 10.855 2.22 11.015 2.34 ;
      RECT 10.855 2.22 11.055 2.325 ;
      RECT 11.095 2.14 11.12 2.305 ;
      RECT 10.815 2.23 11.12 2.3 ;
      RECT 10.935 2.195 11.16 2.29 ;
      RECT 10.815 2.26 11.17 2.285 ;
      RECT 10.895 2.205 11.16 2.29 ;
      RECT 10.975 2.18 11.12 2.305 ;
      RECT 11.055 2.155 11.095 2.315 ;
      RECT 11.015 2.165 11.12 2.305 ;
      RECT 10.855 6 10.935 6.15 ;
      RECT 10.855 6 10.975 6.135 ;
      RECT 10.855 6 11.015 6.12 ;
      RECT 10.855 6 11.055 6.105 ;
      RECT 11.095 5.92 11.12 6.085 ;
      RECT 10.815 6.01 11.12 6.08 ;
      RECT 10.935 5.975 11.16 6.07 ;
      RECT 10.815 6.04 11.17 6.065 ;
      RECT 10.895 5.985 11.16 6.07 ;
      RECT 10.975 5.96 11.12 6.085 ;
      RECT 11.055 5.935 11.095 6.095 ;
      RECT 11.015 5.945 11.12 6.085 ;
      RECT 10.78 2.705 10.82 2.975 ;
      RECT 10.74 2.78 10.86 2.95 ;
      RECT 10.74 2.855 10.9 2.93 ;
      RECT 10.74 2.895 10.91 2.915 ;
      RECT 10.7 2.645 10.74 2.88 ;
      RECT 10.66 2.665 10.78 2.805 ;
      RECT 10.62 2.685 10.78 2.735 ;
      RECT 10.7 2.65 10.78 2.88 ;
      RECT 10.78 6.485 10.82 6.755 ;
      RECT 10.74 6.56 10.86 6.73 ;
      RECT 10.74 6.635 10.9 6.71 ;
      RECT 10.74 6.675 10.91 6.695 ;
      RECT 10.7 6.425 10.74 6.66 ;
      RECT 10.66 6.445 10.78 6.585 ;
      RECT 10.62 6.465 10.78 6.515 ;
      RECT 10.7 6.43 10.78 6.66 ;
      RECT 10.615 1.465 10.655 1.64 ;
      RECT 10.575 1.49 10.655 1.625 ;
      RECT 10.575 1.49 10.695 1.62 ;
      RECT 10.575 1.49 10.735 1.595 ;
      RECT 10.535 1.51 10.775 1.565 ;
      RECT 10.775 1.375 10.815 1.55 ;
      RECT 10.775 1.395 10.855 1.525 ;
      RECT 10.615 1.465 10.89 1.51 ;
      RECT 10.655 1.445 10.855 1.525 ;
      RECT 10.735 1.4 10.775 1.57 ;
      RECT 10.695 1.42 10.855 1.525 ;
      RECT 10.615 5.245 10.655 5.42 ;
      RECT 10.575 5.27 10.655 5.405 ;
      RECT 10.575 5.27 10.695 5.4 ;
      RECT 10.575 5.27 10.735 5.375 ;
      RECT 10.535 5.29 10.775 5.345 ;
      RECT 10.775 5.155 10.815 5.33 ;
      RECT 10.775 5.175 10.855 5.305 ;
      RECT 10.615 5.245 10.89 5.29 ;
      RECT 10.655 5.225 10.855 5.305 ;
      RECT 10.735 5.18 10.775 5.35 ;
      RECT 10.695 5.2 10.855 5.305 ;
      RECT 10.17 1.115 10.19 1.46 ;
      RECT 10.17 1.175 10.23 1.445 ;
      RECT 10.13 1.295 10.27 1.435 ;
      RECT 10.13 1.39 10.29 1.425 ;
      RECT 10.09 1.14 10.19 1.345 ;
      RECT 10.05 1.15 10.19 1.22 ;
      RECT 10.13 1.125 10.19 1.435 ;
      RECT 10.17 4.895 10.19 5.24 ;
      RECT 10.17 4.955 10.23 5.225 ;
      RECT 10.13 5.075 10.27 5.215 ;
      RECT 10.13 5.17 10.29 5.205 ;
      RECT 10.09 4.92 10.19 5.125 ;
      RECT 10.05 4.93 10.19 5 ;
      RECT 10.13 4.905 10.19 5.215 ;
      RECT 10.02 2.92 10.04 3.26 ;
      RECT 10.02 2.98 10.08 3.25 ;
      RECT 9.98 3.1 10.12 3.24 ;
      RECT 9.98 3.195 10.14 3.23 ;
      RECT 9.94 2.945 10.04 3.16 ;
      RECT 9.9 2.955 10.04 3.035 ;
      RECT 9.98 2.93 10.04 3.24 ;
      RECT 10.02 6.7 10.04 7.04 ;
      RECT 10.02 6.76 10.08 7.03 ;
      RECT 9.98 6.88 10.12 7.02 ;
      RECT 9.98 6.975 10.14 7.01 ;
      RECT 9.94 6.725 10.04 6.94 ;
      RECT 9.9 6.735 10.04 6.815 ;
      RECT 9.98 6.71 10.04 7.02 ;
      RECT 9.375 2.82 9.415 2.99 ;
      RECT 9.335 2.84 9.415 2.975 ;
      RECT 9.335 2.84 9.455 2.97 ;
      RECT 9.335 2.84 9.535 2.93 ;
      RECT 9.295 2.865 9.535 2.915 ;
      RECT 9.295 2.865 9.575 2.905 ;
      RECT 9.575 2.72 9.585 2.895 ;
      RECT 9.495 2.755 9.625 2.88 ;
      RECT 9.375 2.82 9.655 2.86 ;
      RECT 9.415 2.8 9.625 2.88 ;
      RECT 9.455 2.78 9.495 2.95 ;
      RECT 9.535 2.735 9.585 2.895 ;
      RECT 9.375 6.6 9.415 6.77 ;
      RECT 9.335 6.62 9.415 6.755 ;
      RECT 9.335 6.62 9.455 6.75 ;
      RECT 9.335 6.62 9.535 6.71 ;
      RECT 9.295 6.645 9.535 6.695 ;
      RECT 9.295 6.645 9.575 6.685 ;
      RECT 9.575 6.5 9.585 6.675 ;
      RECT 9.495 6.535 9.625 6.66 ;
      RECT 9.375 6.6 9.655 6.64 ;
      RECT 9.415 6.58 9.625 6.66 ;
      RECT 9.455 6.56 9.495 6.73 ;
      RECT 9.535 6.515 9.585 6.675 ;
      RECT 9.42 1.48 9.46 1.745 ;
      RECT 9.38 1.555 9.5 1.72 ;
      RECT 9.38 1.625 9.54 1.7 ;
      RECT 9.38 1.665 9.55 1.685 ;
      RECT 9.34 1.415 9.38 1.65 ;
      RECT 9.3 1.44 9.42 1.58 ;
      RECT 9.26 1.46 9.42 1.51 ;
      RECT 9.34 1.425 9.42 1.65 ;
      RECT 9.42 5.26 9.46 5.525 ;
      RECT 9.38 5.335 9.5 5.5 ;
      RECT 9.38 5.405 9.54 5.48 ;
      RECT 9.38 5.445 9.55 5.465 ;
      RECT 9.34 5.195 9.38 5.43 ;
      RECT 9.3 5.22 9.42 5.36 ;
      RECT 9.26 5.24 9.42 5.29 ;
      RECT 9.34 5.205 9.42 5.43 ;
      RECT 9.045 2.08 9.085 2.23 ;
      RECT 9.045 2.08 9.125 2.225 ;
      RECT 9.045 2.08 9.165 2.21 ;
      RECT 9.045 2.08 9.205 2.2 ;
      RECT 9.285 2 9.31 2.17 ;
      RECT 9.005 2.09 9.31 2.165 ;
      RECT 9.125 2.06 9.35 2.155 ;
      RECT 9.005 2.135 9.355 2.145 ;
      RECT 9.085 2.065 9.35 2.155 ;
      RECT 9.125 2.055 9.31 2.17 ;
      RECT 9.245 2.015 9.285 2.175 ;
      RECT 9.165 2.04 9.31 2.17 ;
      RECT 9.205 2.025 9.245 2.185 ;
      RECT 9.045 5.86 9.085 6.01 ;
      RECT 9.045 5.86 9.125 6.005 ;
      RECT 9.045 5.86 9.165 5.99 ;
      RECT 9.045 5.86 9.205 5.98 ;
      RECT 9.285 5.78 9.31 5.95 ;
      RECT 9.005 5.87 9.31 5.945 ;
      RECT 9.125 5.84 9.35 5.935 ;
      RECT 9.005 5.915 9.355 5.925 ;
      RECT 9.085 5.845 9.35 5.935 ;
      RECT 9.125 5.835 9.31 5.95 ;
      RECT 9.245 5.795 9.285 5.955 ;
      RECT 9.165 5.82 9.31 5.95 ;
      RECT 9.205 5.805 9.245 5.965 ;
      RECT 7.075 2.22 7.155 2.37 ;
      RECT 7.075 2.22 7.195 2.355 ;
      RECT 7.075 2.22 7.235 2.34 ;
      RECT 7.075 2.22 7.275 2.325 ;
      RECT 7.315 2.14 7.34 2.305 ;
      RECT 7.035 2.23 7.34 2.3 ;
      RECT 7.155 2.195 7.38 2.29 ;
      RECT 7.035 2.26 7.39 2.285 ;
      RECT 7.115 2.205 7.38 2.29 ;
      RECT 7.195 2.18 7.34 2.305 ;
      RECT 7.275 2.155 7.315 2.315 ;
      RECT 7.235 2.165 7.34 2.305 ;
      RECT 7.075 6 7.155 6.15 ;
      RECT 7.075 6 7.195 6.135 ;
      RECT 7.075 6 7.235 6.12 ;
      RECT 7.075 6 7.275 6.105 ;
      RECT 7.315 5.92 7.34 6.085 ;
      RECT 7.035 6.01 7.34 6.08 ;
      RECT 7.155 5.975 7.38 6.07 ;
      RECT 7.035 6.04 7.39 6.065 ;
      RECT 7.115 5.985 7.38 6.07 ;
      RECT 7.195 5.96 7.34 6.085 ;
      RECT 7.275 5.935 7.315 6.095 ;
      RECT 7.235 5.945 7.34 6.085 ;
      RECT 7 2.705 7.04 2.975 ;
      RECT 6.96 2.78 7.08 2.95 ;
      RECT 6.96 2.855 7.12 2.93 ;
      RECT 6.96 2.895 7.13 2.915 ;
      RECT 6.92 2.645 6.96 2.88 ;
      RECT 6.88 2.665 7 2.805 ;
      RECT 6.84 2.685 7 2.735 ;
      RECT 6.92 2.65 7 2.88 ;
      RECT 7 6.485 7.04 6.755 ;
      RECT 6.96 6.56 7.08 6.73 ;
      RECT 6.96 6.635 7.12 6.71 ;
      RECT 6.96 6.675 7.13 6.695 ;
      RECT 6.92 6.425 6.96 6.66 ;
      RECT 6.88 6.445 7 6.585 ;
      RECT 6.84 6.465 7 6.515 ;
      RECT 6.92 6.43 7 6.66 ;
      RECT 6.835 1.465 6.875 1.64 ;
      RECT 6.795 1.49 6.875 1.625 ;
      RECT 6.795 1.49 6.915 1.62 ;
      RECT 6.795 1.49 6.955 1.595 ;
      RECT 6.755 1.51 6.995 1.565 ;
      RECT 6.995 1.375 7.035 1.55 ;
      RECT 6.995 1.395 7.075 1.525 ;
      RECT 6.835 1.465 7.11 1.51 ;
      RECT 6.875 1.445 7.075 1.525 ;
      RECT 6.955 1.4 6.995 1.57 ;
      RECT 6.915 1.42 7.075 1.525 ;
      RECT 6.835 5.245 6.875 5.42 ;
      RECT 6.795 5.27 6.875 5.405 ;
      RECT 6.795 5.27 6.915 5.4 ;
      RECT 6.795 5.27 6.955 5.375 ;
      RECT 6.755 5.29 6.995 5.345 ;
      RECT 6.995 5.155 7.035 5.33 ;
      RECT 6.995 5.175 7.075 5.305 ;
      RECT 6.835 5.245 7.11 5.29 ;
      RECT 6.875 5.225 7.075 5.305 ;
      RECT 6.955 5.18 6.995 5.35 ;
      RECT 6.915 5.2 7.075 5.305 ;
      RECT 6.39 1.115 6.41 1.46 ;
      RECT 6.39 1.175 6.45 1.445 ;
      RECT 6.35 1.295 6.49 1.435 ;
      RECT 6.35 1.39 6.51 1.425 ;
      RECT 6.31 1.14 6.41 1.345 ;
      RECT 6.27 1.15 6.41 1.22 ;
      RECT 6.35 1.125 6.41 1.435 ;
      RECT 6.39 4.895 6.41 5.24 ;
      RECT 6.39 4.955 6.45 5.225 ;
      RECT 6.35 5.075 6.49 5.215 ;
      RECT 6.35 5.17 6.51 5.205 ;
      RECT 6.31 4.92 6.41 5.125 ;
      RECT 6.27 4.93 6.41 5 ;
      RECT 6.35 4.905 6.41 5.215 ;
      RECT 6.24 2.92 6.26 3.26 ;
      RECT 6.24 2.98 6.3 3.25 ;
      RECT 6.2 3.1 6.34 3.24 ;
      RECT 6.2 3.195 6.36 3.23 ;
      RECT 6.16 2.945 6.26 3.16 ;
      RECT 6.12 2.955 6.26 3.035 ;
      RECT 6.2 2.93 6.26 3.24 ;
      RECT 6.24 6.7 6.26 7.04 ;
      RECT 6.24 6.76 6.3 7.03 ;
      RECT 6.2 6.88 6.34 7.02 ;
      RECT 6.2 6.975 6.36 7.01 ;
      RECT 6.16 6.725 6.26 6.94 ;
      RECT 6.12 6.735 6.26 6.815 ;
      RECT 6.2 6.71 6.26 7.02 ;
      RECT 5.595 2.82 5.635 2.99 ;
      RECT 5.555 2.84 5.635 2.975 ;
      RECT 5.555 2.84 5.675 2.97 ;
      RECT 5.555 2.84 5.755 2.93 ;
      RECT 5.515 2.865 5.755 2.915 ;
      RECT 5.515 2.865 5.795 2.905 ;
      RECT 5.795 2.72 5.805 2.895 ;
      RECT 5.715 2.755 5.845 2.88 ;
      RECT 5.595 2.82 5.875 2.86 ;
      RECT 5.635 2.8 5.845 2.88 ;
      RECT 5.675 2.78 5.715 2.95 ;
      RECT 5.755 2.735 5.805 2.895 ;
      RECT 5.595 6.6 5.635 6.77 ;
      RECT 5.555 6.62 5.635 6.755 ;
      RECT 5.555 6.62 5.675 6.75 ;
      RECT 5.555 6.62 5.755 6.71 ;
      RECT 5.515 6.645 5.755 6.695 ;
      RECT 5.515 6.645 5.795 6.685 ;
      RECT 5.795 6.5 5.805 6.675 ;
      RECT 5.715 6.535 5.845 6.66 ;
      RECT 5.595 6.6 5.875 6.64 ;
      RECT 5.635 6.58 5.845 6.66 ;
      RECT 5.675 6.56 5.715 6.73 ;
      RECT 5.755 6.515 5.805 6.675 ;
      RECT 5.64 1.48 5.68 1.745 ;
      RECT 5.6 1.555 5.72 1.72 ;
      RECT 5.6 1.625 5.76 1.7 ;
      RECT 5.6 1.665 5.77 1.685 ;
      RECT 5.56 1.415 5.6 1.65 ;
      RECT 5.52 1.44 5.64 1.58 ;
      RECT 5.48 1.46 5.64 1.51 ;
      RECT 5.56 1.425 5.64 1.65 ;
      RECT 5.64 5.26 5.68 5.525 ;
      RECT 5.6 5.335 5.72 5.5 ;
      RECT 5.6 5.405 5.76 5.48 ;
      RECT 5.6 5.445 5.77 5.465 ;
      RECT 5.56 5.195 5.6 5.43 ;
      RECT 5.52 5.22 5.64 5.36 ;
      RECT 5.48 5.24 5.64 5.29 ;
      RECT 5.56 5.205 5.64 5.43 ;
      RECT 5.265 2.08 5.305 2.23 ;
      RECT 5.265 2.08 5.345 2.225 ;
      RECT 5.265 2.08 5.385 2.21 ;
      RECT 5.265 2.08 5.425 2.2 ;
      RECT 5.505 2 5.53 2.17 ;
      RECT 5.225 2.09 5.53 2.165 ;
      RECT 5.345 2.06 5.57 2.155 ;
      RECT 5.225 2.135 5.575 2.145 ;
      RECT 5.305 2.065 5.57 2.155 ;
      RECT 5.345 2.055 5.53 2.17 ;
      RECT 5.465 2.015 5.505 2.175 ;
      RECT 5.385 2.04 5.53 2.17 ;
      RECT 5.425 2.025 5.465 2.185 ;
      RECT 5.265 5.86 5.305 6.01 ;
      RECT 5.265 5.86 5.345 6.005 ;
      RECT 5.265 5.86 5.385 5.99 ;
      RECT 5.265 5.86 5.425 5.98 ;
      RECT 5.505 5.78 5.53 5.95 ;
      RECT 5.225 5.87 5.53 5.945 ;
      RECT 5.345 5.84 5.57 5.935 ;
      RECT 5.225 5.915 5.575 5.925 ;
      RECT 5.305 5.845 5.57 5.935 ;
      RECT 5.345 5.835 5.53 5.95 ;
      RECT 5.465 5.795 5.505 5.955 ;
      RECT 5.385 5.82 5.53 5.95 ;
      RECT 5.425 5.805 5.465 5.965 ;
      RECT 3.295 2.22 3.375 2.37 ;
      RECT 3.295 2.22 3.415 2.355 ;
      RECT 3.295 2.22 3.455 2.34 ;
      RECT 3.295 2.22 3.495 2.325 ;
      RECT 3.535 2.14 3.56 2.305 ;
      RECT 3.255 2.23 3.56 2.3 ;
      RECT 3.375 2.195 3.6 2.29 ;
      RECT 3.255 2.26 3.61 2.285 ;
      RECT 3.335 2.205 3.6 2.29 ;
      RECT 3.415 2.18 3.56 2.305 ;
      RECT 3.495 2.155 3.535 2.315 ;
      RECT 3.455 2.165 3.56 2.305 ;
      RECT 3.295 6 3.375 6.15 ;
      RECT 3.295 6 3.415 6.135 ;
      RECT 3.295 6 3.455 6.12 ;
      RECT 3.295 6 3.495 6.105 ;
      RECT 3.535 5.92 3.56 6.085 ;
      RECT 3.255 6.01 3.56 6.08 ;
      RECT 3.375 5.975 3.6 6.07 ;
      RECT 3.255 6.04 3.61 6.065 ;
      RECT 3.335 5.985 3.6 6.07 ;
      RECT 3.415 5.96 3.56 6.085 ;
      RECT 3.495 5.935 3.535 6.095 ;
      RECT 3.455 5.945 3.56 6.085 ;
      RECT 3.22 2.705 3.26 2.975 ;
      RECT 3.18 2.78 3.3 2.95 ;
      RECT 3.18 2.855 3.34 2.93 ;
      RECT 3.18 2.895 3.35 2.915 ;
      RECT 3.14 2.645 3.18 2.88 ;
      RECT 3.1 2.665 3.22 2.805 ;
      RECT 3.06 2.685 3.22 2.735 ;
      RECT 3.14 2.65 3.22 2.88 ;
      RECT 3.22 6.485 3.26 6.755 ;
      RECT 3.18 6.56 3.3 6.73 ;
      RECT 3.18 6.635 3.34 6.71 ;
      RECT 3.18 6.675 3.35 6.695 ;
      RECT 3.14 6.425 3.18 6.66 ;
      RECT 3.1 6.445 3.22 6.585 ;
      RECT 3.06 6.465 3.22 6.515 ;
      RECT 3.14 6.43 3.22 6.66 ;
      RECT 3.055 1.465 3.095 1.64 ;
      RECT 3.015 1.49 3.095 1.625 ;
      RECT 3.015 1.49 3.135 1.62 ;
      RECT 3.015 1.49 3.175 1.595 ;
      RECT 2.975 1.51 3.215 1.565 ;
      RECT 3.215 1.375 3.255 1.55 ;
      RECT 3.215 1.395 3.295 1.525 ;
      RECT 3.055 1.465 3.33 1.51 ;
      RECT 3.095 1.445 3.295 1.525 ;
      RECT 3.175 1.4 3.215 1.57 ;
      RECT 3.135 1.42 3.295 1.525 ;
      RECT 3.055 5.245 3.095 5.42 ;
      RECT 3.015 5.27 3.095 5.405 ;
      RECT 3.015 5.27 3.135 5.4 ;
      RECT 3.015 5.27 3.175 5.375 ;
      RECT 2.975 5.29 3.215 5.345 ;
      RECT 3.215 5.155 3.255 5.33 ;
      RECT 3.215 5.175 3.295 5.305 ;
      RECT 3.055 5.245 3.33 5.29 ;
      RECT 3.095 5.225 3.295 5.305 ;
      RECT 3.175 5.18 3.215 5.35 ;
      RECT 3.135 5.2 3.295 5.305 ;
      RECT 2.61 1.115 2.63 1.46 ;
      RECT 2.61 1.175 2.67 1.445 ;
      RECT 2.57 1.295 2.71 1.435 ;
      RECT 2.57 1.39 2.73 1.425 ;
      RECT 2.53 1.14 2.63 1.345 ;
      RECT 2.49 1.15 2.63 1.22 ;
      RECT 2.57 1.125 2.63 1.435 ;
      RECT 2.61 4.895 2.63 5.24 ;
      RECT 2.61 4.955 2.67 5.225 ;
      RECT 2.57 5.075 2.71 5.215 ;
      RECT 2.57 5.17 2.73 5.205 ;
      RECT 2.53 4.92 2.63 5.125 ;
      RECT 2.49 4.93 2.63 5 ;
      RECT 2.57 4.905 2.63 5.215 ;
      RECT 2.46 2.92 2.48 3.26 ;
      RECT 2.46 2.98 2.52 3.25 ;
      RECT 2.42 3.1 2.56 3.24 ;
      RECT 2.42 3.195 2.58 3.23 ;
      RECT 2.38 2.945 2.48 3.16 ;
      RECT 2.34 2.955 2.48 3.035 ;
      RECT 2.42 2.93 2.48 3.24 ;
      RECT 2.46 6.7 2.48 7.04 ;
      RECT 2.46 6.76 2.52 7.03 ;
      RECT 2.42 6.88 2.56 7.02 ;
      RECT 2.42 6.975 2.58 7.01 ;
      RECT 2.38 6.725 2.48 6.94 ;
      RECT 2.34 6.735 2.48 6.815 ;
      RECT 2.42 6.71 2.48 7.02 ;
      RECT 1.815 2.82 1.855 2.99 ;
      RECT 1.775 2.84 1.855 2.975 ;
      RECT 1.775 2.84 1.895 2.97 ;
      RECT 1.775 2.84 1.975 2.93 ;
      RECT 1.735 2.865 1.975 2.915 ;
      RECT 1.735 2.865 2.015 2.905 ;
      RECT 2.015 2.72 2.025 2.895 ;
      RECT 1.935 2.755 2.065 2.88 ;
      RECT 1.815 2.82 2.095 2.86 ;
      RECT 1.855 2.8 2.065 2.88 ;
      RECT 1.895 2.78 1.935 2.95 ;
      RECT 1.975 2.735 2.025 2.895 ;
      RECT 1.815 6.6 1.855 6.77 ;
      RECT 1.775 6.62 1.855 6.755 ;
      RECT 1.775 6.62 1.895 6.75 ;
      RECT 1.775 6.62 1.975 6.71 ;
      RECT 1.735 6.645 1.975 6.695 ;
      RECT 1.735 6.645 2.015 6.685 ;
      RECT 2.015 6.5 2.025 6.675 ;
      RECT 1.935 6.535 2.065 6.66 ;
      RECT 1.815 6.6 2.095 6.64 ;
      RECT 1.855 6.58 2.065 6.66 ;
      RECT 1.895 6.56 1.935 6.73 ;
      RECT 1.975 6.515 2.025 6.675 ;
      RECT 1.86 1.48 1.9 1.745 ;
      RECT 1.82 1.555 1.94 1.72 ;
      RECT 1.82 1.625 1.98 1.7 ;
      RECT 1.82 1.665 1.99 1.685 ;
      RECT 1.78 1.415 1.82 1.65 ;
      RECT 1.74 1.44 1.86 1.58 ;
      RECT 1.7 1.46 1.86 1.51 ;
      RECT 1.78 1.425 1.86 1.65 ;
      RECT 1.86 5.26 1.9 5.525 ;
      RECT 1.82 5.335 1.94 5.5 ;
      RECT 1.82 5.405 1.98 5.48 ;
      RECT 1.82 5.445 1.99 5.465 ;
      RECT 1.78 5.195 1.82 5.43 ;
      RECT 1.74 5.22 1.86 5.36 ;
      RECT 1.7 5.24 1.86 5.29 ;
      RECT 1.78 5.205 1.86 5.43 ;
      RECT 1.485 2.08 1.525 2.23 ;
      RECT 1.485 2.08 1.565 2.225 ;
      RECT 1.485 2.08 1.605 2.21 ;
      RECT 1.485 2.08 1.645 2.2 ;
      RECT 1.725 2 1.75 2.17 ;
      RECT 1.445 2.09 1.75 2.165 ;
      RECT 1.565 2.06 1.79 2.155 ;
      RECT 1.445 2.135 1.795 2.145 ;
      RECT 1.525 2.065 1.79 2.155 ;
      RECT 1.565 2.055 1.75 2.17 ;
      RECT 1.685 2.015 1.725 2.175 ;
      RECT 1.605 2.04 1.75 2.17 ;
      RECT 1.645 2.025 1.685 2.185 ;
      RECT 1.485 5.86 1.525 6.01 ;
      RECT 1.485 5.86 1.565 6.005 ;
      RECT 1.485 5.86 1.605 5.99 ;
      RECT 1.485 5.86 1.645 5.98 ;
      RECT 1.725 5.78 1.75 5.95 ;
      RECT 1.445 5.87 1.75 5.945 ;
      RECT 1.565 5.84 1.79 5.935 ;
      RECT 1.445 5.915 1.795 5.925 ;
      RECT 1.525 5.845 1.79 5.935 ;
      RECT 1.565 5.835 1.75 5.95 ;
      RECT 1.685 5.795 1.725 5.955 ;
      RECT 1.605 5.82 1.75 5.95 ;
      RECT 1.645 5.805 1.685 5.965 ;
    LAYER NEMBODY ;
      RECT 19.24 7.56 19.84 8.16 ;
      RECT 15.46 7.56 16.06 8.16 ;
      RECT 15.86 4.58 16.06 8.16 ;
      RECT 11.68 7.56 12.28 8.16 ;
      RECT 12.08 4.58 12.28 8.16 ;
      RECT 7.9 7.56 8.5 8.16 ;
      RECT 8.3 4.58 8.5 8.16 ;
      RECT 4.12 7.56 4.72 8.16 ;
      RECT 4.52 4.58 4.72 8.16 ;
      RECT 0.34 7.56 0.94 8.16 ;
      RECT 0.74 4.58 0.94 8.16 ;
      RECT 16.26 7.56 19.84 7.76 ;
      RECT 12.48 7.56 16.06 7.76 ;
      RECT 8.7 7.56 12.28 7.76 ;
      RECT 4.92 7.56 8.5 7.76 ;
      RECT 1.14 7.56 4.72 7.76 ;
      RECT 16.26 4.58 16.46 7.76 ;
      RECT 12.48 4.58 12.68 7.76 ;
      RECT 8.7 4.58 8.9 7.76 ;
      RECT 4.92 4.58 5.12 7.76 ;
      RECT 1.14 4.58 1.34 7.76 ;
      RECT 16.26 7.16 19.44 7.36 ;
      RECT 19.24 3.78 19.44 7.36 ;
      RECT 12.48 7.16 15.66 7.36 ;
      RECT 15.46 3.78 15.66 7.36 ;
      RECT 8.7 7.16 11.88 7.36 ;
      RECT 11.68 3.78 11.88 7.36 ;
      RECT 4.92 7.16 8.1 7.36 ;
      RECT 7.9 3.78 8.1 7.36 ;
      RECT 1.14 7.16 4.32 7.36 ;
      RECT 4.12 3.78 4.32 7.36 ;
      RECT 16.26 4.58 19.04 7.36 ;
      RECT 18.84 4.18 19.04 7.36 ;
      RECT 12.48 4.58 15.26 7.36 ;
      RECT 15.06 4.18 15.26 7.36 ;
      RECT 8.7 4.58 11.48 7.36 ;
      RECT 11.28 4.18 11.48 7.36 ;
      RECT 4.92 4.58 7.7 7.36 ;
      RECT 7.5 4.18 7.7 7.36 ;
      RECT 1.14 4.58 3.92 7.36 ;
      RECT 3.72 4.18 3.92 7.36 ;
      RECT 15.86 4.58 19.04 4.78 ;
      RECT 12.08 4.58 15.26 4.78 ;
      RECT 8.3 4.58 11.48 4.78 ;
      RECT 4.52 4.58 7.7 4.78 ;
      RECT 0.74 4.58 3.92 4.78 ;
      RECT 19.24 3.78 19.84 4.38 ;
      RECT 15.46 4.18 19.04 4.38 ;
      RECT 11.68 4.18 15.26 4.38 ;
      RECT 7.9 4.18 11.48 4.38 ;
      RECT 4.12 4.18 7.7 4.38 ;
      RECT 0.34 4.18 3.92 4.38 ;
      RECT 15.46 3.78 16.06 4.38 ;
      RECT 15.86 0.8 16.06 4.38 ;
      RECT 11.68 3.78 12.28 4.38 ;
      RECT 12.08 0.8 12.28 4.38 ;
      RECT 7.9 3.78 8.5 4.38 ;
      RECT 8.3 0.8 8.5 4.38 ;
      RECT 4.12 3.78 4.72 4.38 ;
      RECT 4.52 0.8 4.72 4.38 ;
      RECT 0.34 3.78 0.94 4.38 ;
      RECT 0.74 0.8 0.94 4.38 ;
      RECT 16.26 3.78 19.84 3.98 ;
      RECT 12.48 3.78 16.06 3.98 ;
      RECT 8.7 3.78 12.28 3.98 ;
      RECT 4.92 3.78 8.5 3.98 ;
      RECT 1.14 3.78 4.72 3.98 ;
      RECT 16.26 0.8 16.46 3.98 ;
      RECT 12.48 0.8 12.68 3.98 ;
      RECT 8.7 0.8 8.9 3.98 ;
      RECT 4.92 0.8 5.12 3.98 ;
      RECT 1.14 0.8 1.34 3.98 ;
      RECT 16.26 3.38 19.44 3.58 ;
      RECT 19.24 0 19.44 3.58 ;
      RECT 12.48 3.38 15.66 3.58 ;
      RECT 15.46 0 15.66 3.58 ;
      RECT 8.7 3.38 11.88 3.58 ;
      RECT 11.68 0 11.88 3.58 ;
      RECT 4.92 3.38 8.1 3.58 ;
      RECT 7.9 0 8.1 3.58 ;
      RECT 1.14 3.38 4.32 3.58 ;
      RECT 4.12 0 4.32 3.58 ;
      RECT 16.26 0.8 19.04 3.58 ;
      RECT 18.84 0.4 19.04 3.58 ;
      RECT 12.48 0.8 15.26 3.58 ;
      RECT 15.06 0.4 15.26 3.58 ;
      RECT 8.7 0.8 11.48 3.58 ;
      RECT 11.28 0.4 11.48 3.58 ;
      RECT 4.92 0.8 7.7 3.58 ;
      RECT 7.5 0.4 7.7 3.58 ;
      RECT 1.14 0.8 3.92 3.58 ;
      RECT 3.72 0.4 3.92 3.58 ;
      RECT 15.86 0.8 19.04 1 ;
      RECT 12.08 0.8 15.26 1 ;
      RECT 8.3 0.8 11.48 1 ;
      RECT 4.52 0.8 7.7 1 ;
      RECT 0.74 0.8 3.92 1 ;
      RECT 19.24 0 19.84 0.6 ;
      RECT 15.46 0.4 19.04 0.6 ;
      RECT 11.68 0.4 15.26 0.6 ;
      RECT 7.9 0.4 11.48 0.6 ;
      RECT 4.12 0.4 7.7 0.6 ;
      RECT 0.34 0.4 3.92 0.6 ;
      RECT 15.46 0 16.06 0.6 ;
      RECT 11.68 0 12.28 0.6 ;
      RECT 7.9 0 8.5 0.6 ;
      RECT 4.12 0 4.72 0.6 ;
      RECT 0.34 0 0.94 0.6 ;
  END
END nem_ohmux_invd2_10i_8b

END LIBRARY
