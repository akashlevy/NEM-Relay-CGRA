###############################################################################
#TSMC Library/IP Product
#Filename: tphn40lpgv2od3_sl_9lm.lef
#Technology: N40
#Product Type: Standard I/O
#Product Name: tphn40lpgv2od3_sl
#Version: 210a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.005 BY 120.000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 120.000 BY 120.000 ;
END corner

MACRO PCLAMP1ANA_G
    CLASS BLOCK ;
    FOREIGN PCLAMP1ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 76.000 BY 53.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        END
    END VSSESD
    PIN VDDESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER VIA2 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 76.000 53.000 ;
    END
END PCLAMP1ANA_G

MACRO PCLAMP2ANA_G
    CLASS BLOCK ;
    FOREIGN PCLAMP2ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 76.000 BY 53.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        END
    END VSSESD
    PIN VDDESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER VIA2 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 76.000 53.000 ;
    END
END PCLAMP2ANA_G

MACRO PCLAMPAC_G
    CLASS BLOCK ;
    FOREIGN PCLAMPAC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 76.000 BY 53.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        END
    END VSSESD
    PIN VDDESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER VIA2 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 76.000 53.000 ;
    END
END PCLAMPAC_G

MACRO PCLAMPA_G
    CLASS BLOCK ;
    FOREIGN PCLAMPA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 76.000 BY 53.000 ;
    SYMMETRY X Y R90 ;
    PIN VSSESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M3 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        END
    END VSSESD
    PIN VDDESD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        END
    END VDDESD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 76.000 53.000 ;
        LAYER VIA2 ;
        RECT  71.385 0.000 74.385 53.000 ;
        RECT  66.685 0.000 70.385 53.000 ;
        RECT  61.985 0.000 65.685 53.000 ;
        RECT  57.285 0.000 60.985 53.000 ;
        RECT  52.585 0.000 56.285 53.000 ;
        RECT  47.885 0.000 51.585 53.000 ;
        RECT  44.380 0.000 46.885 53.000 ;
        RECT  37.650 0.000 41.375 53.000 ;
        RECT  30.875 0.000 35.375 53.000 ;
        RECT  24.875 0.000 29.375 53.000 ;
        RECT  19.625 0.000 23.375 53.000 ;
        RECT  13.870 0.000 17.870 53.000 ;
        RECT  7.870 0.000 11.870 53.000 ;
        RECT  1.615 0.000 5.615 53.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 76.000 53.000 ;
    END
END PCLAMPA_G

MACRO PCORNERA_G
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNERA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 120.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE corner ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M6 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M5 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M4 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M3 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  77.530 7.250 120.000 11.750 ;
                POLYGON  36.750 82.120 82.120 36.750 120.000 36.750 120.000 39.290 83.275 39.290
                 39.290 83.275 39.290 120.000 36.750 120.000 ;
                POLYGON  31.250 79.720 79.720 31.250 120.000 31.250 120.000 35.750 81.565 35.750
                 35.750 81.565 35.750 120.000 31.250 120.000 ;
                POLYGON  25.250 76.990 25.575 76.665 25.575 76.585 25.655 76.585 76.585 25.655
                 76.585 25.575 76.665 25.575 76.990 25.250 120.000 25.250 120.000 29.750
                 78.835 29.750 29.750 78.835 29.750 120.000 25.250 120.000 ;
                POLYGON  19.250 74.260 74.260 19.250 120.000 19.250 120.000 23.750 76.105 23.750
                 23.750 76.105 23.750 120.000 19.250 120.000 ;
                POLYGON  13.250 71.530 71.530 13.250 120.000 13.250 120.000 17.750 73.375 17.750
                 17.750 73.375 17.750 120.000 13.250 120.000 ;
        RECT  7.250 77.530 11.750 120.000 ;
                POLYGON  1.250 74.800 74.800 1.250 120.000 1.250 120.000 5.750 76.645 5.750
                 5.750 76.645 5.750 120.000 1.250 120.000 ;
        LAYER M6 ;
        RECT  77.530 7.250 120.000 11.750 ;
                POLYGON  36.750 82.120 82.120 36.750 120.000 36.750 120.000 39.290 83.275 39.290
                 39.290 83.275 39.290 120.000 36.750 120.000 ;
                POLYGON  31.250 79.720 79.720 31.250 120.000 31.250 120.000 35.750 81.565 35.750
                 35.750 81.565 35.750 120.000 31.250 120.000 ;
                POLYGON  25.250 76.990 25.575 76.665 25.575 76.585 25.655 76.585 76.585 25.655
                 76.585 25.575 76.665 25.575 76.990 25.250 120.000 25.250 120.000 29.750
                 78.835 29.750 29.750 78.835 29.750 120.000 25.250 120.000 ;
                POLYGON  19.250 74.260 74.260 19.250 120.000 19.250 120.000 23.750 76.105 23.750
                 23.750 76.105 23.750 120.000 19.250 120.000 ;
                POLYGON  13.250 71.530 71.530 13.250 120.000 13.250 120.000 17.750 73.375 17.750
                 17.750 73.375 17.750 120.000 13.250 120.000 ;
        RECT  7.250 77.530 11.750 120.000 ;
                POLYGON  1.250 74.800 74.800 1.250 120.000 1.250 120.000 5.750 76.645 5.750
                 5.750 76.645 5.750 120.000 1.250 120.000 ;
        LAYER M5 ;
        RECT  77.530 7.250 120.000 11.750 ;
                POLYGON  36.750 82.120 82.120 36.750 120.000 36.750 120.000 39.290 83.275 39.290
                 39.290 83.275 39.290 120.000 36.750 120.000 ;
                POLYGON  31.250 79.720 79.720 31.250 120.000 31.250 120.000 35.750 81.565 35.750
                 35.750 81.565 35.750 120.000 31.250 120.000 ;
                POLYGON  25.250 76.990 25.575 76.665 25.575 76.585 25.655 76.585 76.585 25.655
                 76.585 25.575 76.665 25.575 76.990 25.250 120.000 25.250 120.000 29.750
                 78.835 29.750 29.750 78.835 29.750 120.000 25.250 120.000 ;
                POLYGON  19.250 74.260 74.260 19.250 120.000 19.250 120.000 23.750 76.105 23.750
                 23.750 76.105 23.750 120.000 19.250 120.000 ;
                POLYGON  13.250 71.530 71.530 13.250 120.000 13.250 120.000 17.750 73.375 17.750
                 17.750 73.375 17.750 120.000 13.250 120.000 ;
        RECT  7.250 77.530 11.750 120.000 ;
                POLYGON  1.250 74.800 74.800 1.250 120.000 1.250 120.000 5.750 76.645 5.750
                 5.750 76.645 5.750 120.000 1.250 120.000 ;
        LAYER M4 ;
        RECT  77.530 7.250 120.000 11.750 ;
                POLYGON  36.750 82.120 82.120 36.750 120.000 36.750 120.000 39.290 83.275 39.290
                 39.290 83.275 39.290 120.000 36.750 120.000 ;
                POLYGON  31.250 79.720 79.720 31.250 120.000 31.250 120.000 35.750 81.565 35.750
                 35.750 81.565 35.750 120.000 31.250 120.000 ;
                POLYGON  25.250 76.990 25.575 76.665 25.575 76.585 25.655 76.585 76.585 25.655
                 76.585 25.575 76.665 25.575 76.990 25.250 120.000 25.250 120.000 29.750
                 78.835 29.750 29.750 78.835 29.750 120.000 25.250 120.000 ;
                POLYGON  19.250 74.260 74.260 19.250 120.000 19.250 120.000 23.750 76.105 23.750
                 23.750 76.105 23.750 120.000 19.250 120.000 ;
                POLYGON  13.250 71.530 71.530 13.250 120.000 13.250 120.000 17.750 73.375 17.750
                 17.750 73.375 17.750 120.000 13.250 120.000 ;
        RECT  7.250 77.530 11.750 120.000 ;
                POLYGON  1.250 74.800 74.800 1.250 120.000 1.250 120.000 5.750 76.645 5.750
                 5.750 76.645 5.750 120.000 1.250 120.000 ;
        LAYER M3 ;
        RECT  77.530 7.250 120.000 11.750 ;
                POLYGON  36.750 82.120 82.120 36.750 120.000 36.750 120.000 39.290 83.275 39.290
                 39.290 83.275 39.290 120.000 36.750 120.000 ;
                POLYGON  31.250 79.720 79.720 31.250 120.000 31.250 120.000 35.750 81.565 35.750
                 35.750 81.565 35.750 120.000 31.250 120.000 ;
                POLYGON  25.250 76.990 25.575 76.665 25.575 76.585 25.655 76.585 76.585 25.655
                 76.585 25.575 76.665 25.575 76.990 25.250 120.000 25.250 120.000 29.750
                 78.835 29.750 29.750 78.835 29.750 120.000 25.250 120.000 ;
                POLYGON  19.250 74.260 74.260 19.250 120.000 19.250 120.000 23.750 76.105 23.750
                 23.750 76.105 23.750 120.000 19.250 120.000 ;
                POLYGON  13.250 71.530 71.530 13.250 120.000 13.250 120.000 17.750 73.375 17.750
                 17.750 73.375 17.750 120.000 13.250 120.000 ;
        RECT  7.250 77.530 11.750 120.000 ;
                POLYGON  1.250 74.800 74.800 1.250 120.000 1.250 120.000 5.750 76.645 5.750
                 5.750 76.645 5.750 120.000 1.250 120.000 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M6 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M5 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M4 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M3 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA1 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 120.000 120.000 ;
    END
END PCORNERA_G

MACRO PCORNER_G
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNER_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 120.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE corner ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  1.250 115.500 5.750 115.500 5.750 68.515 68.515 5.750 115.500 5.750
                 115.500 1.250 120.000 1.250 120.000 4.750 118.000 4.750 118.000 5.750
                 120.000 5.750 120.000 9.250 118.000 9.250 118.000 10.250 120.000 10.250
                 120.000 13.750 118.000 13.750 118.000 14.750 120.000 14.750
                 120.000 18.250 118.000 18.250 118.000 19.250 120.000 19.250
                 120.000 22.750 118.000 22.750 118.000 23.750 120.000 23.750
                 120.000 27.250 118.000 27.250 118.000 28.250 120.000 28.250
                 120.000 31.750 118.000 31.750 118.000 33.080 120.000 33.080
                 120.000 37.580 82.500 37.580 37.580 82.500 37.580 120.000 33.080 120.000
                 33.080 80.650 80.650 33.080 115.500 33.080 115.500 31.750 79.845 31.750
                 31.750 79.845 31.750 115.500 33.080 115.500 33.080 118.000
                 31.750 118.000 31.750 120.000 28.250 120.000 28.250 78.255 78.255 28.250
                 115.500 28.250 115.500 27.250 77.800 27.250 27.250 77.800 27.250 115.500
                 28.250 115.500 28.250 118.000 27.250 118.000 27.250 120.000
                 23.750 120.000 23.750 76.205 76.205 23.750 115.500 23.750 115.500 22.750
                 75.750 22.750 22.750 75.750 22.750 115.500 23.750 115.500 23.750 118.000
                 22.750 118.000 22.750 120.000 19.250 120.000 19.250 74.160 74.160 19.250
                 115.500 19.250 115.500 18.250 73.705 18.250 18.250 73.705 18.250 115.500
                 19.250 115.500 19.250 118.000 18.250 118.000 18.250 120.000
                 14.750 120.000 14.750 72.110 72.110 14.750 115.500 14.750 115.500 13.750
                 71.655 13.750 13.750 71.655 13.750 115.500 14.750 115.500 14.750 118.000
                 13.750 118.000 13.750 120.000 10.250 120.000 10.250 70.065 70.065 10.250
                 115.500 10.250 115.500 9.250 69.610 9.250 9.250 69.610 9.250 115.500
                 10.250 115.500 10.250 118.000 9.250 118.000 9.250 120.000 5.750 120.000
                 5.750 118.000 4.750 118.000 4.750 120.000 1.250 120.000 ;
        LAYER M6 ;
                POLYGON  1.250 115.500 5.750 115.500 5.750 68.515 68.515 5.750 115.500 5.750
                 115.500 1.250 120.000 1.250 120.000 4.750 118.000 4.750 118.000 5.750
                 120.000 5.750 120.000 9.250 118.000 9.250 118.000 10.250 120.000 10.250
                 120.000 13.750 118.000 13.750 118.000 14.750 120.000 14.750
                 120.000 18.250 118.000 18.250 118.000 19.250 120.000 19.250
                 120.000 22.750 118.000 22.750 118.000 23.750 120.000 23.750
                 120.000 27.250 118.000 27.250 118.000 28.250 120.000 28.250
                 120.000 31.750 118.000 31.750 118.000 33.080 120.000 33.080
                 120.000 37.580 82.500 37.580 37.580 82.500 37.580 120.000 33.080 120.000
                 33.080 80.650 80.650 33.080 115.500 33.080 115.500 31.750 79.845 31.750
                 31.750 79.845 31.750 115.500 33.080 115.500 33.080 118.000
                 31.750 118.000 31.750 120.000 28.250 120.000 28.250 78.255 78.255 28.250
                 115.500 28.250 115.500 27.250 77.800 27.250 27.250 77.800 27.250 115.500
                 28.250 115.500 28.250 118.000 27.250 118.000 27.250 120.000
                 23.750 120.000 23.750 76.205 76.205 23.750 115.500 23.750 115.500 22.750
                 75.750 22.750 22.750 75.750 22.750 115.500 23.750 115.500 23.750 118.000
                 22.750 118.000 22.750 120.000 19.250 120.000 19.250 74.160 74.160 19.250
                 115.500 19.250 115.500 18.250 73.705 18.250 18.250 73.705 18.250 115.500
                 19.250 115.500 19.250 118.000 18.250 118.000 18.250 120.000
                 14.750 120.000 14.750 72.110 72.110 14.750 115.500 14.750 115.500 13.750
                 71.655 13.750 13.750 71.655 13.750 115.500 14.750 115.500 14.750 118.000
                 13.750 118.000 13.750 120.000 10.250 120.000 10.250 70.065 70.065 10.250
                 115.500 10.250 115.500 9.250 69.610 9.250 9.250 69.610 9.250 115.500
                 10.250 115.500 10.250 118.000 9.250 118.000 9.250 120.000 5.750 120.000
                 5.750 118.000 4.750 118.000 4.750 120.000 1.250 120.000 ;
        LAYER M5 ;
                POLYGON  1.250 115.500 5.750 115.500 5.750 68.515 68.515 5.750 115.500 5.750
                 115.500 1.250 120.000 1.250 120.000 4.750 118.000 4.750 118.000 5.750
                 120.000 5.750 120.000 9.250 118.000 9.250 118.000 10.250 120.000 10.250
                 120.000 13.750 118.000 13.750 118.000 14.750 120.000 14.750
                 120.000 18.250 118.000 18.250 118.000 19.250 120.000 19.250
                 120.000 22.750 118.000 22.750 118.000 23.750 120.000 23.750
                 120.000 27.250 118.000 27.250 118.000 28.250 120.000 28.250
                 120.000 31.750 118.000 31.750 118.000 33.080 120.000 33.080
                 120.000 37.580 82.500 37.580 37.580 82.500 37.580 120.000 33.080 120.000
                 33.080 80.650 80.650 33.080 115.500 33.080 115.500 31.750 79.845 31.750
                 31.750 79.845 31.750 115.500 33.080 115.500 33.080 118.000
                 31.750 118.000 31.750 120.000 28.250 120.000 28.250 78.255 78.255 28.250
                 115.500 28.250 115.500 27.250 77.800 27.250 27.250 77.800 27.250 115.500
                 28.250 115.500 28.250 118.000 27.250 118.000 27.250 120.000
                 23.750 120.000 23.750 76.205 76.205 23.750 115.500 23.750 115.500 22.750
                 75.750 22.750 22.750 75.750 22.750 115.500 23.750 115.500 23.750 118.000
                 22.750 118.000 22.750 120.000 19.250 120.000 19.250 74.160 74.160 19.250
                 115.500 19.250 115.500 18.250 73.705 18.250 18.250 73.705 18.250 115.500
                 19.250 115.500 19.250 118.000 18.250 118.000 18.250 120.000
                 14.750 120.000 14.750 72.110 72.110 14.750 115.500 14.750 115.500 13.750
                 71.655 13.750 13.750 71.655 13.750 115.500 14.750 115.500 14.750 118.000
                 13.750 118.000 13.750 120.000 10.250 120.000 10.250 70.065 70.065 10.250
                 115.500 10.250 115.500 9.250 69.610 9.250 9.250 69.610 9.250 115.500
                 10.250 115.500 10.250 118.000 9.250 118.000 9.250 120.000 5.750 120.000
                 5.750 118.000 4.750 118.000 4.750 120.000 1.250 120.000 ;
        LAYER M4 ;
                POLYGON  1.250 115.500 5.750 115.500 5.750 68.515 68.515 5.750 115.500 5.750
                 115.500 1.250 120.000 1.250 120.000 4.750 118.000 4.750 118.000 5.750
                 120.000 5.750 120.000 9.250 118.000 9.250 118.000 10.250 120.000 10.250
                 120.000 13.750 118.000 13.750 118.000 14.750 120.000 14.750
                 120.000 18.250 118.000 18.250 118.000 19.250 120.000 19.250
                 120.000 22.750 118.000 22.750 118.000 23.750 120.000 23.750
                 120.000 27.250 118.000 27.250 118.000 28.250 120.000 28.250
                 120.000 31.750 118.000 31.750 118.000 33.080 120.000 33.080
                 120.000 37.580 82.500 37.580 37.580 82.500 37.580 120.000 33.080 120.000
                 33.080 80.650 80.650 33.080 115.500 33.080 115.500 31.750 79.845 31.750
                 31.750 79.845 31.750 115.500 33.080 115.500 33.080 118.000
                 31.750 118.000 31.750 120.000 28.250 120.000 28.250 78.255 78.255 28.250
                 115.500 28.250 115.500 27.250 77.800 27.250 27.250 77.800 27.250 115.500
                 28.250 115.500 28.250 118.000 27.250 118.000 27.250 120.000
                 23.750 120.000 23.750 76.205 76.205 23.750 115.500 23.750 115.500 22.750
                 75.750 22.750 22.750 75.750 22.750 115.500 23.750 115.500 23.750 118.000
                 22.750 118.000 22.750 120.000 19.250 120.000 19.250 74.160 74.160 19.250
                 115.500 19.250 115.500 18.250 73.705 18.250 18.250 73.705 18.250 115.500
                 19.250 115.500 19.250 118.000 18.250 118.000 18.250 120.000
                 14.750 120.000 14.750 72.110 72.110 14.750 115.500 14.750 115.500 13.750
                 71.655 13.750 13.750 71.655 13.750 115.500 14.750 115.500 14.750 118.000
                 13.750 118.000 13.750 120.000 10.250 120.000 10.250 70.065 70.065 10.250
                 115.500 10.250 115.500 9.250 69.610 9.250 9.250 69.610 9.250 115.500
                 10.250 115.500 10.250 118.000 9.250 118.000 9.250 120.000 5.750 120.000
                 5.750 118.000 4.750 118.000 4.750 120.000 1.250 120.000 ;
        LAYER M3 ;
                POLYGON  1.250 115.500 5.750 115.500 5.750 68.515 68.515 5.750 115.500 5.750
                 115.500 1.250 120.000 1.250 120.000 4.750 118.000 4.750 118.000 5.750
                 120.000 5.750 120.000 9.250 118.000 9.250 118.000 10.250 120.000 10.250
                 120.000 13.750 118.000 13.750 118.000 14.750 120.000 14.750
                 120.000 18.250 118.000 18.250 118.000 19.250 120.000 19.250
                 120.000 22.750 118.000 22.750 118.000 23.750 120.000 23.750
                 120.000 27.250 118.000 27.250 118.000 28.250 120.000 28.250
                 120.000 31.750 118.000 31.750 118.000 33.080 120.000 33.080
                 120.000 37.580 82.500 37.580 37.580 82.500 37.580 120.000 33.080 120.000
                 33.080 80.650 80.650 33.080 115.500 33.080 115.500 31.750 79.845 31.750
                 31.750 79.845 31.750 115.500 33.080 115.500 33.080 118.000
                 31.750 118.000 31.750 120.000 28.250 120.000 28.250 78.255 78.255 28.250
                 115.500 28.250 115.500 27.250 77.800 27.250 27.250 77.800 27.250 115.500
                 28.250 115.500 28.250 118.000 27.250 118.000 27.250 120.000
                 23.750 120.000 23.750 76.205 76.205 23.750 115.500 23.750 115.500 22.750
                 75.750 22.750 22.750 75.750 22.750 115.500 23.750 115.500 23.750 118.000
                 22.750 118.000 22.750 120.000 19.250 120.000 19.250 74.160 74.160 19.250
                 115.500 19.250 115.500 18.250 73.705 18.250 18.250 73.705 18.250 115.500
                 19.250 115.500 19.250 118.000 18.250 118.000 18.250 120.000
                 14.750 120.000 14.750 72.110 72.110 14.750 115.500 14.750 115.500 13.750
                 71.655 13.750 13.750 71.655 13.750 115.500 14.750 115.500 14.750 118.000
                 13.750 118.000 13.750 120.000 10.250 120.000 10.250 70.065 70.065 10.250
                 115.500 10.250 115.500 9.250 69.610 9.250 9.250 69.610 9.250 115.500
                 10.250 115.500 10.250 118.000 9.250 118.000 9.250 120.000 5.750 120.000
                 5.750 118.000 4.750 118.000 4.750 120.000 1.250 120.000 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
        LAYER M5 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
        LAYER M6 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
        LAYER M7 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
        LAYER M4 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
        LAYER M5 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
        LAYER M6 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
        LAYER M7 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
        LAYER M3 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
        LAYER M4 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
        LAYER M5 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
        LAYER M6 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
        LAYER M7 ;
                POLYGON  88.020 105.450 105.450 88.020 120.000 88.020 120.000 91.520
                 107.040 91.520 91.520 107.040 91.520 120.000 88.020 120.000 ;
        LAYER M3 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
        LAYER M4 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
        LAYER M5 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
        LAYER M6 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
        LAYER M7 ;
                POLYGON  92.370 107.430 107.430 92.370 120.000 92.370 120.000 95.870
                 109.020 95.870 95.870 109.020 95.870 120.000 92.370 120.000 ;
                POLYGON  96.720 109.410 109.410 96.720 120.000 96.720 120.000 100.220
                 111.000 100.220 100.220 111.000 100.220 120.000 96.720 120.000 ;
                POLYGON  101.070 111.385 111.385 101.070 120.000 101.070 120.000 104.570
                 112.980 104.570 104.570 112.980 104.570 120.000 101.070 120.000 ;
                POLYGON  105.420 113.365 113.365 105.420 120.000 105.420 120.000 108.920
                 114.960 108.920 108.920 114.960 108.920 120.000 105.420 120.000 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M6 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M5 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M4 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        LAYER M3 ;
                POLYGON  83.670 103.470 103.470 83.670 120.000 83.670 120.000 87.170
                 105.060 87.170 87.170 105.060 87.170 120.000 83.670 120.000 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M6 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M5 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M4 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        LAYER M3 ;
                POLYGON  79.975 101.790 101.790 79.975 120.000 79.975 120.000 82.975
                 103.155 82.975 82.975 103.155 82.975 120.000 79.975 120.000 ;
                POLYGON  72.475 98.375 98.375 72.475 120.000 72.475 120.000 75.975 99.970 75.975
                 75.975 99.970 75.975 120.000 72.475 120.000 ;
                POLYGON  67.975 96.330 96.330 67.975 120.000 67.975 120.000 71.475 97.920 71.475
                 71.475 97.920 71.475 120.000 67.975 120.000 ;
                POLYGON  63.475 94.280 94.280 63.475 120.000 63.475 120.000 66.975 95.875 66.975
                 66.975 95.875 66.975 120.000 63.475 120.000 ;
                POLYGON  58.975 92.235 92.235 58.975 120.000 58.975 120.000 62.475 93.825 62.475
                 62.475 93.825 62.475 120.000 58.975 120.000 ;
                POLYGON  54.475 90.185 90.185 54.475 120.000 54.475 120.000 57.975 91.780 57.975
                 57.975 91.780 57.975 120.000 54.475 120.000 ;
                POLYGON  49.975 88.140 88.140 49.975 120.000 49.975 120.000 53.475 89.730 53.475
                 53.475 89.730 53.475 120.000 49.975 120.000 ;
                POLYGON  45.475 86.090 86.090 45.475 120.000 45.475 120.000 48.975 87.685 48.975
                 48.975 87.685 48.975 120.000 45.475 120.000 ;
                POLYGON  40.975 84.045 84.045 40.975 120.000 40.975 120.000 44.475 85.635 44.475
                 44.475 85.635 44.475 120.000 40.975 120.000 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  114.010 117.275 117.275 114.010 120.000 114.010 120.000 117.510
                 118.865 117.510 117.510 118.865 117.510 120.000 114.010 120.000 ;
                POLYGON  109.770 115.345 115.345 109.770 120.000 109.770 120.000 113.270
                 116.940 113.270 113.270 116.940 113.270 120.000 109.770 120.000 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  118.010 119.095 119.095 118.010 120.000 118.010 120.000 118.500
                 119.320 118.500 118.500 119.320 118.500 120.000 118.010 120.000 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA1 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 0.000 120.000 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 120.000 120.000 ;
    END
END PCORNER_G

MACRO PDB3AC_G
    CLASS PAD ;
    FOREIGN PDB3AC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AIO
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M2 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        LAYER M1 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        END
        ANTENNADIFFAREA 300.0000 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 1442.2320 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 257.2500 LAYER VIA1 ;
        ANTENNADIFFAREA 300.0000 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 1442.2320 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 6.1740 LAYER VIA2 ;
        ANTENNADIFFAREA 300.0000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.7200 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 300.0000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 300.0000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 300.0000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 300.0000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END AIO
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TACVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TACVSS
    PIN TACVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TACVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDB3AC_G

MACRO PDB3A_G
    CLASS PAD ;
    FOREIGN PDB3A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN AIO
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M2 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        LAYER M1 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        END
        ANTENNADIFFAREA 300.0000 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 1442.2320 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 257.2500 LAYER VIA1 ;
        ANTENNADIFFAREA 300.0000 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 1442.2320 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 6.1740 LAYER VIA2 ;
        ANTENNADIFFAREA 300.0000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.7200 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 300.0000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 300.0000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 300.0000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 300.0000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END AIO
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  20.220 118.200 22.620 120.000 ;
        RECT  15.760 118.200 18.160 120.000 ;
        RECT  11.300 118.200 13.700 120.000 ;
        RECT  6.840 118.200 9.240 120.000 ;
        RECT  2.380 118.200 4.780 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDB3A_G

MACRO PDDW04DGZ_G
    CLASS PAD ;
    FOREIGN PDDW04DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW04DGZ_G

MACRO PDDW04SDGZ_G
    CLASS PAD ;
    FOREIGN PDDW04SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW04SDGZ_G

MACRO PDDW08DGZ_G
    CLASS PAD ;
    FOREIGN PDDW08DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW08DGZ_G

MACRO PDDW08SDGZ_G
    CLASS PAD ;
    FOREIGN PDDW08SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW08SDGZ_G

MACRO PDDW12DGZ_G
    CLASS PAD ;
    FOREIGN PDDW12DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW12DGZ_G

MACRO PDDW12SDGZ_G
    CLASS PAD ;
    FOREIGN PDDW12SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW12SDGZ_G

MACRO PDDW16DGZ_G
    CLASS PAD ;
    FOREIGN PDDW16DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW16DGZ_G

MACRO PDDW16SDGZ_G
    CLASS PAD ;
    FOREIGN PDDW16SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDDW16SDGZ_G

MACRO PDUW04DGZ_G
    CLASS PAD ;
    FOREIGN PDUW04DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW04DGZ_G

MACRO PDUW04SDGZ_G
    CLASS PAD ;
    FOREIGN PDUW04SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW04SDGZ_G

MACRO PDUW08DGZ_G
    CLASS PAD ;
    FOREIGN PDUW08DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW08DGZ_G

MACRO PDUW08SDGZ_G
    CLASS PAD ;
    FOREIGN PDUW08SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW08SDGZ_G

MACRO PDUW12DGZ_G
    CLASS PAD ;
    FOREIGN PDUW12DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW12DGZ_G

MACRO PDUW12SDGZ_G
    CLASS PAD ;
    FOREIGN PDUW12SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW12SDGZ_G

MACRO PDUW16DGZ_G
    CLASS PAD ;
    FOREIGN PDUW16DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW16DGZ_G

MACRO PDUW16SDGZ_G
    CLASS PAD ;
    FOREIGN PDUW16SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PDUW16SDGZ_G

MACRO PDXOE1DG_G
    CLASS PAD ;
    FOREIGN PDXOE1DG_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M6 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M5 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M4 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M3 ;
        RECT  27.385 76.475 47.615 79.475 ;
        END
        ANTENNAGATEAREA 18.2600 LAYER M3 ;
        ANTENNADIFFAREA 702.1490 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAMAXAREACAR 55.3522 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.7971 LAYER VIA3 ;
        ANTENNAGATEAREA 18.2600 LAYER M4 ;
        ANTENNADIFFAREA 702.1490 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 58.6758 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4057 LAYER VIA4 ;
        ANTENNAGATEAREA 18.2600 LAYER M5 ;
        ANTENNADIFFAREA 702.1490 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 61.9995 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.0143 LAYER VIA5 ;
        ANTENNAGATEAREA 18.2600 LAYER M6 ;
        ANTENNADIFFAREA 702.1490 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 65.3232 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.6229 LAYER VIA6 ;
        ANTENNAGATEAREA 18.2600 LAYER M7 ;
        ANTENNADIFFAREA 702.1490 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 68.6468 LAYER M7 ;
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNAGATEAREA 88.2000 LAYER M3 ;
        ANTENNADIFFAREA 906.5000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 62.5945 LAYER M3 ;
        ANTENNAMAXAREACAR 1.3120 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.1269 LAYER VIA3 ;
        ANTENNAGATEAREA 88.2000 LAYER M4 ;
        ANTENNADIFFAREA 906.5000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 2.0001 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.2529 LAYER VIA4 ;
        ANTENNAGATEAREA 88.2000 LAYER M5 ;
        ANTENNADIFFAREA 906.5000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 2.6882 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.3789 LAYER VIA5 ;
        ANTENNAGATEAREA 88.2000 LAYER M6 ;
        ANTENNADIFFAREA 906.5000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 3.3763 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.5049 LAYER VIA6 ;
        ANTENNAGATEAREA 88.2000 LAYER M7 ;
        ANTENNADIFFAREA 906.5000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 4.0644 LAYER M7 ;
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M6 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M5 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M4 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M3 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M2 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        END
        ANTENNADIFFAREA 4.1300 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.7417 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5782 LAYER VIA1 ;
        ANTENNADIFFAREA 4.1300 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.5038 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 4.1300 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 4.1300 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 4.1300 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 4.1300 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 4.1300 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M6 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M5 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M4 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M3 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M1 ;
        RECT  26.525 119.000 29.415 120.000 ;
        END
        ANTENNAGATEAREA 8.3000 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 9.6527 LAYER M1 ;
        ANTENNAMAXAREACAR 1.1630 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNAMAXAREACAR 0.0638 LAYER VIA1 ;
        ANTENNAGATEAREA 8.3000 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAMAXAREACAR 1.5112 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 0.1275 LAYER VIA2 ;
        ANTENNAGATEAREA 8.3000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 1.8594 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.1913 LAYER VIA3 ;
        ANTENNAGATEAREA 8.3000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 2.2076 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.2550 LAYER VIA4 ;
        ANTENNAGATEAREA 8.3000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 2.5558 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.3188 LAYER VIA5 ;
        ANTENNAGATEAREA 8.3000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 2.9039 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.3826 LAYER VIA6 ;
        ANTENNAGATEAREA 8.3000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 3.2521 LAYER M7 ;
    END E
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 36.120 31.750 36.120 4.750 13.880 4.750
                 13.880 5.750 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250
                 36.120 10.250 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750
                 36.120 18.250 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750
                 13.880 22.750 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250
                 13.880 28.250 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080
                 50.000 33.080 50.000 37.580 49.075 37.580 49.075 40.710 48.745 40.710
                 48.745 37.580 45.445 37.580 45.445 40.230 44.955 40.230 44.955 37.580
                 39.285 37.580 39.285 40.230 38.795 40.230 38.795 37.580 33.125 37.580
                 33.125 40.230 32.635 40.230 32.635 37.580 25.735 37.580 25.735 40.710
                 25.565 40.710 25.565 37.580 24.085 37.580 24.085 40.710 23.755 40.710
                 23.755 37.580 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580
                 14.285 37.580 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580
                 8.125 40.230 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710
                 0.945 40.710 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080
                 11.120 31.750 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250
                 0.000 27.250 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750
                 0.000 19.250 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750
                 11.120 14.750 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250
                 11.120 9.250 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 36.120 108.920 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 29.555 40.975 29.555 39.450 30.045 39.450 30.045 40.975
                 35.715 40.975 35.715 39.450 36.205 39.450 36.205 40.975 41.875 40.975
                 41.875 39.450 42.365 39.450 42.365 40.975 49.225 40.975 49.225 39.450
                 49.395 39.450 49.395 40.975 50.000 40.975 50.000 44.475 38.880 44.475
                 38.880 45.475 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975
                 50.000 49.975 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475
                 50.000 57.975 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475
                 38.880 62.475 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975
                 38.880 67.975 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475
                 50.000 72.475 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475
                 13.880 45.475 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975
                 36.120 49.975 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475
                 36.120 57.975 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475
                 13.880 62.475 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975
                 13.880 67.975 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475
                 36.120 72.475 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 50.000 109.770 50.000 113.270 38.880 113.270
                 38.880 114.010 50.000 114.010 50.000 117.510 36.120 117.510
                 36.120 113.270 13.880 113.270 13.880 114.010 36.120 114.010
                 36.120 117.510 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270
                 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 50.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA2 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  0.000 118.010 50.000 118.500 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.795 33.080 39.285 40.230 ;
        RECT  36.120 1.250 38.880 31.750 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 108.920 ;
        RECT  36.120 109.770 38.880 117.510 ;
        RECT  33.125 33.080 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA3 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.880 33.080 39.285 40.230 ;
        RECT  38.795 1.250 38.880 40.230 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  36.120 1.250 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  33.125 33.080 36.120 37.580 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA4 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA5 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA6 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 50.000 120.000 ;
    END
END PDXOE1DG_G

MACRO PDXOE2DG_G
    CLASS PAD ;
    FOREIGN PDXOE2DG_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M6 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M5 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M4 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M3 ;
        RECT  27.385 76.475 47.615 79.475 ;
        END
        ANTENNAGATEAREA 18.2600 LAYER M3 ;
        ANTENNADIFFAREA 702.1490 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAMAXAREACAR 55.3522 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.7971 LAYER VIA3 ;
        ANTENNAGATEAREA 18.2600 LAYER M4 ;
        ANTENNADIFFAREA 702.1490 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 58.6758 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4057 LAYER VIA4 ;
        ANTENNAGATEAREA 18.2600 LAYER M5 ;
        ANTENNADIFFAREA 702.1490 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 61.9995 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.0143 LAYER VIA5 ;
        ANTENNAGATEAREA 18.2600 LAYER M6 ;
        ANTENNADIFFAREA 702.1490 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 65.3232 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.6229 LAYER VIA6 ;
        ANTENNAGATEAREA 18.2600 LAYER M7 ;
        ANTENNADIFFAREA 702.1490 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 68.6468 LAYER M7 ;
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNAGATEAREA 161.0000 LAYER M3 ;
        ANTENNADIFFAREA 906.5000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 64.1587 LAYER M3 ;
        ANTENNAMAXAREACAR 0.9328 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.0700 LAYER VIA3 ;
        ANTENNAGATEAREA 161.0000 LAYER M4 ;
        ANTENNADIFFAREA 906.5000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 1.3097 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.1390 LAYER VIA4 ;
        ANTENNAGATEAREA 161.0000 LAYER M5 ;
        ANTENNADIFFAREA 906.5000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 1.6867 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.2080 LAYER VIA5 ;
        ANTENNAGATEAREA 161.0000 LAYER M6 ;
        ANTENNADIFFAREA 906.5000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 2.0636 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.2770 LAYER VIA6 ;
        ANTENNAGATEAREA 161.0000 LAYER M7 ;
        ANTENNADIFFAREA 906.5000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 2.4406 LAYER M7 ;
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M6 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M5 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M4 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M3 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M2 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        END
        ANTENNADIFFAREA 4.1300 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.7417 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5782 LAYER VIA1 ;
        ANTENNADIFFAREA 4.1300 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.5038 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 4.1300 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 4.1300 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 4.1300 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 4.1300 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 4.1300 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M6 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M5 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M4 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M3 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M1 ;
        RECT  26.525 119.000 29.415 120.000 ;
        END
        ANTENNAGATEAREA 8.3000 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 9.6527 LAYER M1 ;
        ANTENNAMAXAREACAR 1.1630 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNAMAXAREACAR 0.0638 LAYER VIA1 ;
        ANTENNAGATEAREA 8.3000 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAMAXAREACAR 1.5112 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 0.1275 LAYER VIA2 ;
        ANTENNAGATEAREA 8.3000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 1.8594 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.1913 LAYER VIA3 ;
        ANTENNAGATEAREA 8.3000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 2.2076 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.2550 LAYER VIA4 ;
        ANTENNAGATEAREA 8.3000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 2.5558 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.3188 LAYER VIA5 ;
        ANTENNAGATEAREA 8.3000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 2.9039 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.3826 LAYER VIA6 ;
        ANTENNAGATEAREA 8.3000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 3.2521 LAYER M7 ;
    END E
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 36.120 31.750 36.120 4.750 13.880 4.750
                 13.880 5.750 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250
                 36.120 10.250 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750
                 36.120 18.250 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750
                 13.880 22.750 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250
                 13.880 28.250 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080
                 50.000 33.080 50.000 37.580 49.075 37.580 49.075 40.710 48.745 40.710
                 48.745 37.580 45.445 37.580 45.445 40.230 44.955 40.230 44.955 37.580
                 39.285 37.580 39.285 40.230 38.795 40.230 38.795 37.580 33.125 37.580
                 33.125 40.230 32.635 40.230 32.635 37.580 25.735 37.580 25.735 40.710
                 25.565 40.710 25.565 37.580 24.085 37.580 24.085 40.710 23.755 40.710
                 23.755 37.580 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580
                 14.285 37.580 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580
                 8.125 40.230 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710
                 0.945 40.710 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080
                 11.120 31.750 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250
                 0.000 27.250 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750
                 0.000 19.250 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750
                 11.120 14.750 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250
                 11.120 9.250 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 36.120 108.920 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 29.555 40.975 29.555 39.450 30.045 39.450 30.045 40.975
                 35.715 40.975 35.715 39.450 36.205 39.450 36.205 40.975 41.875 40.975
                 41.875 39.450 42.365 39.450 42.365 40.975 49.225 40.975 49.225 39.450
                 49.395 39.450 49.395 40.975 50.000 40.975 50.000 44.475 38.880 44.475
                 38.880 45.475 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975
                 50.000 49.975 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475
                 50.000 57.975 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475
                 38.880 62.475 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975
                 38.880 67.975 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475
                 50.000 72.475 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475
                 13.880 45.475 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975
                 36.120 49.975 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475
                 36.120 57.975 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475
                 13.880 62.475 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975
                 13.880 67.975 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475
                 36.120 72.475 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 50.000 109.770 50.000 113.270 38.880 113.270
                 38.880 114.010 50.000 114.010 50.000 117.510 36.120 117.510
                 36.120 113.270 13.880 113.270 13.880 114.010 36.120 114.010
                 36.120 117.510 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270
                 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 50.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA2 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  0.000 118.010 50.000 118.500 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.795 33.080 39.285 40.230 ;
        RECT  36.120 1.250 38.880 31.750 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 108.920 ;
        RECT  36.120 109.770 38.880 117.510 ;
        RECT  33.125 33.080 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA3 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.880 33.080 39.285 40.230 ;
        RECT  38.795 1.250 38.880 40.230 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  36.120 1.250 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  33.125 33.080 36.120 37.580 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA4 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA5 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA6 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 50.000 120.000 ;
    END
END PDXOE2DG_G

MACRO PDXOE3DG_G
    CLASS PAD ;
    FOREIGN PDXOE3DG_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN XOUT
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M6 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M5 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M4 ;
        RECT  27.385 76.475 47.615 79.475 ;
        LAYER M3 ;
        RECT  27.385 76.475 47.615 79.475 ;
        END
        ANTENNAGATEAREA 18.2600 LAYER M3 ;
        ANTENNADIFFAREA 702.1490 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAMAXAREACAR 55.3522 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.7971 LAYER VIA3 ;
        ANTENNAGATEAREA 18.2600 LAYER M4 ;
        ANTENNADIFFAREA 702.1490 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 58.6758 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4057 LAYER VIA4 ;
        ANTENNAGATEAREA 18.2600 LAYER M5 ;
        ANTENNADIFFAREA 702.1490 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 61.9995 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.0143 LAYER VIA5 ;
        ANTENNAGATEAREA 18.2600 LAYER M6 ;
        ANTENNADIFFAREA 702.1490 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 65.3232 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.6229 LAYER VIA6 ;
        ANTENNAGATEAREA 18.2600 LAYER M7 ;
        ANTENNADIFFAREA 702.1490 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 68.6468 LAYER M7 ;
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNAGATEAREA 249.2000 LAYER M3 ;
        ANTENNADIFFAREA 906.5000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 65.7229 LAYER M3 ;
        ANTENNAMAXAREACAR 0.7524 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.0455 LAYER VIA3 ;
        ANTENNAGATEAREA 249.2000 LAYER M4 ;
        ANTENNADIFFAREA 906.5000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAMAXAREACAR 0.9960 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.0901 LAYER VIA4 ;
        ANTENNAGATEAREA 249.2000 LAYER M5 ;
        ANTENNADIFFAREA 906.5000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAMAXAREACAR 1.2395 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.1347 LAYER VIA5 ;
        ANTENNAGATEAREA 249.2000 LAYER M6 ;
        ANTENNADIFFAREA 906.5000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAMAXAREACAR 1.4831 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.1793 LAYER VIA6 ;
        ANTENNAGATEAREA 249.2000 LAYER M7 ;
        ANTENNADIFFAREA 906.5000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
        ANTENNAMAXAREACAR 1.7266 LAYER M7 ;
    END XIN
    PIN XC
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M6 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M5 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M4 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M3 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M2 ;
        RECT  34.665 119.000 37.555 120.000 ;
        LAYER M1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        END
        ANTENNADIFFAREA 4.1300 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.7417 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5782 LAYER VIA1 ;
        ANTENNADIFFAREA 4.1300 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.5038 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 4.1300 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 4.1300 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 4.1300 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 4.1300 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 4.1300 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END XC
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M6 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M5 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M4 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M3 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M1 ;
        RECT  26.525 119.000 29.415 120.000 ;
        END
        ANTENNAGATEAREA 8.3000 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 9.6527 LAYER M1 ;
        ANTENNAMAXAREACAR 1.1630 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNAMAXAREACAR 0.0638 LAYER VIA1 ;
        ANTENNAGATEAREA 8.3000 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAMAXAREACAR 1.5112 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 0.1275 LAYER VIA2 ;
        ANTENNAGATEAREA 8.3000 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 1.8594 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 0.1913 LAYER VIA3 ;
        ANTENNAGATEAREA 8.3000 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 2.2076 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 0.2550 LAYER VIA4 ;
        ANTENNAGATEAREA 8.3000 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 2.5558 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 0.3188 LAYER VIA5 ;
        ANTENNAGATEAREA 8.3000 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 2.9039 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 0.3826 LAYER VIA6 ;
        ANTENNAGATEAREA 8.3000 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 3.2521 LAYER M7 ;
    END E
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 38.880 31.750 38.880 33.080 50.000 33.080
                 50.000 37.580 36.120 37.580 36.120 4.750 13.880 4.750 13.880 5.750
                 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250 36.120 10.250
                 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750 36.120 18.250
                 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750 13.880 22.750
                 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250 13.880 28.250
                 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080 36.120 33.080
                 36.120 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 50.000 1.250 50.000 4.750 38.880 4.750 38.880 5.750
                 50.000 5.750 50.000 9.250 38.880 9.250 38.880 10.250 50.000 10.250
                 50.000 13.750 38.880 13.750 38.880 14.750 50.000 14.750 50.000 18.250
                 38.880 18.250 38.880 19.250 50.000 19.250 50.000 22.750 38.880 22.750
                 38.880 23.750 50.000 23.750 50.000 27.250 38.880 27.250 38.880 28.250
                 50.000 28.250 50.000 31.750 36.120 31.750 36.120 4.750 13.880 4.750
                 13.880 5.750 36.120 5.750 36.120 9.250 13.880 9.250 13.880 10.250
                 36.120 10.250 36.120 13.750 13.880 13.750 13.880 14.750 36.120 14.750
                 36.120 18.250 13.880 18.250 13.880 19.250 36.120 19.250 36.120 22.750
                 13.880 22.750 13.880 23.750 36.120 23.750 36.120 27.250 13.880 27.250
                 13.880 28.250 36.120 28.250 36.120 31.750 13.880 31.750 13.880 33.080
                 50.000 33.080 50.000 37.580 49.075 37.580 49.075 40.710 48.745 40.710
                 48.745 37.580 45.445 37.580 45.445 40.230 44.955 40.230 44.955 37.580
                 39.285 37.580 39.285 40.230 38.795 40.230 38.795 37.580 33.125 37.580
                 33.125 40.230 32.635 40.230 32.635 37.580 25.735 37.580 25.735 40.710
                 25.565 40.710 25.565 37.580 24.085 37.580 24.085 40.710 23.755 40.710
                 23.755 37.580 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580
                 14.285 37.580 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580
                 8.125 40.230 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710
                 0.945 40.710 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080
                 11.120 31.750 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250
                 0.000 27.250 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750
                 0.000 19.250 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750
                 11.120 14.750 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250
                 11.120 9.250 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 38.880 108.920 38.880 109.770 50.000 109.770 50.000 113.270
                 38.880 113.270 38.880 114.010 50.000 114.010 50.000 117.510
                 36.120 117.510 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 13.880 108.920
                 13.880 109.770 36.120 109.770 36.120 113.270 13.880 113.270
                 13.880 114.010 36.120 114.010 36.120 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 0.000 109.770 11.120 109.770
                 11.120 108.920 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570
                 0.000 104.570 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220
                 0.000 96.720 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370
                 11.120 92.370 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020
                 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 50.000 83.670 50.000 87.170 38.880 87.170 38.880 88.020
                 50.000 88.020 50.000 91.520 38.880 91.520 38.880 92.370 50.000 92.370
                 50.000 95.870 38.880 95.870 38.880 96.720 50.000 96.720 50.000 100.220
                 38.880 100.220 38.880 101.070 50.000 101.070 50.000 104.570
                 38.880 104.570 38.880 105.420 50.000 105.420 50.000 108.920
                 36.120 108.920 36.120 87.170 13.880 87.170 13.880 88.020 36.120 88.020
                 36.120 91.520 13.880 91.520 13.880 92.370 36.120 92.370 36.120 95.870
                 13.880 95.870 13.880 96.720 36.120 96.720 36.120 100.220 13.880 100.220
                 13.880 101.070 36.120 101.070 36.120 104.570 13.880 104.570
                 13.880 105.420 36.120 105.420 36.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 50.000 40.975 50.000 44.475 38.880 44.475 38.880 45.475
                 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975 50.000 49.975
                 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475 50.000 57.975
                 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475 38.880 62.475
                 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975 38.880 67.975
                 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475 50.000 72.475
                 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475 13.880 45.475
                 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975 36.120 49.975
                 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475 36.120 57.975
                 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475 13.880 62.475
                 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975 13.880 67.975
                 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475 36.120 72.475
                 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 50.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 29.555 40.975 29.555 39.450 30.045 39.450 30.045 40.975
                 35.715 40.975 35.715 39.450 36.205 39.450 36.205 40.975 41.875 40.975
                 41.875 39.450 42.365 39.450 42.365 40.975 49.225 40.975 49.225 39.450
                 49.395 39.450 49.395 40.975 50.000 40.975 50.000 44.475 38.880 44.475
                 38.880 45.475 50.000 45.475 50.000 48.975 38.880 48.975 38.880 49.975
                 50.000 49.975 50.000 53.475 38.880 53.475 38.880 54.475 50.000 54.475
                 50.000 57.975 38.880 57.975 38.880 58.975 50.000 58.975 50.000 62.475
                 38.880 62.475 38.880 63.475 50.000 63.475 50.000 66.975 38.880 66.975
                 38.880 67.975 50.000 67.975 50.000 71.475 38.880 71.475 38.880 72.475
                 50.000 72.475 50.000 75.975 36.120 75.975 36.120 44.475 13.880 44.475
                 13.880 45.475 36.120 45.475 36.120 48.975 13.880 48.975 13.880 49.975
                 36.120 49.975 36.120 53.475 13.880 53.475 13.880 54.475 36.120 54.475
                 36.120 57.975 13.880 57.975 13.880 58.975 36.120 58.975 36.120 62.475
                 13.880 62.475 13.880 63.475 36.120 63.475 36.120 66.975 13.880 66.975
                 13.880 67.975 36.120 67.975 36.120 71.475 13.880 71.475 13.880 72.475
                 36.120 72.475 36.120 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 50.000 109.770 50.000 113.270 38.880 113.270
                 38.880 114.010 50.000 114.010 50.000 117.510 36.120 117.510
                 36.120 113.270 13.880 113.270 13.880 114.010 36.120 114.010
                 36.120 117.510 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270
                 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 50.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA1 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  26.525 119.000 29.415 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA2 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  0.000 118.010 50.000 118.500 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.795 33.080 39.285 40.230 ;
        RECT  36.120 1.250 38.880 31.750 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 108.920 ;
        RECT  36.120 109.770 38.880 117.510 ;
        RECT  33.125 33.080 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA3 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  49.075 33.080 50.000 37.580 ;
        RECT  49.395 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  49.225 39.450 49.395 44.475 ;
        RECT  42.365 40.975 49.225 44.475 ;
        RECT  48.745 33.080 49.075 40.710 ;
        RECT  45.445 33.080 48.745 37.580 ;
        RECT  44.955 33.080 45.445 40.230 ;
        RECT  39.285 33.080 44.955 37.580 ;
        RECT  41.875 39.450 42.365 44.475 ;
        RECT  38.880 40.975 41.875 44.475 ;
        RECT  38.880 33.080 39.285 40.230 ;
        RECT  38.795 1.250 38.880 40.230 ;
        RECT  36.205 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  36.120 1.250 38.795 37.580 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  36.120 39.450 36.205 75.975 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  33.125 33.080 36.120 37.580 ;
        RECT  35.715 39.450 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  30.045 40.975 35.715 44.475 ;
        RECT  32.635 33.080 33.125 40.230 ;
        RECT  25.735 33.080 32.635 37.580 ;
        RECT  29.555 39.450 30.045 44.475 ;
        RECT  23.605 40.975 29.555 44.475 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  25.565 33.080 25.735 40.710 ;
        RECT  24.085 33.080 25.565 37.580 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA4 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA5 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 50.000 120.000 ;
        LAYER VIA6 ;
        RECT  38.880 1.250 50.000 4.750 ;
        RECT  38.880 5.750 50.000 9.250 ;
        RECT  38.880 10.250 50.000 13.750 ;
        RECT  38.880 14.750 50.000 18.250 ;
        RECT  38.880 19.250 50.000 22.750 ;
        RECT  38.880 23.750 50.000 27.250 ;
        RECT  38.880 28.250 50.000 31.750 ;
        RECT  38.880 33.080 50.000 37.580 ;
        RECT  38.880 40.975 50.000 44.475 ;
        RECT  38.880 45.475 50.000 48.975 ;
        RECT  38.880 49.975 50.000 53.475 ;
        RECT  38.880 54.475 50.000 57.975 ;
        RECT  38.880 58.975 50.000 62.475 ;
        RECT  38.880 63.475 50.000 66.975 ;
        RECT  38.880 67.975 50.000 71.475 ;
        RECT  38.880 72.475 50.000 75.975 ;
        RECT  0.000 79.975 50.000 82.975 ;
        RECT  38.880 83.670 50.000 87.170 ;
        RECT  38.880 88.020 50.000 91.520 ;
        RECT  38.880 92.370 50.000 95.870 ;
        RECT  38.880 96.720 50.000 100.220 ;
        RECT  38.880 101.070 50.000 104.570 ;
        RECT  38.880 105.420 50.000 108.920 ;
        RECT  38.880 109.770 50.000 113.270 ;
        RECT  38.880 114.010 50.000 117.510 ;
        RECT  36.120 1.250 38.880 37.580 ;
        RECT  36.120 40.975 38.880 75.975 ;
        RECT  36.120 83.670 38.880 117.510 ;
        RECT  34.665 119.000 37.555 120.000 ;
        RECT  13.880 1.250 36.120 4.750 ;
        RECT  13.880 5.750 36.120 9.250 ;
        RECT  13.880 10.250 36.120 13.750 ;
        RECT  13.880 14.750 36.120 18.250 ;
        RECT  13.880 19.250 36.120 22.750 ;
        RECT  13.880 23.750 36.120 27.250 ;
        RECT  13.880 28.250 36.120 31.750 ;
        RECT  13.880 33.080 36.120 37.580 ;
        RECT  13.880 40.975 36.120 44.475 ;
        RECT  13.880 45.475 36.120 48.975 ;
        RECT  13.880 49.975 36.120 53.475 ;
        RECT  13.880 54.475 36.120 57.975 ;
        RECT  13.880 58.975 36.120 62.475 ;
        RECT  13.880 63.475 36.120 66.975 ;
        RECT  13.880 67.975 36.120 71.475 ;
        RECT  13.880 72.475 36.120 75.975 ;
        RECT  13.880 83.670 36.120 87.170 ;
        RECT  13.880 88.020 36.120 91.520 ;
        RECT  13.880 92.370 36.120 95.870 ;
        RECT  13.880 96.720 36.120 100.220 ;
        RECT  13.880 101.070 36.120 104.570 ;
        RECT  13.880 105.420 36.120 108.920 ;
        RECT  13.880 109.770 36.120 113.270 ;
        RECT  13.880 114.010 36.120 117.510 ;
        RECT  26.525 119.000 29.415 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 50.000 120.000 ;
    END
END PDXOE3DG_G

MACRO PENDCAPA_G
    CLASS PAD ;
    FOREIGN PENDCAPA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.500 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M5 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M6 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M7 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M4 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M5 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M6 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M7 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M4 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M5 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M6 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M7 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M3 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M4 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M5 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M6 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M7 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M3 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M4 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M5 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M6 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M7 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M3 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M4 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M5 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M6 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M7 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M3 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M4 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M5 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M6 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M7 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M6 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M5 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M4 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M3 ;
        RECT  0.000 105.420 12.500 108.920 ;
        END
    END VSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M3 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M4 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M5 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M6 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 40.975 5.760 44.475 ;
        RECT  0.000 45.475 5.760 48.975 ;
        RECT  0.000 49.975 5.760 53.475 ;
        RECT  0.000 54.475 5.760 57.975 ;
        RECT  0.000 58.975 5.760 62.475 ;
        RECT  0.000 63.475 5.760 66.975 ;
        RECT  0.000 67.975 5.760 71.475 ;
        RECT  0.000 72.475 5.760 75.975 ;
        RECT  0.000 79.975 5.760 82.975 ;
        LAYER M7 ;
        RECT  0.000 0.000 12.500 120.000 ;
    END
END PENDCAPA_G

MACRO PENDCAP_G
    CLASS PAD ;
    FOREIGN PENDCAP_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.500 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        LAYER M6 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        LAYER M5 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        LAYER M4 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        LAYER M3 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M5 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M6 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M7 ;
        RECT  0.000 109.770 12.500 113.270 ;
        LAYER M4 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M5 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M6 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M7 ;
        RECT  0.000 114.010 12.500 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M4 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M5 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M6 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M7 ;
        RECT  0.000 83.670 12.500 87.170 ;
        LAYER M3 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M4 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M5 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M6 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M7 ;
        RECT  0.000 88.020 12.500 91.520 ;
        LAYER M3 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M4 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M5 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M6 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M7 ;
        RECT  0.000 92.370 12.500 95.870 ;
        LAYER M3 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M4 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M5 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M6 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M7 ;
        RECT  0.000 96.720 12.500 100.220 ;
        LAYER M3 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M4 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M5 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M6 ;
        RECT  0.000 101.070 12.500 104.570 ;
        LAYER M7 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M6 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M5 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M4 ;
        RECT  0.000 105.420 12.500 108.920 ;
        LAYER M3 ;
        RECT  0.000 105.420 12.500 108.920 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 109.770 7.500 113.270 ;
        RECT  0.000 114.010 7.500 117.510 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 7.500 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M3 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M4 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M5 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M6 ;
        RECT  0.000 0.000 12.500 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 83.670 12.500 87.170 ;
        RECT  0.000 88.020 12.500 91.520 ;
        RECT  0.000 92.370 12.500 95.870 ;
        RECT  0.000 96.720 12.500 100.220 ;
        RECT  0.000 101.070 12.500 104.570 ;
        RECT  0.000 105.420 12.500 108.920 ;
        RECT  0.000 109.770 12.500 113.270 ;
        RECT  0.000 114.010 12.500 117.510 ;
        RECT  0.000 1.250 7.500 4.750 ;
        RECT  0.000 5.750 7.500 9.250 ;
        RECT  0.000 10.250 7.500 13.750 ;
        RECT  0.000 14.750 7.500 18.250 ;
        RECT  0.000 19.250 7.500 22.750 ;
        RECT  0.000 23.750 7.500 27.250 ;
        RECT  0.000 28.250 7.500 31.750 ;
        RECT  0.000 33.080 7.500 37.580 ;
        RECT  0.000 40.975 7.500 44.475 ;
        RECT  0.000 45.475 7.500 48.975 ;
        RECT  0.000 49.975 7.500 53.475 ;
        RECT  0.000 54.475 7.500 57.975 ;
        RECT  0.000 58.975 7.500 62.475 ;
        RECT  0.000 63.475 7.500 66.975 ;
        RECT  0.000 67.975 7.500 71.475 ;
        RECT  0.000 72.475 7.500 75.975 ;
        RECT  0.000 79.975 7.500 82.975 ;
        LAYER M7 ;
        RECT  0.000 0.000 12.500 120.000 ;
    END
END PENDCAP_G

MACRO PFILLER0005A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER0005A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.005 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 0.005 5.750 ;
        RECT  0.000 7.250 0.005 11.750 ;
        RECT  0.000 13.250 0.005 17.750 ;
        RECT  0.000 19.250 0.005 23.750 ;
        RECT  0.000 25.250 0.005 29.750 ;
        RECT  0.000 31.250 0.005 35.750 ;
        RECT  0.000 36.750 0.005 39.290 ;
        LAYER M6 ;
        RECT  0.000 1.250 0.005 5.750 ;
        RECT  0.000 7.250 0.005 11.750 ;
        RECT  0.000 13.250 0.005 17.750 ;
        RECT  0.000 19.250 0.005 23.750 ;
        RECT  0.000 25.250 0.005 29.750 ;
        RECT  0.000 31.250 0.005 35.750 ;
        RECT  0.000 36.750 0.005 39.290 ;
        LAYER M5 ;
        RECT  0.000 1.250 0.005 5.750 ;
        RECT  0.000 7.250 0.005 11.750 ;
        RECT  0.000 13.250 0.005 17.750 ;
        RECT  0.000 19.250 0.005 23.750 ;
        RECT  0.000 25.250 0.005 29.750 ;
        RECT  0.000 31.250 0.005 35.750 ;
        RECT  0.000 36.750 0.005 39.290 ;
        LAYER M4 ;
        RECT  0.000 1.250 0.005 5.750 ;
        RECT  0.000 7.250 0.005 11.750 ;
        RECT  0.000 13.250 0.005 17.750 ;
        RECT  0.000 19.250 0.005 23.750 ;
        RECT  0.000 25.250 0.005 29.750 ;
        RECT  0.000 31.250 0.005 35.750 ;
        RECT  0.000 36.750 0.005 39.290 ;
        LAYER M3 ;
        RECT  0.000 1.250 0.005 5.750 ;
        RECT  0.000 7.250 0.005 11.750 ;
        RECT  0.000 13.250 0.005 17.750 ;
        RECT  0.000 19.250 0.005 23.750 ;
        RECT  0.000 25.250 0.005 29.750 ;
        RECT  0.000 31.250 0.005 35.750 ;
        RECT  0.000 36.750 0.005 39.290 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.005 120.000 ;
    END
END PFILLER0005A_G

MACRO PFILLER0005_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER0005_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.005 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 0.005 4.750 ;
        RECT  0.000 5.750 0.005 9.250 ;
        RECT  0.000 10.250 0.005 13.750 ;
        RECT  0.000 14.750 0.005 18.250 ;
        RECT  0.000 19.250 0.005 22.750 ;
        RECT  0.000 23.750 0.005 27.250 ;
        RECT  0.000 28.250 0.005 31.750 ;
        RECT  0.000 33.080 0.005 37.580 ;
        LAYER M6 ;
        RECT  0.000 1.250 0.005 4.750 ;
        RECT  0.000 5.750 0.005 9.250 ;
        RECT  0.000 10.250 0.005 13.750 ;
        RECT  0.000 14.750 0.005 18.250 ;
        RECT  0.000 19.250 0.005 22.750 ;
        RECT  0.000 23.750 0.005 27.250 ;
        RECT  0.000 28.250 0.005 31.750 ;
        RECT  0.000 33.080 0.005 37.580 ;
        LAYER M5 ;
        RECT  0.000 1.250 0.005 4.750 ;
        RECT  0.000 5.750 0.005 9.250 ;
        RECT  0.000 10.250 0.005 13.750 ;
        RECT  0.000 14.750 0.005 18.250 ;
        RECT  0.000 19.250 0.005 22.750 ;
        RECT  0.000 23.750 0.005 27.250 ;
        RECT  0.000 28.250 0.005 31.750 ;
        RECT  0.000 33.080 0.005 37.580 ;
        LAYER M4 ;
        RECT  0.000 1.250 0.005 4.750 ;
        RECT  0.000 5.750 0.005 9.250 ;
        RECT  0.000 10.250 0.005 13.750 ;
        RECT  0.000 14.750 0.005 18.250 ;
        RECT  0.000 19.250 0.005 22.750 ;
        RECT  0.000 23.750 0.005 27.250 ;
        RECT  0.000 28.250 0.005 31.750 ;
        RECT  0.000 33.080 0.005 37.580 ;
        LAYER M3 ;
        RECT  0.000 1.250 0.005 4.750 ;
        RECT  0.000 5.750 0.005 9.250 ;
        RECT  0.000 10.250 0.005 13.750 ;
        RECT  0.000 14.750 0.005 18.250 ;
        RECT  0.000 19.250 0.005 22.750 ;
        RECT  0.000 23.750 0.005 27.250 ;
        RECT  0.000 28.250 0.005 31.750 ;
        RECT  0.000 33.080 0.005 37.580 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 0.005 87.170 ;
        RECT  0.000 88.020 0.005 91.520 ;
        RECT  0.000 92.370 0.005 95.870 ;
        RECT  0.000 96.720 0.005 100.220 ;
        RECT  0.000 101.070 0.005 104.570 ;
        RECT  0.000 105.420 0.005 108.920 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 0.005 44.475 ;
        RECT  0.000 45.475 0.005 48.975 ;
        RECT  0.000 49.975 0.005 53.475 ;
        RECT  0.000 54.475 0.005 57.975 ;
        RECT  0.000 58.975 0.005 62.475 ;
        RECT  0.000 63.475 0.005 66.975 ;
        RECT  0.000 67.975 0.005 71.475 ;
        RECT  0.000 72.475 0.005 75.975 ;
        RECT  0.000 79.975 0.005 82.975 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 109.770 0.005 113.270 ;
        RECT  0.000 114.010 0.005 117.510 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 0.005 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.005 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.005 120.000 ;
    END
END PFILLER0005_G

MACRO PFILLER05A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER05A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.500 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 0.500 5.750 ;
        RECT  0.000 7.250 0.500 11.750 ;
        RECT  0.000 13.250 0.500 17.750 ;
        RECT  0.000 19.250 0.500 23.750 ;
        RECT  0.000 25.250 0.500 29.750 ;
        RECT  0.000 31.250 0.500 35.750 ;
        RECT  0.000 36.750 0.500 39.290 ;
        LAYER M6 ;
        RECT  0.000 1.250 0.500 5.750 ;
        RECT  0.000 7.250 0.500 11.750 ;
        RECT  0.000 13.250 0.500 17.750 ;
        RECT  0.000 19.250 0.500 23.750 ;
        RECT  0.000 25.250 0.500 29.750 ;
        RECT  0.000 31.250 0.500 35.750 ;
        RECT  0.000 36.750 0.500 39.290 ;
        LAYER M5 ;
        RECT  0.000 1.250 0.500 5.750 ;
        RECT  0.000 7.250 0.500 11.750 ;
        RECT  0.000 13.250 0.500 17.750 ;
        RECT  0.000 19.250 0.500 23.750 ;
        RECT  0.000 25.250 0.500 29.750 ;
        RECT  0.000 31.250 0.500 35.750 ;
        RECT  0.000 36.750 0.500 39.290 ;
        LAYER M4 ;
        RECT  0.000 1.250 0.500 5.750 ;
        RECT  0.000 7.250 0.500 11.750 ;
        RECT  0.000 13.250 0.500 17.750 ;
        RECT  0.000 19.250 0.500 23.750 ;
        RECT  0.000 25.250 0.500 29.750 ;
        RECT  0.000 31.250 0.500 35.750 ;
        RECT  0.000 36.750 0.500 39.290 ;
        LAYER M3 ;
        RECT  0.000 1.250 0.500 5.750 ;
        RECT  0.000 7.250 0.500 11.750 ;
        RECT  0.000 13.250 0.500 17.750 ;
        RECT  0.000 19.250 0.500 23.750 ;
        RECT  0.000 25.250 0.500 29.750 ;
        RECT  0.000 31.250 0.500 35.750 ;
        RECT  0.000 36.750 0.500 39.290 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.500 120.000 ;
    END
END PFILLER05A_G

MACRO PFILLER05_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER05_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.500 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 0.500 4.750 ;
        RECT  0.000 5.750 0.500 9.250 ;
        RECT  0.000 10.250 0.500 13.750 ;
        RECT  0.000 14.750 0.500 18.250 ;
        RECT  0.000 19.250 0.500 22.750 ;
        RECT  0.000 23.750 0.500 27.250 ;
        RECT  0.000 28.250 0.500 31.750 ;
        RECT  0.000 33.080 0.500 37.580 ;
        LAYER M6 ;
        RECT  0.000 1.250 0.500 4.750 ;
        RECT  0.000 5.750 0.500 9.250 ;
        RECT  0.000 10.250 0.500 13.750 ;
        RECT  0.000 14.750 0.500 18.250 ;
        RECT  0.000 19.250 0.500 22.750 ;
        RECT  0.000 23.750 0.500 27.250 ;
        RECT  0.000 28.250 0.500 31.750 ;
        RECT  0.000 33.080 0.500 37.580 ;
        LAYER M5 ;
        RECT  0.000 1.250 0.500 4.750 ;
        RECT  0.000 5.750 0.500 9.250 ;
        RECT  0.000 10.250 0.500 13.750 ;
        RECT  0.000 14.750 0.500 18.250 ;
        RECT  0.000 19.250 0.500 22.750 ;
        RECT  0.000 23.750 0.500 27.250 ;
        RECT  0.000 28.250 0.500 31.750 ;
        RECT  0.000 33.080 0.500 37.580 ;
        LAYER M4 ;
        RECT  0.000 1.250 0.500 4.750 ;
        RECT  0.000 5.750 0.500 9.250 ;
        RECT  0.000 10.250 0.500 13.750 ;
        RECT  0.000 14.750 0.500 18.250 ;
        RECT  0.000 19.250 0.500 22.750 ;
        RECT  0.000 23.750 0.500 27.250 ;
        RECT  0.000 28.250 0.500 31.750 ;
        RECT  0.000 33.080 0.500 37.580 ;
        LAYER M3 ;
        RECT  0.000 1.250 0.500 4.750 ;
        RECT  0.000 5.750 0.500 9.250 ;
        RECT  0.000 10.250 0.500 13.750 ;
        RECT  0.000 14.750 0.500 18.250 ;
        RECT  0.000 19.250 0.500 22.750 ;
        RECT  0.000 23.750 0.500 27.250 ;
        RECT  0.000 28.250 0.500 31.750 ;
        RECT  0.000 33.080 0.500 37.580 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 0.500 87.170 ;
        RECT  0.000 88.020 0.500 91.520 ;
        RECT  0.000 92.370 0.500 95.870 ;
        RECT  0.000 96.720 0.500 100.220 ;
        RECT  0.000 101.070 0.500 104.570 ;
        RECT  0.000 105.420 0.500 108.920 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 0.500 44.475 ;
        RECT  0.000 45.475 0.500 48.975 ;
        RECT  0.000 49.975 0.500 53.475 ;
        RECT  0.000 54.475 0.500 57.975 ;
        RECT  0.000 58.975 0.500 62.475 ;
        RECT  0.000 63.475 0.500 66.975 ;
        RECT  0.000 67.975 0.500 71.475 ;
        RECT  0.000 72.475 0.500 75.975 ;
        RECT  0.000 79.975 0.500 82.975 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 109.770 0.500 113.270 ;
        RECT  0.000 114.010 0.500 117.510 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 0.500 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 0.500 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 0.500 120.000 ;
    END
END PFILLER05_G

MACRO PFILLER10A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER10A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 6.380 87.170 6.380 88.020
                 10.000 88.020 10.000 91.520 6.380 91.520 6.380 92.370 10.000 92.370
                 10.000 95.870 6.380 95.870 6.380 96.720 10.000 96.720 10.000 100.220
                 6.380 100.220 6.380 101.070 10.000 101.070 10.000 104.570 6.380 104.570
                 6.380 105.420 10.000 105.420 10.000 108.920 6.380 108.920 6.380 109.770
                 10.000 109.770 10.000 113.270 6.380 113.270 6.380 114.010 10.000 114.010
                 10.000 117.510 0.000 117.510 0.000 114.010 3.620 114.010 3.620 113.270
                 0.000 113.270 0.000 109.770 3.620 109.770 3.620 108.920 0.000 108.920
                 0.000 105.420 3.620 105.420 3.620 104.570 0.000 104.570 0.000 101.070
                 3.620 101.070 3.620 100.220 0.000 100.220 0.000 96.720 3.620 96.720
                 3.620 95.870 0.000 95.870 0.000 92.370 3.620 92.370 3.620 91.520
                 0.000 91.520 0.000 88.020 3.620 88.020 3.620 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 6.380 87.170 6.380 88.020
                 10.000 88.020 10.000 91.520 6.380 91.520 6.380 92.370 10.000 92.370
                 10.000 95.870 6.380 95.870 6.380 96.720 10.000 96.720 10.000 100.220
                 6.380 100.220 6.380 101.070 10.000 101.070 10.000 104.570 6.380 104.570
                 6.380 105.420 10.000 105.420 10.000 108.920 6.380 108.920 6.380 109.770
                 10.000 109.770 10.000 113.270 6.380 113.270 6.380 114.010 10.000 114.010
                 10.000 117.510 0.000 117.510 0.000 114.010 3.620 114.010 3.620 113.270
                 0.000 113.270 0.000 109.770 3.620 109.770 3.620 108.920 0.000 108.920
                 0.000 105.420 3.620 105.420 3.620 104.570 0.000 104.570 0.000 101.070
                 3.620 101.070 3.620 100.220 0.000 100.220 0.000 96.720 3.620 96.720
                 3.620 95.870 0.000 95.870 0.000 92.370 3.620 92.370 3.620 91.520
                 0.000 91.520 0.000 88.020 3.620 88.020 3.620 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 6.380 87.170 6.380 88.020
                 10.000 88.020 10.000 91.520 6.380 91.520 6.380 92.370 10.000 92.370
                 10.000 95.870 6.380 95.870 6.380 96.720 10.000 96.720 10.000 100.220
                 6.380 100.220 6.380 101.070 10.000 101.070 10.000 104.570 6.380 104.570
                 6.380 105.420 10.000 105.420 10.000 108.920 6.380 108.920 6.380 109.770
                 10.000 109.770 10.000 113.270 6.380 113.270 6.380 114.010 10.000 114.010
                 10.000 117.510 0.000 117.510 0.000 114.010 3.620 114.010 3.620 113.270
                 0.000 113.270 0.000 109.770 3.620 109.770 3.620 108.920 0.000 108.920
                 0.000 105.420 3.620 105.420 3.620 104.570 0.000 104.570 0.000 101.070
                 3.620 101.070 3.620 100.220 0.000 100.220 0.000 96.720 3.620 96.720
                 3.620 95.870 0.000 95.870 0.000 92.370 3.620 92.370 3.620 91.520
                 0.000 91.520 0.000 88.020 3.620 88.020 3.620 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 6.380 87.170 6.380 88.020
                 10.000 88.020 10.000 91.520 6.380 91.520 6.380 92.370 10.000 92.370
                 10.000 95.870 6.380 95.870 6.380 96.720 10.000 96.720 10.000 100.220
                 6.380 100.220 6.380 101.070 10.000 101.070 10.000 104.570 6.380 104.570
                 6.380 105.420 10.000 105.420 10.000 108.920 6.380 108.920 6.380 109.770
                 10.000 109.770 10.000 113.270 6.380 113.270 6.380 114.010 10.000 114.010
                 10.000 117.510 0.000 117.510 0.000 114.010 3.620 114.010 3.620 113.270
                 0.000 113.270 0.000 109.770 3.620 109.770 3.620 108.920 0.000 108.920
                 0.000 105.420 3.620 105.420 3.620 104.570 0.000 104.570 0.000 101.070
                 3.620 101.070 3.620 100.220 0.000 100.220 0.000 96.720 3.620 96.720
                 3.620 95.870 0.000 95.870 0.000 92.370 3.620 92.370 3.620 91.520
                 0.000 91.520 0.000 88.020 3.620 88.020 3.620 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 6.380 87.170 6.380 88.020
                 10.000 88.020 10.000 91.520 6.380 91.520 6.380 92.370 10.000 92.370
                 10.000 95.870 6.380 95.870 6.380 96.720 10.000 96.720 10.000 100.220
                 6.380 100.220 6.380 101.070 10.000 101.070 10.000 104.570 6.380 104.570
                 6.380 105.420 10.000 105.420 10.000 108.920 6.380 108.920 6.380 109.770
                 10.000 109.770 10.000 113.270 6.380 113.270 6.380 114.010 10.000 114.010
                 10.000 117.510 0.000 117.510 0.000 114.010 3.620 114.010 3.620 113.270
                 0.000 113.270 0.000 109.770 3.620 109.770 3.620 108.920 0.000 108.920
                 0.000 105.420 3.620 105.420 3.620 104.570 0.000 104.570 0.000 101.070
                 3.620 101.070 3.620 100.220 0.000 100.220 0.000 96.720 3.620 96.720
                 3.620 95.870 0.000 95.870 0.000 92.370 3.620 92.370 3.620 91.520
                 0.000 91.520 0.000 88.020 3.620 88.020 3.620 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 5.750 6.380 5.750 6.380 7.250 10.000 7.250
                 10.000 11.750 6.380 11.750 6.380 13.250 10.000 13.250 10.000 17.750
                 6.380 17.750 6.380 19.250 10.000 19.250 10.000 23.750 6.380 23.750
                 6.380 25.250 10.000 25.250 10.000 29.750 6.380 29.750 6.380 31.250
                 10.000 31.250 10.000 35.750 6.380 35.750 6.380 36.750 10.000 36.750
                 10.000 39.290 0.000 39.290 0.000 36.750 3.620 36.750 3.620 35.750
                 0.000 35.750 0.000 31.250 3.620 31.250 3.620 29.750 0.000 29.750
                 0.000 25.250 3.620 25.250 3.620 23.750 0.000 23.750 0.000 19.250
                 3.620 19.250 3.620 17.750 0.000 17.750 0.000 13.250 3.620 13.250
                 3.620 11.750 0.000 11.750 0.000 7.250 3.620 7.250 3.620 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 5.750 6.380 5.750 6.380 7.250 10.000 7.250
                 10.000 11.750 6.380 11.750 6.380 13.250 10.000 13.250 10.000 17.750
                 6.380 17.750 6.380 19.250 10.000 19.250 10.000 23.750 6.380 23.750
                 6.380 25.250 10.000 25.250 10.000 29.750 6.380 29.750 6.380 31.250
                 10.000 31.250 10.000 35.750 6.380 35.750 6.380 36.750 10.000 36.750
                 10.000 39.290 0.000 39.290 0.000 36.750 3.620 36.750 3.620 35.750
                 0.000 35.750 0.000 31.250 3.620 31.250 3.620 29.750 0.000 29.750
                 0.000 25.250 3.620 25.250 3.620 23.750 0.000 23.750 0.000 19.250
                 3.620 19.250 3.620 17.750 0.000 17.750 0.000 13.250 3.620 13.250
                 3.620 11.750 0.000 11.750 0.000 7.250 3.620 7.250 3.620 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 5.750 6.380 5.750 6.380 7.250 10.000 7.250
                 10.000 11.750 6.380 11.750 6.380 13.250 10.000 13.250 10.000 17.750
                 6.380 17.750 6.380 19.250 10.000 19.250 10.000 23.750 6.380 23.750
                 6.380 25.250 10.000 25.250 10.000 29.750 6.380 29.750 6.380 31.250
                 10.000 31.250 10.000 35.750 6.380 35.750 6.380 36.750 10.000 36.750
                 10.000 39.290 0.000 39.290 0.000 36.750 3.620 36.750 3.620 35.750
                 0.000 35.750 0.000 31.250 3.620 31.250 3.620 29.750 0.000 29.750
                 0.000 25.250 3.620 25.250 3.620 23.750 0.000 23.750 0.000 19.250
                 3.620 19.250 3.620 17.750 0.000 17.750 0.000 13.250 3.620 13.250
                 3.620 11.750 0.000 11.750 0.000 7.250 3.620 7.250 3.620 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 5.750 6.380 5.750 6.380 7.250 10.000 7.250
                 10.000 11.750 6.380 11.750 6.380 13.250 10.000 13.250 10.000 17.750
                 6.380 17.750 6.380 19.250 10.000 19.250 10.000 23.750 6.380 23.750
                 6.380 25.250 10.000 25.250 10.000 29.750 6.380 29.750 6.380 31.250
                 10.000 31.250 10.000 35.750 6.380 35.750 6.380 36.750 10.000 36.750
                 10.000 39.290 0.000 39.290 0.000 36.750 3.620 36.750 3.620 35.750
                 0.000 35.750 0.000 31.250 3.620 31.250 3.620 29.750 0.000 29.750
                 0.000 25.250 3.620 25.250 3.620 23.750 0.000 23.750 0.000 19.250
                 3.620 19.250 3.620 17.750 0.000 17.750 0.000 13.250 3.620 13.250
                 3.620 11.750 0.000 11.750 0.000 7.250 3.620 7.250 3.620 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 5.750 6.380 5.750 6.380 7.250 10.000 7.250
                 10.000 11.750 6.380 11.750 6.380 13.250 10.000 13.250 10.000 17.750
                 6.380 17.750 6.380 19.250 10.000 19.250 10.000 23.750 6.380 23.750
                 6.380 25.250 10.000 25.250 10.000 29.750 6.380 29.750 6.380 31.250
                 10.000 31.250 10.000 35.750 6.380 35.750 6.380 36.750 10.000 36.750
                 10.000 39.290 0.000 39.290 0.000 36.750 3.620 36.750 3.620 35.750
                 0.000 35.750 0.000 31.250 3.620 31.250 3.620 29.750 0.000 29.750
                 0.000 25.250 3.620 25.250 3.620 23.750 0.000 23.750 0.000 19.250
                 3.620 19.250 3.620 17.750 0.000 17.750 0.000 13.250 3.620 13.250
                 3.620 11.750 0.000 11.750 0.000 7.250 3.620 7.250 3.620 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 6.380 44.475 6.380 45.475
                 10.000 45.475 10.000 48.975 6.380 48.975 6.380 49.975 10.000 49.975
                 10.000 53.475 6.380 53.475 6.380 54.475 10.000 54.475 10.000 57.975
                 6.380 57.975 6.380 58.975 10.000 58.975 10.000 62.475 6.380 62.475
                 6.380 63.475 10.000 63.475 10.000 66.975 6.380 66.975 6.380 67.975
                 10.000 67.975 10.000 71.475 6.380 71.475 6.380 72.475 10.000 72.475
                 10.000 75.975 0.000 75.975 0.000 72.475 3.620 72.475 3.620 71.475
                 0.000 71.475 0.000 67.975 3.620 67.975 3.620 66.975 0.000 66.975
                 0.000 63.475 3.620 63.475 3.620 62.475 0.000 62.475 0.000 58.975
                 3.620 58.975 3.620 57.975 0.000 57.975 0.000 54.475 3.620 54.475
                 3.620 53.475 0.000 53.475 0.000 49.975 3.620 49.975 3.620 48.975
                 0.000 48.975 0.000 45.475 3.620 45.475 3.620 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 6.380 44.475 6.380 45.475
                 10.000 45.475 10.000 48.975 6.380 48.975 6.380 49.975 10.000 49.975
                 10.000 53.475 6.380 53.475 6.380 54.475 10.000 54.475 10.000 57.975
                 6.380 57.975 6.380 58.975 10.000 58.975 10.000 62.475 6.380 62.475
                 6.380 63.475 10.000 63.475 10.000 66.975 6.380 66.975 6.380 67.975
                 10.000 67.975 10.000 71.475 6.380 71.475 6.380 72.475 10.000 72.475
                 10.000 75.975 0.000 75.975 0.000 72.475 3.620 72.475 3.620 71.475
                 0.000 71.475 0.000 67.975 3.620 67.975 3.620 66.975 0.000 66.975
                 0.000 63.475 3.620 63.475 3.620 62.475 0.000 62.475 0.000 58.975
                 3.620 58.975 3.620 57.975 0.000 57.975 0.000 54.475 3.620 54.475
                 3.620 53.475 0.000 53.475 0.000 49.975 3.620 49.975 3.620 48.975
                 0.000 48.975 0.000 45.475 3.620 45.475 3.620 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 6.380 44.475 6.380 45.475
                 10.000 45.475 10.000 48.975 6.380 48.975 6.380 49.975 10.000 49.975
                 10.000 53.475 6.380 53.475 6.380 54.475 10.000 54.475 10.000 57.975
                 6.380 57.975 6.380 58.975 10.000 58.975 10.000 62.475 6.380 62.475
                 6.380 63.475 10.000 63.475 10.000 66.975 6.380 66.975 6.380 67.975
                 10.000 67.975 10.000 71.475 6.380 71.475 6.380 72.475 10.000 72.475
                 10.000 75.975 0.000 75.975 0.000 72.475 3.620 72.475 3.620 71.475
                 0.000 71.475 0.000 67.975 3.620 67.975 3.620 66.975 0.000 66.975
                 0.000 63.475 3.620 63.475 3.620 62.475 0.000 62.475 0.000 58.975
                 3.620 58.975 3.620 57.975 0.000 57.975 0.000 54.475 3.620 54.475
                 3.620 53.475 0.000 53.475 0.000 49.975 3.620 49.975 3.620 48.975
                 0.000 48.975 0.000 45.475 3.620 45.475 3.620 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 6.380 44.475 6.380 45.475
                 10.000 45.475 10.000 48.975 6.380 48.975 6.380 49.975 10.000 49.975
                 10.000 53.475 6.380 53.475 6.380 54.475 10.000 54.475 10.000 57.975
                 6.380 57.975 6.380 58.975 10.000 58.975 10.000 62.475 6.380 62.475
                 6.380 63.475 10.000 63.475 10.000 66.975 6.380 66.975 6.380 67.975
                 10.000 67.975 10.000 71.475 6.380 71.475 6.380 72.475 10.000 72.475
                 10.000 75.975 0.000 75.975 0.000 72.475 3.620 72.475 3.620 71.475
                 0.000 71.475 0.000 67.975 3.620 67.975 3.620 66.975 0.000 66.975
                 0.000 63.475 3.620 63.475 3.620 62.475 0.000 62.475 0.000 58.975
                 3.620 58.975 3.620 57.975 0.000 57.975 0.000 54.475 3.620 54.475
                 3.620 53.475 0.000 53.475 0.000 49.975 3.620 49.975 3.620 48.975
                 0.000 48.975 0.000 45.475 3.620 45.475 3.620 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 6.380 44.475 6.380 45.475
                 10.000 45.475 10.000 48.975 6.380 48.975 6.380 49.975 10.000 49.975
                 10.000 53.475 6.380 53.475 6.380 54.475 10.000 54.475 10.000 57.975
                 6.380 57.975 6.380 58.975 10.000 58.975 10.000 62.475 6.380 62.475
                 6.380 63.475 10.000 63.475 10.000 66.975 6.380 66.975 6.380 67.975
                 10.000 67.975 10.000 71.475 6.380 71.475 6.380 72.475 10.000 72.475
                 10.000 75.975 0.000 75.975 0.000 72.475 3.620 72.475 3.620 71.475
                 0.000 71.475 0.000 67.975 3.620 67.975 3.620 66.975 0.000 66.975
                 0.000 63.475 3.620 63.475 3.620 62.475 0.000 62.475 0.000 58.975
                 3.620 58.975 3.620 57.975 0.000 57.975 0.000 54.475 3.620 54.475
                 3.620 53.475 0.000 53.475 0.000 49.975 3.620 49.975 3.620 48.975
                 0.000 48.975 0.000 45.475 3.620 45.475 3.620 44.475 0.000 44.475 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA2 ;
        RECT  6.380 1.250 10.000 5.750 ;
        RECT  6.380 7.250 10.000 11.750 ;
        RECT  6.380 13.250 10.000 17.750 ;
        RECT  6.380 19.250 10.000 23.750 ;
        RECT  6.380 25.250 10.000 29.750 ;
        RECT  6.380 31.250 10.000 35.750 ;
        RECT  6.380 36.750 10.000 39.290 ;
        RECT  6.380 40.975 10.000 44.475 ;
        RECT  6.380 45.475 10.000 48.975 ;
        RECT  6.380 49.975 10.000 53.475 ;
        RECT  6.380 54.475 10.000 57.975 ;
        RECT  6.380 58.975 10.000 62.475 ;
        RECT  6.380 63.475 10.000 66.975 ;
        RECT  6.380 67.975 10.000 71.475 ;
        RECT  6.380 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  6.380 83.670 10.000 87.170 ;
        RECT  6.380 88.020 10.000 91.520 ;
        RECT  6.380 92.370 10.000 95.870 ;
        RECT  6.380 96.720 10.000 100.220 ;
        RECT  6.380 101.070 10.000 104.570 ;
        RECT  6.380 105.420 10.000 108.920 ;
        RECT  6.380 109.770 10.000 113.270 ;
        RECT  6.380 114.010 10.000 117.510 ;
        RECT  3.620 1.250 6.380 39.290 ;
        RECT  3.620 40.975 6.380 75.975 ;
        RECT  3.620 83.670 6.380 117.510 ;
        RECT  0.000 1.250 3.620 5.750 ;
        RECT  0.000 7.250 3.620 11.750 ;
        RECT  0.000 13.250 3.620 17.750 ;
        RECT  0.000 19.250 3.620 23.750 ;
        RECT  0.000 25.250 3.620 29.750 ;
        RECT  0.000 31.250 3.620 35.750 ;
        RECT  0.000 36.750 3.620 39.290 ;
        RECT  0.000 40.975 3.620 44.475 ;
        RECT  0.000 45.475 3.620 48.975 ;
        RECT  0.000 49.975 3.620 53.475 ;
        RECT  0.000 54.475 3.620 57.975 ;
        RECT  0.000 58.975 3.620 62.475 ;
        RECT  0.000 63.475 3.620 66.975 ;
        RECT  0.000 67.975 3.620 71.475 ;
        RECT  0.000 72.475 3.620 75.975 ;
        RECT  0.000 83.670 3.620 87.170 ;
        RECT  0.000 88.020 3.620 91.520 ;
        RECT  0.000 92.370 3.620 95.870 ;
        RECT  0.000 96.720 3.620 100.220 ;
        RECT  0.000 101.070 3.620 104.570 ;
        RECT  0.000 105.420 3.620 108.920 ;
        RECT  0.000 109.770 3.620 113.270 ;
        RECT  0.000 114.010 3.620 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA3 ;
        RECT  6.380 1.250 10.000 5.750 ;
        RECT  6.380 7.250 10.000 11.750 ;
        RECT  6.380 13.250 10.000 17.750 ;
        RECT  6.380 19.250 10.000 23.750 ;
        RECT  6.380 25.250 10.000 29.750 ;
        RECT  6.380 31.250 10.000 35.750 ;
        RECT  6.380 36.750 10.000 39.290 ;
        RECT  6.380 40.975 10.000 44.475 ;
        RECT  6.380 45.475 10.000 48.975 ;
        RECT  6.380 49.975 10.000 53.475 ;
        RECT  6.380 54.475 10.000 57.975 ;
        RECT  6.380 58.975 10.000 62.475 ;
        RECT  6.380 63.475 10.000 66.975 ;
        RECT  6.380 67.975 10.000 71.475 ;
        RECT  6.380 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  6.380 83.670 10.000 87.170 ;
        RECT  6.380 88.020 10.000 91.520 ;
        RECT  6.380 92.370 10.000 95.870 ;
        RECT  6.380 96.720 10.000 100.220 ;
        RECT  6.380 101.070 10.000 104.570 ;
        RECT  6.380 105.420 10.000 108.920 ;
        RECT  6.380 109.770 10.000 113.270 ;
        RECT  6.380 114.010 10.000 117.510 ;
        RECT  3.620 1.250 6.380 39.290 ;
        RECT  3.620 40.975 6.380 75.975 ;
        RECT  3.620 83.670 6.380 117.510 ;
        RECT  0.000 1.250 3.620 5.750 ;
        RECT  0.000 7.250 3.620 11.750 ;
        RECT  0.000 13.250 3.620 17.750 ;
        RECT  0.000 19.250 3.620 23.750 ;
        RECT  0.000 25.250 3.620 29.750 ;
        RECT  0.000 31.250 3.620 35.750 ;
        RECT  0.000 36.750 3.620 39.290 ;
        RECT  0.000 40.975 3.620 44.475 ;
        RECT  0.000 45.475 3.620 48.975 ;
        RECT  0.000 49.975 3.620 53.475 ;
        RECT  0.000 54.475 3.620 57.975 ;
        RECT  0.000 58.975 3.620 62.475 ;
        RECT  0.000 63.475 3.620 66.975 ;
        RECT  0.000 67.975 3.620 71.475 ;
        RECT  0.000 72.475 3.620 75.975 ;
        RECT  0.000 83.670 3.620 87.170 ;
        RECT  0.000 88.020 3.620 91.520 ;
        RECT  0.000 92.370 3.620 95.870 ;
        RECT  0.000 96.720 3.620 100.220 ;
        RECT  0.000 101.070 3.620 104.570 ;
        RECT  0.000 105.420 3.620 108.920 ;
        RECT  0.000 109.770 3.620 113.270 ;
        RECT  0.000 114.010 3.620 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA4 ;
        RECT  6.380 1.250 10.000 5.750 ;
        RECT  6.380 7.250 10.000 11.750 ;
        RECT  6.380 13.250 10.000 17.750 ;
        RECT  6.380 19.250 10.000 23.750 ;
        RECT  6.380 25.250 10.000 29.750 ;
        RECT  6.380 31.250 10.000 35.750 ;
        RECT  6.380 36.750 10.000 39.290 ;
        RECT  6.380 40.975 10.000 44.475 ;
        RECT  6.380 45.475 10.000 48.975 ;
        RECT  6.380 49.975 10.000 53.475 ;
        RECT  6.380 54.475 10.000 57.975 ;
        RECT  6.380 58.975 10.000 62.475 ;
        RECT  6.380 63.475 10.000 66.975 ;
        RECT  6.380 67.975 10.000 71.475 ;
        RECT  6.380 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  6.380 83.670 10.000 87.170 ;
        RECT  6.380 88.020 10.000 91.520 ;
        RECT  6.380 92.370 10.000 95.870 ;
        RECT  6.380 96.720 10.000 100.220 ;
        RECT  6.380 101.070 10.000 104.570 ;
        RECT  6.380 105.420 10.000 108.920 ;
        RECT  6.380 109.770 10.000 113.270 ;
        RECT  6.380 114.010 10.000 117.510 ;
        RECT  3.620 1.250 6.380 39.290 ;
        RECT  3.620 40.975 6.380 75.975 ;
        RECT  3.620 83.670 6.380 117.510 ;
        RECT  0.000 1.250 3.620 5.750 ;
        RECT  0.000 7.250 3.620 11.750 ;
        RECT  0.000 13.250 3.620 17.750 ;
        RECT  0.000 19.250 3.620 23.750 ;
        RECT  0.000 25.250 3.620 29.750 ;
        RECT  0.000 31.250 3.620 35.750 ;
        RECT  0.000 36.750 3.620 39.290 ;
        RECT  0.000 40.975 3.620 44.475 ;
        RECT  0.000 45.475 3.620 48.975 ;
        RECT  0.000 49.975 3.620 53.475 ;
        RECT  0.000 54.475 3.620 57.975 ;
        RECT  0.000 58.975 3.620 62.475 ;
        RECT  0.000 63.475 3.620 66.975 ;
        RECT  0.000 67.975 3.620 71.475 ;
        RECT  0.000 72.475 3.620 75.975 ;
        RECT  0.000 83.670 3.620 87.170 ;
        RECT  0.000 88.020 3.620 91.520 ;
        RECT  0.000 92.370 3.620 95.870 ;
        RECT  0.000 96.720 3.620 100.220 ;
        RECT  0.000 101.070 3.620 104.570 ;
        RECT  0.000 105.420 3.620 108.920 ;
        RECT  0.000 109.770 3.620 113.270 ;
        RECT  0.000 114.010 3.620 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA5 ;
        RECT  6.380 1.250 10.000 5.750 ;
        RECT  6.380 7.250 10.000 11.750 ;
        RECT  6.380 13.250 10.000 17.750 ;
        RECT  6.380 19.250 10.000 23.750 ;
        RECT  6.380 25.250 10.000 29.750 ;
        RECT  6.380 31.250 10.000 35.750 ;
        RECT  6.380 36.750 10.000 39.290 ;
        RECT  6.380 40.975 10.000 44.475 ;
        RECT  6.380 45.475 10.000 48.975 ;
        RECT  6.380 49.975 10.000 53.475 ;
        RECT  6.380 54.475 10.000 57.975 ;
        RECT  6.380 58.975 10.000 62.475 ;
        RECT  6.380 63.475 10.000 66.975 ;
        RECT  6.380 67.975 10.000 71.475 ;
        RECT  6.380 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  6.380 83.670 10.000 87.170 ;
        RECT  6.380 88.020 10.000 91.520 ;
        RECT  6.380 92.370 10.000 95.870 ;
        RECT  6.380 96.720 10.000 100.220 ;
        RECT  6.380 101.070 10.000 104.570 ;
        RECT  6.380 105.420 10.000 108.920 ;
        RECT  6.380 109.770 10.000 113.270 ;
        RECT  6.380 114.010 10.000 117.510 ;
        RECT  3.620 1.250 6.380 39.290 ;
        RECT  3.620 40.975 6.380 75.975 ;
        RECT  3.620 83.670 6.380 117.510 ;
        RECT  0.000 1.250 3.620 5.750 ;
        RECT  0.000 7.250 3.620 11.750 ;
        RECT  0.000 13.250 3.620 17.750 ;
        RECT  0.000 19.250 3.620 23.750 ;
        RECT  0.000 25.250 3.620 29.750 ;
        RECT  0.000 31.250 3.620 35.750 ;
        RECT  0.000 36.750 3.620 39.290 ;
        RECT  0.000 40.975 3.620 44.475 ;
        RECT  0.000 45.475 3.620 48.975 ;
        RECT  0.000 49.975 3.620 53.475 ;
        RECT  0.000 54.475 3.620 57.975 ;
        RECT  0.000 58.975 3.620 62.475 ;
        RECT  0.000 63.475 3.620 66.975 ;
        RECT  0.000 67.975 3.620 71.475 ;
        RECT  0.000 72.475 3.620 75.975 ;
        RECT  0.000 83.670 3.620 87.170 ;
        RECT  0.000 88.020 3.620 91.520 ;
        RECT  0.000 92.370 3.620 95.870 ;
        RECT  0.000 96.720 3.620 100.220 ;
        RECT  0.000 101.070 3.620 104.570 ;
        RECT  0.000 105.420 3.620 108.920 ;
        RECT  0.000 109.770 3.620 113.270 ;
        RECT  0.000 114.010 3.620 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA6 ;
        RECT  6.380 1.250 10.000 5.750 ;
        RECT  6.380 7.250 10.000 11.750 ;
        RECT  6.380 13.250 10.000 17.750 ;
        RECT  6.380 19.250 10.000 23.750 ;
        RECT  6.380 25.250 10.000 29.750 ;
        RECT  6.380 31.250 10.000 35.750 ;
        RECT  6.380 36.750 10.000 39.290 ;
        RECT  6.380 40.975 10.000 44.475 ;
        RECT  6.380 45.475 10.000 48.975 ;
        RECT  6.380 49.975 10.000 53.475 ;
        RECT  6.380 54.475 10.000 57.975 ;
        RECT  6.380 58.975 10.000 62.475 ;
        RECT  6.380 63.475 10.000 66.975 ;
        RECT  6.380 67.975 10.000 71.475 ;
        RECT  6.380 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  6.380 83.670 10.000 87.170 ;
        RECT  6.380 88.020 10.000 91.520 ;
        RECT  6.380 92.370 10.000 95.870 ;
        RECT  6.380 96.720 10.000 100.220 ;
        RECT  6.380 101.070 10.000 104.570 ;
        RECT  6.380 105.420 10.000 108.920 ;
        RECT  6.380 109.770 10.000 113.270 ;
        RECT  6.380 114.010 10.000 117.510 ;
        RECT  3.620 1.250 6.380 39.290 ;
        RECT  3.620 40.975 6.380 75.975 ;
        RECT  3.620 83.670 6.380 117.510 ;
        RECT  0.000 1.250 3.620 5.750 ;
        RECT  0.000 7.250 3.620 11.750 ;
        RECT  0.000 13.250 3.620 17.750 ;
        RECT  0.000 19.250 3.620 23.750 ;
        RECT  0.000 25.250 3.620 29.750 ;
        RECT  0.000 31.250 3.620 35.750 ;
        RECT  0.000 36.750 3.620 39.290 ;
        RECT  0.000 40.975 3.620 44.475 ;
        RECT  0.000 45.475 3.620 48.975 ;
        RECT  0.000 49.975 3.620 53.475 ;
        RECT  0.000 54.475 3.620 57.975 ;
        RECT  0.000 58.975 3.620 62.475 ;
        RECT  0.000 63.475 3.620 66.975 ;
        RECT  0.000 67.975 3.620 71.475 ;
        RECT  0.000 72.475 3.620 75.975 ;
        RECT  0.000 83.670 3.620 87.170 ;
        RECT  0.000 88.020 3.620 91.520 ;
        RECT  0.000 92.370 3.620 95.870 ;
        RECT  0.000 96.720 3.620 100.220 ;
        RECT  0.000 101.070 3.620 104.570 ;
        RECT  0.000 105.420 3.620 108.920 ;
        RECT  0.000 109.770 3.620 113.270 ;
        RECT  0.000 114.010 3.620 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 10.000 120.000 ;
    END
END PFILLER10A_G

MACRO PFILLER10_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER10_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 4.750 8.000 4.750 8.000 5.750 10.000 5.750
                 10.000 9.250 8.000 9.250 8.000 10.250 10.000 10.250 10.000 13.750
                 8.000 13.750 8.000 14.750 10.000 14.750 10.000 18.250 8.000 18.250
                 8.000 19.250 10.000 19.250 10.000 22.750 8.000 22.750 8.000 23.750
                 10.000 23.750 10.000 27.250 8.000 27.250 8.000 28.250 10.000 28.250
                 10.000 31.750 8.000 31.750 8.000 33.080 10.000 33.080 10.000 37.580
                 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750 7.000 9.250
                 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750 3.000 13.750
                 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250 3.000 19.250
                 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750 7.000 23.750
                 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250 7.000 31.750
                 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580 0.000 37.580
                 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750 0.000 28.250
                 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750 2.000 23.750
                 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250 2.000 18.250
                 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750 0.000 13.750
                 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750 2.000 5.750
                 2.000 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 4.750 8.000 4.750 8.000 5.750 10.000 5.750
                 10.000 9.250 8.000 9.250 8.000 10.250 10.000 10.250 10.000 13.750
                 8.000 13.750 8.000 14.750 10.000 14.750 10.000 18.250 8.000 18.250
                 8.000 19.250 10.000 19.250 10.000 22.750 8.000 22.750 8.000 23.750
                 10.000 23.750 10.000 27.250 8.000 27.250 8.000 28.250 10.000 28.250
                 10.000 31.750 8.000 31.750 8.000 33.080 10.000 33.080 10.000 37.580
                 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750 7.000 9.250
                 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750 3.000 13.750
                 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250 3.000 19.250
                 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750 7.000 23.750
                 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250 7.000 31.750
                 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580 0.000 37.580
                 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750 0.000 28.250
                 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750 2.000 23.750
                 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250 2.000 18.250
                 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750 0.000 13.750
                 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750 2.000 5.750
                 2.000 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 4.750 8.000 4.750 8.000 5.750 10.000 5.750
                 10.000 9.250 8.000 9.250 8.000 10.250 10.000 10.250 10.000 13.750
                 8.000 13.750 8.000 14.750 10.000 14.750 10.000 18.250 8.000 18.250
                 8.000 19.250 10.000 19.250 10.000 22.750 8.000 22.750 8.000 23.750
                 10.000 23.750 10.000 27.250 8.000 27.250 8.000 28.250 10.000 28.250
                 10.000 31.750 8.000 31.750 8.000 33.080 10.000 33.080 10.000 37.580
                 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750 7.000 9.250
                 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750 3.000 13.750
                 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250 3.000 19.250
                 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750 7.000 23.750
                 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250 7.000 31.750
                 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580 0.000 37.580
                 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750 0.000 28.250
                 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750 2.000 23.750
                 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250 2.000 18.250
                 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750 0.000 13.750
                 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750 2.000 5.750
                 2.000 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 4.750 8.000 4.750 8.000 5.750 10.000 5.750
                 10.000 9.250 8.000 9.250 8.000 10.250 10.000 10.250 10.000 13.750
                 8.000 13.750 8.000 14.750 10.000 14.750 10.000 18.250 8.000 18.250
                 8.000 19.250 10.000 19.250 10.000 22.750 8.000 22.750 8.000 23.750
                 10.000 23.750 10.000 27.250 8.000 27.250 8.000 28.250 10.000 28.250
                 10.000 31.750 8.000 31.750 8.000 33.080 10.000 33.080 10.000 37.580
                 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750 7.000 9.250
                 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750 3.000 13.750
                 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250 3.000 19.250
                 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750 7.000 23.750
                 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250 7.000 31.750
                 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580 0.000 37.580
                 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750 0.000 28.250
                 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750 2.000 23.750
                 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250 2.000 18.250
                 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750 0.000 13.750
                 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750 2.000 5.750
                 2.000 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 10.000 1.250 10.000 4.750 8.000 4.750 8.000 5.750 10.000 5.750
                 10.000 9.250 8.000 9.250 8.000 10.250 10.000 10.250 10.000 13.750
                 8.000 13.750 8.000 14.750 10.000 14.750 10.000 18.250 8.000 18.250
                 8.000 19.250 10.000 19.250 10.000 22.750 8.000 22.750 8.000 23.750
                 10.000 23.750 10.000 27.250 8.000 27.250 8.000 28.250 10.000 28.250
                 10.000 31.750 8.000 31.750 8.000 33.080 10.000 33.080 10.000 37.580
                 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750 7.000 9.250
                 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750 3.000 13.750
                 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250 3.000 19.250
                 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750 7.000 23.750
                 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250 7.000 31.750
                 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580 0.000 37.580
                 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750 0.000 28.250
                 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750 2.000 23.750
                 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250 2.000 18.250
                 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750 0.000 13.750
                 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750 2.000 5.750
                 2.000 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 8.000 87.170 8.000 88.020
                 10.000 88.020 10.000 91.520 8.000 91.520 8.000 92.370 10.000 92.370
                 10.000 95.870 8.000 95.870 8.000 96.720 10.000 96.720 10.000 100.220
                 8.000 100.220 8.000 101.070 10.000 101.070 10.000 104.570 8.000 104.570
                 8.000 105.420 10.000 105.420 10.000 108.920 8.000 108.920 8.000 109.770
                 10.000 109.770 10.000 113.270 8.000 113.270 8.000 114.010 10.000 114.010
                 10.000 117.510 7.000 117.510 7.000 87.170 3.000 87.170 3.000 88.020
                 7.000 88.020 7.000 91.520 3.000 91.520 3.000 92.370 7.000 92.370
                 7.000 95.870 3.000 95.870 3.000 96.720 7.000 96.720 7.000 100.220
                 3.000 100.220 3.000 101.070 7.000 101.070 7.000 104.570 3.000 104.570
                 3.000 105.420 7.000 105.420 7.000 108.920 3.000 108.920 3.000 109.770
                 7.000 109.770 7.000 113.270 3.000 113.270 3.000 114.010 7.000 114.010
                 7.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 8.000 87.170 8.000 88.020
                 10.000 88.020 10.000 91.520 8.000 91.520 8.000 92.370 10.000 92.370
                 10.000 95.870 8.000 95.870 8.000 96.720 10.000 96.720 10.000 100.220
                 8.000 100.220 8.000 101.070 10.000 101.070 10.000 104.570 8.000 104.570
                 8.000 105.420 10.000 105.420 10.000 108.920 8.000 108.920 8.000 109.770
                 10.000 109.770 10.000 113.270 8.000 113.270 8.000 114.010 10.000 114.010
                 10.000 117.510 7.000 117.510 7.000 87.170 3.000 87.170 3.000 88.020
                 7.000 88.020 7.000 91.520 3.000 91.520 3.000 92.370 7.000 92.370
                 7.000 95.870 3.000 95.870 3.000 96.720 7.000 96.720 7.000 100.220
                 3.000 100.220 3.000 101.070 7.000 101.070 7.000 104.570 3.000 104.570
                 3.000 105.420 7.000 105.420 7.000 108.920 3.000 108.920 3.000 109.770
                 7.000 109.770 7.000 113.270 3.000 113.270 3.000 114.010 7.000 114.010
                 7.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 8.000 87.170 8.000 88.020
                 10.000 88.020 10.000 91.520 8.000 91.520 8.000 92.370 10.000 92.370
                 10.000 95.870 8.000 95.870 8.000 96.720 10.000 96.720 10.000 100.220
                 8.000 100.220 8.000 101.070 10.000 101.070 10.000 104.570 8.000 104.570
                 8.000 105.420 10.000 105.420 10.000 108.920 8.000 108.920 8.000 109.770
                 10.000 109.770 10.000 113.270 8.000 113.270 8.000 114.010 10.000 114.010
                 10.000 117.510 7.000 117.510 7.000 87.170 3.000 87.170 3.000 88.020
                 7.000 88.020 7.000 91.520 3.000 91.520 3.000 92.370 7.000 92.370
                 7.000 95.870 3.000 95.870 3.000 96.720 7.000 96.720 7.000 100.220
                 3.000 100.220 3.000 101.070 7.000 101.070 7.000 104.570 3.000 104.570
                 3.000 105.420 7.000 105.420 7.000 108.920 3.000 108.920 3.000 109.770
                 7.000 109.770 7.000 113.270 3.000 113.270 3.000 114.010 7.000 114.010
                 7.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 8.000 87.170 8.000 88.020
                 10.000 88.020 10.000 91.520 8.000 91.520 8.000 92.370 10.000 92.370
                 10.000 95.870 8.000 95.870 8.000 96.720 10.000 96.720 10.000 100.220
                 8.000 100.220 8.000 101.070 10.000 101.070 10.000 104.570 8.000 104.570
                 8.000 105.420 10.000 105.420 10.000 108.920 8.000 108.920 8.000 109.770
                 10.000 109.770 10.000 113.270 8.000 113.270 8.000 114.010 10.000 114.010
                 10.000 117.510 7.000 117.510 7.000 87.170 3.000 87.170 3.000 88.020
                 7.000 88.020 7.000 91.520 3.000 91.520 3.000 92.370 7.000 92.370
                 7.000 95.870 3.000 95.870 3.000 96.720 7.000 96.720 7.000 100.220
                 3.000 100.220 3.000 101.070 7.000 101.070 7.000 104.570 3.000 104.570
                 3.000 105.420 7.000 105.420 7.000 108.920 3.000 108.920 3.000 109.770
                 7.000 109.770 7.000 113.270 3.000 113.270 3.000 114.010 7.000 114.010
                 7.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 10.000 83.670 10.000 87.170 8.000 87.170 8.000 88.020
                 10.000 88.020 10.000 91.520 8.000 91.520 8.000 92.370 10.000 92.370
                 10.000 95.870 8.000 95.870 8.000 96.720 10.000 96.720 10.000 100.220
                 8.000 100.220 8.000 101.070 10.000 101.070 10.000 104.570 8.000 104.570
                 8.000 105.420 10.000 105.420 10.000 108.920 7.000 108.920 7.000 87.170
                 3.000 87.170 3.000 88.020 7.000 88.020 7.000 91.520 3.000 91.520
                 3.000 92.370 7.000 92.370 7.000 95.870 3.000 95.870 3.000 96.720
                 7.000 96.720 7.000 100.220 3.000 100.220 3.000 101.070 7.000 101.070
                 7.000 104.570 3.000 104.570 3.000 105.420 7.000 105.420 7.000 108.920
                 0.000 108.920 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570
                 0.000 101.070 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720
                 2.000 96.720 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370
                 2.000 91.520 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 8.000 44.475 8.000 45.475
                 10.000 45.475 10.000 48.975 8.000 48.975 8.000 49.975 10.000 49.975
                 10.000 53.475 8.000 53.475 8.000 54.475 10.000 54.475 10.000 57.975
                 8.000 57.975 8.000 58.975 10.000 58.975 10.000 62.475 8.000 62.475
                 8.000 63.475 10.000 63.475 10.000 66.975 8.000 66.975 8.000 67.975
                 10.000 67.975 10.000 71.475 8.000 71.475 8.000 72.475 10.000 72.475
                 10.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 8.000 44.475 8.000 45.475
                 10.000 45.475 10.000 48.975 8.000 48.975 8.000 49.975 10.000 49.975
                 10.000 53.475 8.000 53.475 8.000 54.475 10.000 54.475 10.000 57.975
                 8.000 57.975 8.000 58.975 10.000 58.975 10.000 62.475 8.000 62.475
                 8.000 63.475 10.000 63.475 10.000 66.975 8.000 66.975 8.000 67.975
                 10.000 67.975 10.000 71.475 8.000 71.475 8.000 72.475 10.000 72.475
                 10.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 8.000 44.475 8.000 45.475
                 10.000 45.475 10.000 48.975 8.000 48.975 8.000 49.975 10.000 49.975
                 10.000 53.475 8.000 53.475 8.000 54.475 10.000 54.475 10.000 57.975
                 8.000 57.975 8.000 58.975 10.000 58.975 10.000 62.475 8.000 62.475
                 8.000 63.475 10.000 63.475 10.000 66.975 8.000 66.975 8.000 67.975
                 10.000 67.975 10.000 71.475 8.000 71.475 8.000 72.475 10.000 72.475
                 10.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 8.000 44.475 8.000 45.475
                 10.000 45.475 10.000 48.975 8.000 48.975 8.000 49.975 10.000 49.975
                 10.000 53.475 8.000 53.475 8.000 54.475 10.000 54.475 10.000 57.975
                 8.000 57.975 8.000 58.975 10.000 58.975 10.000 62.475 8.000 62.475
                 8.000 63.475 10.000 63.475 10.000 66.975 8.000 66.975 8.000 67.975
                 10.000 67.975 10.000 71.475 8.000 71.475 8.000 72.475 10.000 72.475
                 10.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 10.000 82.975 ;
                POLYGON  0.000 40.975 10.000 40.975 10.000 44.475 8.000 44.475 8.000 45.475
                 10.000 45.475 10.000 48.975 8.000 48.975 8.000 49.975 10.000 49.975
                 10.000 53.475 8.000 53.475 8.000 54.475 10.000 54.475 10.000 57.975
                 8.000 57.975 8.000 58.975 10.000 58.975 10.000 62.475 8.000 62.475
                 8.000 63.475 10.000 63.475 10.000 66.975 8.000 66.975 8.000 67.975
                 10.000 67.975 10.000 71.475 8.000 71.475 8.000 72.475 10.000 72.475
                 10.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 10.000 109.770 10.000 113.270 8.000 113.270 8.000 114.010
                 10.000 114.010 10.000 117.510 7.000 117.510 7.000 113.270 3.000 113.270
                 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510 0.000 114.010
                 2.000 114.010 2.000 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 10.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA2 ;
        RECT  8.000 1.250 10.000 4.750 ;
        RECT  8.000 5.750 10.000 9.250 ;
        RECT  8.000 10.250 10.000 13.750 ;
        RECT  8.000 14.750 10.000 18.250 ;
        RECT  8.000 19.250 10.000 22.750 ;
        RECT  8.000 23.750 10.000 27.250 ;
        RECT  8.000 28.250 10.000 31.750 ;
        RECT  8.000 33.080 10.000 37.580 ;
        RECT  8.000 40.975 10.000 44.475 ;
        RECT  8.000 45.475 10.000 48.975 ;
        RECT  8.000 49.975 10.000 53.475 ;
        RECT  8.000 54.475 10.000 57.975 ;
        RECT  8.000 58.975 10.000 62.475 ;
        RECT  8.000 63.475 10.000 66.975 ;
        RECT  8.000 67.975 10.000 71.475 ;
        RECT  8.000 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  8.000 83.670 10.000 87.170 ;
        RECT  8.000 88.020 10.000 91.520 ;
        RECT  8.000 92.370 10.000 95.870 ;
        RECT  8.000 96.720 10.000 100.220 ;
        RECT  8.000 101.070 10.000 104.570 ;
        RECT  8.000 105.420 10.000 108.920 ;
        RECT  8.000 109.770 10.000 113.270 ;
        RECT  8.000 114.010 10.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 108.920 ;
        RECT  7.000 109.770 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 108.920 ;
        RECT  2.000 109.770 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA3 ;
        RECT  8.000 1.250 10.000 4.750 ;
        RECT  8.000 5.750 10.000 9.250 ;
        RECT  8.000 10.250 10.000 13.750 ;
        RECT  8.000 14.750 10.000 18.250 ;
        RECT  8.000 19.250 10.000 22.750 ;
        RECT  8.000 23.750 10.000 27.250 ;
        RECT  8.000 28.250 10.000 31.750 ;
        RECT  8.000 33.080 10.000 37.580 ;
        RECT  8.000 40.975 10.000 44.475 ;
        RECT  8.000 45.475 10.000 48.975 ;
        RECT  8.000 49.975 10.000 53.475 ;
        RECT  8.000 54.475 10.000 57.975 ;
        RECT  8.000 58.975 10.000 62.475 ;
        RECT  8.000 63.475 10.000 66.975 ;
        RECT  8.000 67.975 10.000 71.475 ;
        RECT  8.000 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  8.000 83.670 10.000 87.170 ;
        RECT  8.000 88.020 10.000 91.520 ;
        RECT  8.000 92.370 10.000 95.870 ;
        RECT  8.000 96.720 10.000 100.220 ;
        RECT  8.000 101.070 10.000 104.570 ;
        RECT  8.000 105.420 10.000 108.920 ;
        RECT  8.000 109.770 10.000 113.270 ;
        RECT  8.000 114.010 10.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA4 ;
        RECT  8.000 1.250 10.000 4.750 ;
        RECT  8.000 5.750 10.000 9.250 ;
        RECT  8.000 10.250 10.000 13.750 ;
        RECT  8.000 14.750 10.000 18.250 ;
        RECT  8.000 19.250 10.000 22.750 ;
        RECT  8.000 23.750 10.000 27.250 ;
        RECT  8.000 28.250 10.000 31.750 ;
        RECT  8.000 33.080 10.000 37.580 ;
        RECT  8.000 40.975 10.000 44.475 ;
        RECT  8.000 45.475 10.000 48.975 ;
        RECT  8.000 49.975 10.000 53.475 ;
        RECT  8.000 54.475 10.000 57.975 ;
        RECT  8.000 58.975 10.000 62.475 ;
        RECT  8.000 63.475 10.000 66.975 ;
        RECT  8.000 67.975 10.000 71.475 ;
        RECT  8.000 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  8.000 83.670 10.000 87.170 ;
        RECT  8.000 88.020 10.000 91.520 ;
        RECT  8.000 92.370 10.000 95.870 ;
        RECT  8.000 96.720 10.000 100.220 ;
        RECT  8.000 101.070 10.000 104.570 ;
        RECT  8.000 105.420 10.000 108.920 ;
        RECT  8.000 109.770 10.000 113.270 ;
        RECT  8.000 114.010 10.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA5 ;
        RECT  8.000 1.250 10.000 4.750 ;
        RECT  8.000 5.750 10.000 9.250 ;
        RECT  8.000 10.250 10.000 13.750 ;
        RECT  8.000 14.750 10.000 18.250 ;
        RECT  8.000 19.250 10.000 22.750 ;
        RECT  8.000 23.750 10.000 27.250 ;
        RECT  8.000 28.250 10.000 31.750 ;
        RECT  8.000 33.080 10.000 37.580 ;
        RECT  8.000 40.975 10.000 44.475 ;
        RECT  8.000 45.475 10.000 48.975 ;
        RECT  8.000 49.975 10.000 53.475 ;
        RECT  8.000 54.475 10.000 57.975 ;
        RECT  8.000 58.975 10.000 62.475 ;
        RECT  8.000 63.475 10.000 66.975 ;
        RECT  8.000 67.975 10.000 71.475 ;
        RECT  8.000 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  8.000 83.670 10.000 87.170 ;
        RECT  8.000 88.020 10.000 91.520 ;
        RECT  8.000 92.370 10.000 95.870 ;
        RECT  8.000 96.720 10.000 100.220 ;
        RECT  8.000 101.070 10.000 104.570 ;
        RECT  8.000 105.420 10.000 108.920 ;
        RECT  8.000 109.770 10.000 113.270 ;
        RECT  8.000 114.010 10.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 10.000 120.000 ;
        LAYER VIA6 ;
        RECT  8.000 1.250 10.000 4.750 ;
        RECT  8.000 5.750 10.000 9.250 ;
        RECT  8.000 10.250 10.000 13.750 ;
        RECT  8.000 14.750 10.000 18.250 ;
        RECT  8.000 19.250 10.000 22.750 ;
        RECT  8.000 23.750 10.000 27.250 ;
        RECT  8.000 28.250 10.000 31.750 ;
        RECT  8.000 33.080 10.000 37.580 ;
        RECT  8.000 40.975 10.000 44.475 ;
        RECT  8.000 45.475 10.000 48.975 ;
        RECT  8.000 49.975 10.000 53.475 ;
        RECT  8.000 54.475 10.000 57.975 ;
        RECT  8.000 58.975 10.000 62.475 ;
        RECT  8.000 63.475 10.000 66.975 ;
        RECT  8.000 67.975 10.000 71.475 ;
        RECT  8.000 72.475 10.000 75.975 ;
        RECT  0.000 79.975 10.000 82.975 ;
        RECT  8.000 83.670 10.000 87.170 ;
        RECT  8.000 88.020 10.000 91.520 ;
        RECT  8.000 92.370 10.000 95.870 ;
        RECT  8.000 96.720 10.000 100.220 ;
        RECT  8.000 101.070 10.000 104.570 ;
        RECT  8.000 105.420 10.000 108.920 ;
        RECT  8.000 109.770 10.000 113.270 ;
        RECT  8.000 114.010 10.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 10.000 120.000 ;
    END
END PFILLER10_G

MACRO PFILLER1A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER1A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        LAYER M6 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        LAYER M5 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        LAYER M4 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        LAYER M3 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 1.250 1.000 5.750 ;
        RECT  0.000 7.250 1.000 11.750 ;
        RECT  0.000 13.250 1.000 17.750 ;
        RECT  0.000 19.250 1.000 23.750 ;
        RECT  0.000 25.250 1.000 29.750 ;
        RECT  0.000 31.250 1.000 35.750 ;
        RECT  0.000 36.750 1.000 39.290 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 1.000 120.000 ;
    END
END PFILLER1A_G

MACRO PFILLER1_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER1_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        LAYER M6 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        LAYER M5 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        LAYER M4 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        LAYER M3 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M4 ;
        RECT  0.000 109.770 1.000 113.270 ;
        LAYER M5 ;
        RECT  0.000 109.770 1.000 113.270 ;
        LAYER M6 ;
        RECT  0.000 109.770 1.000 113.270 ;
        LAYER M7 ;
        RECT  0.000 109.770 1.000 113.270 ;
        LAYER M4 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 1.000 87.170 ;
        LAYER M4 ;
        RECT  0.000 83.670 1.000 87.170 ;
        LAYER M5 ;
        RECT  0.000 83.670 1.000 87.170 ;
        LAYER M6 ;
        RECT  0.000 83.670 1.000 87.170 ;
        LAYER M7 ;
        RECT  0.000 83.670 1.000 87.170 ;
        LAYER M3 ;
        RECT  0.000 88.020 1.000 91.520 ;
        LAYER M4 ;
        RECT  0.000 88.020 1.000 91.520 ;
        LAYER M5 ;
        RECT  0.000 88.020 1.000 91.520 ;
        LAYER M6 ;
        RECT  0.000 88.020 1.000 91.520 ;
        LAYER M7 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        LAYER M6 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        LAYER M5 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        LAYER M4 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        LAYER M3 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 1.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        LAYER M4 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 1.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 1.250 1.000 4.750 ;
        RECT  0.000 5.750 1.000 9.250 ;
        RECT  0.000 10.250 1.000 13.750 ;
        RECT  0.000 14.750 1.000 18.250 ;
        RECT  0.000 19.250 1.000 22.750 ;
        RECT  0.000 23.750 1.000 27.250 ;
        RECT  0.000 28.250 1.000 31.750 ;
        RECT  0.000 33.080 1.000 37.580 ;
        RECT  0.000 40.975 1.000 44.475 ;
        RECT  0.000 45.475 1.000 48.975 ;
        RECT  0.000 49.975 1.000 53.475 ;
        RECT  0.000 54.475 1.000 57.975 ;
        RECT  0.000 58.975 1.000 62.475 ;
        RECT  0.000 63.475 1.000 66.975 ;
        RECT  0.000 67.975 1.000 71.475 ;
        RECT  0.000 72.475 1.000 75.975 ;
        RECT  0.000 79.975 1.000 82.975 ;
        RECT  0.000 83.670 1.000 87.170 ;
        RECT  0.000 88.020 1.000 91.520 ;
        RECT  0.000 92.370 1.000 95.870 ;
        RECT  0.000 96.720 1.000 100.220 ;
        RECT  0.000 101.070 1.000 104.570 ;
        RECT  0.000 105.420 1.000 108.920 ;
        RECT  0.000 109.770 1.000 113.270 ;
        RECT  0.000 114.010 1.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 1.000 120.000 ;
    END
END PFILLER1_G

MACRO PFILLER20A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER20A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 11.380 87.170 11.380 88.020
                 20.000 88.020 20.000 91.520 11.380 91.520 11.380 92.370 20.000 92.370
                 20.000 95.870 11.380 95.870 11.380 96.720 20.000 96.720 20.000 100.220
                 11.380 100.220 11.380 101.070 20.000 101.070 20.000 104.570
                 11.380 104.570 11.380 105.420 20.000 105.420 20.000 108.920
                 11.380 108.920 11.380 109.770 20.000 109.770 20.000 113.270
                 11.380 113.270 11.380 114.010 20.000 114.010 20.000 117.510
                 0.000 117.510 0.000 114.010 8.620 114.010 8.620 113.270 0.000 113.270
                 0.000 109.770 8.620 109.770 8.620 108.920 0.000 108.920 0.000 105.420
                 8.620 105.420 8.620 104.570 0.000 104.570 0.000 101.070 8.620 101.070
                 8.620 100.220 0.000 100.220 0.000 96.720 8.620 96.720 8.620 95.870
                 0.000 95.870 0.000 92.370 8.620 92.370 8.620 91.520 0.000 91.520
                 0.000 88.020 8.620 88.020 8.620 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 11.380 87.170 11.380 88.020
                 20.000 88.020 20.000 91.520 11.380 91.520 11.380 92.370 20.000 92.370
                 20.000 95.870 11.380 95.870 11.380 96.720 20.000 96.720 20.000 100.220
                 11.380 100.220 11.380 101.070 20.000 101.070 20.000 104.570
                 11.380 104.570 11.380 105.420 20.000 105.420 20.000 108.920
                 11.380 108.920 11.380 109.770 20.000 109.770 20.000 113.270
                 11.380 113.270 11.380 114.010 20.000 114.010 20.000 117.510
                 0.000 117.510 0.000 114.010 8.620 114.010 8.620 113.270 0.000 113.270
                 0.000 109.770 8.620 109.770 8.620 108.920 0.000 108.920 0.000 105.420
                 8.620 105.420 8.620 104.570 0.000 104.570 0.000 101.070 8.620 101.070
                 8.620 100.220 0.000 100.220 0.000 96.720 8.620 96.720 8.620 95.870
                 0.000 95.870 0.000 92.370 8.620 92.370 8.620 91.520 0.000 91.520
                 0.000 88.020 8.620 88.020 8.620 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 11.380 87.170 11.380 88.020
                 20.000 88.020 20.000 91.520 11.380 91.520 11.380 92.370 20.000 92.370
                 20.000 95.870 11.380 95.870 11.380 96.720 20.000 96.720 20.000 100.220
                 11.380 100.220 11.380 101.070 20.000 101.070 20.000 104.570
                 11.380 104.570 11.380 105.420 20.000 105.420 20.000 108.920
                 11.380 108.920 11.380 109.770 20.000 109.770 20.000 113.270
                 11.380 113.270 11.380 114.010 20.000 114.010 20.000 117.510
                 0.000 117.510 0.000 114.010 8.620 114.010 8.620 113.270 0.000 113.270
                 0.000 109.770 8.620 109.770 8.620 108.920 0.000 108.920 0.000 105.420
                 8.620 105.420 8.620 104.570 0.000 104.570 0.000 101.070 8.620 101.070
                 8.620 100.220 0.000 100.220 0.000 96.720 8.620 96.720 8.620 95.870
                 0.000 95.870 0.000 92.370 8.620 92.370 8.620 91.520 0.000 91.520
                 0.000 88.020 8.620 88.020 8.620 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 11.380 87.170 11.380 88.020
                 20.000 88.020 20.000 91.520 11.380 91.520 11.380 92.370 20.000 92.370
                 20.000 95.870 11.380 95.870 11.380 96.720 20.000 96.720 20.000 100.220
                 11.380 100.220 11.380 101.070 20.000 101.070 20.000 104.570
                 11.380 104.570 11.380 105.420 20.000 105.420 20.000 108.920
                 11.380 108.920 11.380 109.770 20.000 109.770 20.000 113.270
                 11.380 113.270 11.380 114.010 20.000 114.010 20.000 117.510
                 0.000 117.510 0.000 114.010 8.620 114.010 8.620 113.270 0.000 113.270
                 0.000 109.770 8.620 109.770 8.620 108.920 0.000 108.920 0.000 105.420
                 8.620 105.420 8.620 104.570 0.000 104.570 0.000 101.070 8.620 101.070
                 8.620 100.220 0.000 100.220 0.000 96.720 8.620 96.720 8.620 95.870
                 0.000 95.870 0.000 92.370 8.620 92.370 8.620 91.520 0.000 91.520
                 0.000 88.020 8.620 88.020 8.620 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 11.380 87.170 11.380 88.020
                 20.000 88.020 20.000 91.520 11.380 91.520 11.380 92.370 20.000 92.370
                 20.000 95.870 11.380 95.870 11.380 96.720 20.000 96.720 20.000 100.220
                 11.380 100.220 11.380 101.070 20.000 101.070 20.000 104.570
                 11.380 104.570 11.380 105.420 20.000 105.420 20.000 108.920
                 11.380 108.920 11.380 109.770 20.000 109.770 20.000 113.270
                 11.380 113.270 11.380 114.010 20.000 114.010 20.000 117.510
                 0.000 117.510 0.000 114.010 8.620 114.010 8.620 113.270 0.000 113.270
                 0.000 109.770 8.620 109.770 8.620 108.920 0.000 108.920 0.000 105.420
                 8.620 105.420 8.620 104.570 0.000 104.570 0.000 101.070 8.620 101.070
                 8.620 100.220 0.000 100.220 0.000 96.720 8.620 96.720 8.620 95.870
                 0.000 95.870 0.000 92.370 8.620 92.370 8.620 91.520 0.000 91.520
                 0.000 88.020 8.620 88.020 8.620 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 5.750 11.380 5.750 11.380 7.250
                 20.000 7.250 20.000 11.750 11.380 11.750 11.380 13.250 20.000 13.250
                 20.000 17.750 11.380 17.750 11.380 19.250 20.000 19.250 20.000 23.750
                 11.380 23.750 11.380 25.250 20.000 25.250 20.000 29.750 11.380 29.750
                 11.380 31.250 20.000 31.250 20.000 35.750 11.380 35.750 11.380 36.750
                 20.000 36.750 20.000 39.290 0.000 39.290 0.000 36.750 8.620 36.750
                 8.620 35.750 0.000 35.750 0.000 31.250 8.620 31.250 8.620 29.750
                 0.000 29.750 0.000 25.250 8.620 25.250 8.620 23.750 0.000 23.750
                 0.000 19.250 8.620 19.250 8.620 17.750 0.000 17.750 0.000 13.250
                 8.620 13.250 8.620 11.750 0.000 11.750 0.000 7.250 8.620 7.250 8.620 5.750
                 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 5.750 11.380 5.750 11.380 7.250
                 20.000 7.250 20.000 11.750 11.380 11.750 11.380 13.250 20.000 13.250
                 20.000 17.750 11.380 17.750 11.380 19.250 20.000 19.250 20.000 23.750
                 11.380 23.750 11.380 25.250 20.000 25.250 20.000 29.750 11.380 29.750
                 11.380 31.250 20.000 31.250 20.000 35.750 11.380 35.750 11.380 36.750
                 20.000 36.750 20.000 39.290 0.000 39.290 0.000 36.750 8.620 36.750
                 8.620 35.750 0.000 35.750 0.000 31.250 8.620 31.250 8.620 29.750
                 0.000 29.750 0.000 25.250 8.620 25.250 8.620 23.750 0.000 23.750
                 0.000 19.250 8.620 19.250 8.620 17.750 0.000 17.750 0.000 13.250
                 8.620 13.250 8.620 11.750 0.000 11.750 0.000 7.250 8.620 7.250 8.620 5.750
                 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 5.750 11.380 5.750 11.380 7.250
                 20.000 7.250 20.000 11.750 11.380 11.750 11.380 13.250 20.000 13.250
                 20.000 17.750 11.380 17.750 11.380 19.250 20.000 19.250 20.000 23.750
                 11.380 23.750 11.380 25.250 20.000 25.250 20.000 29.750 11.380 29.750
                 11.380 31.250 20.000 31.250 20.000 35.750 11.380 35.750 11.380 36.750
                 20.000 36.750 20.000 39.290 0.000 39.290 0.000 36.750 8.620 36.750
                 8.620 35.750 0.000 35.750 0.000 31.250 8.620 31.250 8.620 29.750
                 0.000 29.750 0.000 25.250 8.620 25.250 8.620 23.750 0.000 23.750
                 0.000 19.250 8.620 19.250 8.620 17.750 0.000 17.750 0.000 13.250
                 8.620 13.250 8.620 11.750 0.000 11.750 0.000 7.250 8.620 7.250 8.620 5.750
                 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 5.750 11.380 5.750 11.380 7.250
                 20.000 7.250 20.000 11.750 11.380 11.750 11.380 13.250 20.000 13.250
                 20.000 17.750 11.380 17.750 11.380 19.250 20.000 19.250 20.000 23.750
                 11.380 23.750 11.380 25.250 20.000 25.250 20.000 29.750 11.380 29.750
                 11.380 31.250 20.000 31.250 20.000 35.750 11.380 35.750 11.380 36.750
                 20.000 36.750 20.000 39.290 0.000 39.290 0.000 36.750 8.620 36.750
                 8.620 35.750 0.000 35.750 0.000 31.250 8.620 31.250 8.620 29.750
                 0.000 29.750 0.000 25.250 8.620 25.250 8.620 23.750 0.000 23.750
                 0.000 19.250 8.620 19.250 8.620 17.750 0.000 17.750 0.000 13.250
                 8.620 13.250 8.620 11.750 0.000 11.750 0.000 7.250 8.620 7.250 8.620 5.750
                 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 5.750 11.380 5.750 11.380 7.250
                 20.000 7.250 20.000 11.750 11.380 11.750 11.380 13.250 20.000 13.250
                 20.000 17.750 11.380 17.750 11.380 19.250 20.000 19.250 20.000 23.750
                 11.380 23.750 11.380 25.250 20.000 25.250 20.000 29.750 11.380 29.750
                 11.380 31.250 20.000 31.250 20.000 35.750 11.380 35.750 11.380 36.750
                 20.000 36.750 20.000 39.290 0.000 39.290 0.000 36.750 8.620 36.750
                 8.620 35.750 0.000 35.750 0.000 31.250 8.620 31.250 8.620 29.750
                 0.000 29.750 0.000 25.250 8.620 25.250 8.620 23.750 0.000 23.750
                 0.000 19.250 8.620 19.250 8.620 17.750 0.000 17.750 0.000 13.250
                 8.620 13.250 8.620 11.750 0.000 11.750 0.000 7.250 8.620 7.250 8.620 5.750
                 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 11.380 44.475 11.380 45.475
                 20.000 45.475 20.000 48.975 11.380 48.975 11.380 49.975 20.000 49.975
                 20.000 53.475 11.380 53.475 11.380 54.475 20.000 54.475 20.000 57.975
                 11.380 57.975 11.380 58.975 20.000 58.975 20.000 62.475 11.380 62.475
                 11.380 63.475 20.000 63.475 20.000 66.975 11.380 66.975 11.380 67.975
                 20.000 67.975 20.000 71.475 11.380 71.475 11.380 72.475 20.000 72.475
                 20.000 75.975 0.000 75.975 0.000 72.475 8.620 72.475 8.620 71.475
                 0.000 71.475 0.000 67.975 8.620 67.975 8.620 66.975 0.000 66.975
                 0.000 63.475 8.620 63.475 8.620 62.475 0.000 62.475 0.000 58.975
                 8.620 58.975 8.620 57.975 0.000 57.975 0.000 54.475 8.620 54.475
                 8.620 53.475 0.000 53.475 0.000 49.975 8.620 49.975 8.620 48.975
                 0.000 48.975 0.000 45.475 8.620 45.475 8.620 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 11.380 44.475 11.380 45.475
                 20.000 45.475 20.000 48.975 11.380 48.975 11.380 49.975 20.000 49.975
                 20.000 53.475 11.380 53.475 11.380 54.475 20.000 54.475 20.000 57.975
                 11.380 57.975 11.380 58.975 20.000 58.975 20.000 62.475 11.380 62.475
                 11.380 63.475 20.000 63.475 20.000 66.975 11.380 66.975 11.380 67.975
                 20.000 67.975 20.000 71.475 11.380 71.475 11.380 72.475 20.000 72.475
                 20.000 75.975 0.000 75.975 0.000 72.475 8.620 72.475 8.620 71.475
                 0.000 71.475 0.000 67.975 8.620 67.975 8.620 66.975 0.000 66.975
                 0.000 63.475 8.620 63.475 8.620 62.475 0.000 62.475 0.000 58.975
                 8.620 58.975 8.620 57.975 0.000 57.975 0.000 54.475 8.620 54.475
                 8.620 53.475 0.000 53.475 0.000 49.975 8.620 49.975 8.620 48.975
                 0.000 48.975 0.000 45.475 8.620 45.475 8.620 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 11.380 44.475 11.380 45.475
                 20.000 45.475 20.000 48.975 11.380 48.975 11.380 49.975 20.000 49.975
                 20.000 53.475 11.380 53.475 11.380 54.475 20.000 54.475 20.000 57.975
                 11.380 57.975 11.380 58.975 20.000 58.975 20.000 62.475 11.380 62.475
                 11.380 63.475 20.000 63.475 20.000 66.975 11.380 66.975 11.380 67.975
                 20.000 67.975 20.000 71.475 11.380 71.475 11.380 72.475 20.000 72.475
                 20.000 75.975 0.000 75.975 0.000 72.475 8.620 72.475 8.620 71.475
                 0.000 71.475 0.000 67.975 8.620 67.975 8.620 66.975 0.000 66.975
                 0.000 63.475 8.620 63.475 8.620 62.475 0.000 62.475 0.000 58.975
                 8.620 58.975 8.620 57.975 0.000 57.975 0.000 54.475 8.620 54.475
                 8.620 53.475 0.000 53.475 0.000 49.975 8.620 49.975 8.620 48.975
                 0.000 48.975 0.000 45.475 8.620 45.475 8.620 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 11.380 44.475 11.380 45.475
                 20.000 45.475 20.000 48.975 11.380 48.975 11.380 49.975 20.000 49.975
                 20.000 53.475 11.380 53.475 11.380 54.475 20.000 54.475 20.000 57.975
                 11.380 57.975 11.380 58.975 20.000 58.975 20.000 62.475 11.380 62.475
                 11.380 63.475 20.000 63.475 20.000 66.975 11.380 66.975 11.380 67.975
                 20.000 67.975 20.000 71.475 11.380 71.475 11.380 72.475 20.000 72.475
                 20.000 75.975 0.000 75.975 0.000 72.475 8.620 72.475 8.620 71.475
                 0.000 71.475 0.000 67.975 8.620 67.975 8.620 66.975 0.000 66.975
                 0.000 63.475 8.620 63.475 8.620 62.475 0.000 62.475 0.000 58.975
                 8.620 58.975 8.620 57.975 0.000 57.975 0.000 54.475 8.620 54.475
                 8.620 53.475 0.000 53.475 0.000 49.975 8.620 49.975 8.620 48.975
                 0.000 48.975 0.000 45.475 8.620 45.475 8.620 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 11.380 44.475 11.380 45.475
                 20.000 45.475 20.000 48.975 11.380 48.975 11.380 49.975 20.000 49.975
                 20.000 53.475 11.380 53.475 11.380 54.475 20.000 54.475 20.000 57.975
                 11.380 57.975 11.380 58.975 20.000 58.975 20.000 62.475 11.380 62.475
                 11.380 63.475 20.000 63.475 20.000 66.975 11.380 66.975 11.380 67.975
                 20.000 67.975 20.000 71.475 11.380 71.475 11.380 72.475 20.000 72.475
                 20.000 75.975 0.000 75.975 0.000 72.475 8.620 72.475 8.620 71.475
                 0.000 71.475 0.000 67.975 8.620 67.975 8.620 66.975 0.000 66.975
                 0.000 63.475 8.620 63.475 8.620 62.475 0.000 62.475 0.000 58.975
                 8.620 58.975 8.620 57.975 0.000 57.975 0.000 54.475 8.620 54.475
                 8.620 53.475 0.000 53.475 0.000 49.975 8.620 49.975 8.620 48.975
                 0.000 48.975 0.000 45.475 8.620 45.475 8.620 44.475 0.000 44.475 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA2 ;
        RECT  11.380 1.250 20.000 5.750 ;
        RECT  11.380 7.250 20.000 11.750 ;
        RECT  11.380 13.250 20.000 17.750 ;
        RECT  11.380 19.250 20.000 23.750 ;
        RECT  11.380 25.250 20.000 29.750 ;
        RECT  11.380 31.250 20.000 35.750 ;
        RECT  11.380 36.750 20.000 39.290 ;
        RECT  11.380 40.975 20.000 44.475 ;
        RECT  11.380 45.475 20.000 48.975 ;
        RECT  11.380 49.975 20.000 53.475 ;
        RECT  11.380 54.475 20.000 57.975 ;
        RECT  11.380 58.975 20.000 62.475 ;
        RECT  11.380 63.475 20.000 66.975 ;
        RECT  11.380 67.975 20.000 71.475 ;
        RECT  11.380 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  11.380 83.670 20.000 87.170 ;
        RECT  11.380 88.020 20.000 91.520 ;
        RECT  11.380 92.370 20.000 95.870 ;
        RECT  11.380 96.720 20.000 100.220 ;
        RECT  11.380 101.070 20.000 104.570 ;
        RECT  11.380 105.420 20.000 108.920 ;
        RECT  11.380 109.770 20.000 113.270 ;
        RECT  11.380 114.010 20.000 117.510 ;
        RECT  8.620 1.250 11.380 39.290 ;
        RECT  8.620 40.975 11.380 75.975 ;
        RECT  8.620 83.670 11.380 117.510 ;
        RECT  0.000 1.250 8.620 5.750 ;
        RECT  0.000 7.250 8.620 11.750 ;
        RECT  0.000 13.250 8.620 17.750 ;
        RECT  0.000 19.250 8.620 23.750 ;
        RECT  0.000 25.250 8.620 29.750 ;
        RECT  0.000 31.250 8.620 35.750 ;
        RECT  0.000 36.750 8.620 39.290 ;
        RECT  0.000 40.975 8.620 44.475 ;
        RECT  0.000 45.475 8.620 48.975 ;
        RECT  0.000 49.975 8.620 53.475 ;
        RECT  0.000 54.475 8.620 57.975 ;
        RECT  0.000 58.975 8.620 62.475 ;
        RECT  0.000 63.475 8.620 66.975 ;
        RECT  0.000 67.975 8.620 71.475 ;
        RECT  0.000 72.475 8.620 75.975 ;
        RECT  0.000 83.670 8.620 87.170 ;
        RECT  0.000 88.020 8.620 91.520 ;
        RECT  0.000 92.370 8.620 95.870 ;
        RECT  0.000 96.720 8.620 100.220 ;
        RECT  0.000 101.070 8.620 104.570 ;
        RECT  0.000 105.420 8.620 108.920 ;
        RECT  0.000 109.770 8.620 113.270 ;
        RECT  0.000 114.010 8.620 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA3 ;
        RECT  11.380 1.250 20.000 5.750 ;
        RECT  11.380 7.250 20.000 11.750 ;
        RECT  11.380 13.250 20.000 17.750 ;
        RECT  11.380 19.250 20.000 23.750 ;
        RECT  11.380 25.250 20.000 29.750 ;
        RECT  11.380 31.250 20.000 35.750 ;
        RECT  11.380 36.750 20.000 39.290 ;
        RECT  11.380 40.975 20.000 44.475 ;
        RECT  11.380 45.475 20.000 48.975 ;
        RECT  11.380 49.975 20.000 53.475 ;
        RECT  11.380 54.475 20.000 57.975 ;
        RECT  11.380 58.975 20.000 62.475 ;
        RECT  11.380 63.475 20.000 66.975 ;
        RECT  11.380 67.975 20.000 71.475 ;
        RECT  11.380 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  11.380 83.670 20.000 87.170 ;
        RECT  11.380 88.020 20.000 91.520 ;
        RECT  11.380 92.370 20.000 95.870 ;
        RECT  11.380 96.720 20.000 100.220 ;
        RECT  11.380 101.070 20.000 104.570 ;
        RECT  11.380 105.420 20.000 108.920 ;
        RECT  11.380 109.770 20.000 113.270 ;
        RECT  11.380 114.010 20.000 117.510 ;
        RECT  8.620 1.250 11.380 39.290 ;
        RECT  8.620 40.975 11.380 75.975 ;
        RECT  8.620 83.670 11.380 117.510 ;
        RECT  0.000 1.250 8.620 5.750 ;
        RECT  0.000 7.250 8.620 11.750 ;
        RECT  0.000 13.250 8.620 17.750 ;
        RECT  0.000 19.250 8.620 23.750 ;
        RECT  0.000 25.250 8.620 29.750 ;
        RECT  0.000 31.250 8.620 35.750 ;
        RECT  0.000 36.750 8.620 39.290 ;
        RECT  0.000 40.975 8.620 44.475 ;
        RECT  0.000 45.475 8.620 48.975 ;
        RECT  0.000 49.975 8.620 53.475 ;
        RECT  0.000 54.475 8.620 57.975 ;
        RECT  0.000 58.975 8.620 62.475 ;
        RECT  0.000 63.475 8.620 66.975 ;
        RECT  0.000 67.975 8.620 71.475 ;
        RECT  0.000 72.475 8.620 75.975 ;
        RECT  0.000 83.670 8.620 87.170 ;
        RECT  0.000 88.020 8.620 91.520 ;
        RECT  0.000 92.370 8.620 95.870 ;
        RECT  0.000 96.720 8.620 100.220 ;
        RECT  0.000 101.070 8.620 104.570 ;
        RECT  0.000 105.420 8.620 108.920 ;
        RECT  0.000 109.770 8.620 113.270 ;
        RECT  0.000 114.010 8.620 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA4 ;
        RECT  11.380 1.250 20.000 5.750 ;
        RECT  11.380 7.250 20.000 11.750 ;
        RECT  11.380 13.250 20.000 17.750 ;
        RECT  11.380 19.250 20.000 23.750 ;
        RECT  11.380 25.250 20.000 29.750 ;
        RECT  11.380 31.250 20.000 35.750 ;
        RECT  11.380 36.750 20.000 39.290 ;
        RECT  11.380 40.975 20.000 44.475 ;
        RECT  11.380 45.475 20.000 48.975 ;
        RECT  11.380 49.975 20.000 53.475 ;
        RECT  11.380 54.475 20.000 57.975 ;
        RECT  11.380 58.975 20.000 62.475 ;
        RECT  11.380 63.475 20.000 66.975 ;
        RECT  11.380 67.975 20.000 71.475 ;
        RECT  11.380 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  11.380 83.670 20.000 87.170 ;
        RECT  11.380 88.020 20.000 91.520 ;
        RECT  11.380 92.370 20.000 95.870 ;
        RECT  11.380 96.720 20.000 100.220 ;
        RECT  11.380 101.070 20.000 104.570 ;
        RECT  11.380 105.420 20.000 108.920 ;
        RECT  11.380 109.770 20.000 113.270 ;
        RECT  11.380 114.010 20.000 117.510 ;
        RECT  8.620 1.250 11.380 39.290 ;
        RECT  8.620 40.975 11.380 75.975 ;
        RECT  8.620 83.670 11.380 117.510 ;
        RECT  0.000 1.250 8.620 5.750 ;
        RECT  0.000 7.250 8.620 11.750 ;
        RECT  0.000 13.250 8.620 17.750 ;
        RECT  0.000 19.250 8.620 23.750 ;
        RECT  0.000 25.250 8.620 29.750 ;
        RECT  0.000 31.250 8.620 35.750 ;
        RECT  0.000 36.750 8.620 39.290 ;
        RECT  0.000 40.975 8.620 44.475 ;
        RECT  0.000 45.475 8.620 48.975 ;
        RECT  0.000 49.975 8.620 53.475 ;
        RECT  0.000 54.475 8.620 57.975 ;
        RECT  0.000 58.975 8.620 62.475 ;
        RECT  0.000 63.475 8.620 66.975 ;
        RECT  0.000 67.975 8.620 71.475 ;
        RECT  0.000 72.475 8.620 75.975 ;
        RECT  0.000 83.670 8.620 87.170 ;
        RECT  0.000 88.020 8.620 91.520 ;
        RECT  0.000 92.370 8.620 95.870 ;
        RECT  0.000 96.720 8.620 100.220 ;
        RECT  0.000 101.070 8.620 104.570 ;
        RECT  0.000 105.420 8.620 108.920 ;
        RECT  0.000 109.770 8.620 113.270 ;
        RECT  0.000 114.010 8.620 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA5 ;
        RECT  11.380 1.250 20.000 5.750 ;
        RECT  11.380 7.250 20.000 11.750 ;
        RECT  11.380 13.250 20.000 17.750 ;
        RECT  11.380 19.250 20.000 23.750 ;
        RECT  11.380 25.250 20.000 29.750 ;
        RECT  11.380 31.250 20.000 35.750 ;
        RECT  11.380 36.750 20.000 39.290 ;
        RECT  11.380 40.975 20.000 44.475 ;
        RECT  11.380 45.475 20.000 48.975 ;
        RECT  11.380 49.975 20.000 53.475 ;
        RECT  11.380 54.475 20.000 57.975 ;
        RECT  11.380 58.975 20.000 62.475 ;
        RECT  11.380 63.475 20.000 66.975 ;
        RECT  11.380 67.975 20.000 71.475 ;
        RECT  11.380 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  11.380 83.670 20.000 87.170 ;
        RECT  11.380 88.020 20.000 91.520 ;
        RECT  11.380 92.370 20.000 95.870 ;
        RECT  11.380 96.720 20.000 100.220 ;
        RECT  11.380 101.070 20.000 104.570 ;
        RECT  11.380 105.420 20.000 108.920 ;
        RECT  11.380 109.770 20.000 113.270 ;
        RECT  11.380 114.010 20.000 117.510 ;
        RECT  8.620 1.250 11.380 39.290 ;
        RECT  8.620 40.975 11.380 75.975 ;
        RECT  8.620 83.670 11.380 117.510 ;
        RECT  0.000 1.250 8.620 5.750 ;
        RECT  0.000 7.250 8.620 11.750 ;
        RECT  0.000 13.250 8.620 17.750 ;
        RECT  0.000 19.250 8.620 23.750 ;
        RECT  0.000 25.250 8.620 29.750 ;
        RECT  0.000 31.250 8.620 35.750 ;
        RECT  0.000 36.750 8.620 39.290 ;
        RECT  0.000 40.975 8.620 44.475 ;
        RECT  0.000 45.475 8.620 48.975 ;
        RECT  0.000 49.975 8.620 53.475 ;
        RECT  0.000 54.475 8.620 57.975 ;
        RECT  0.000 58.975 8.620 62.475 ;
        RECT  0.000 63.475 8.620 66.975 ;
        RECT  0.000 67.975 8.620 71.475 ;
        RECT  0.000 72.475 8.620 75.975 ;
        RECT  0.000 83.670 8.620 87.170 ;
        RECT  0.000 88.020 8.620 91.520 ;
        RECT  0.000 92.370 8.620 95.870 ;
        RECT  0.000 96.720 8.620 100.220 ;
        RECT  0.000 101.070 8.620 104.570 ;
        RECT  0.000 105.420 8.620 108.920 ;
        RECT  0.000 109.770 8.620 113.270 ;
        RECT  0.000 114.010 8.620 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA6 ;
        RECT  11.380 1.250 20.000 5.750 ;
        RECT  11.380 7.250 20.000 11.750 ;
        RECT  11.380 13.250 20.000 17.750 ;
        RECT  11.380 19.250 20.000 23.750 ;
        RECT  11.380 25.250 20.000 29.750 ;
        RECT  11.380 31.250 20.000 35.750 ;
        RECT  11.380 36.750 20.000 39.290 ;
        RECT  11.380 40.975 20.000 44.475 ;
        RECT  11.380 45.475 20.000 48.975 ;
        RECT  11.380 49.975 20.000 53.475 ;
        RECT  11.380 54.475 20.000 57.975 ;
        RECT  11.380 58.975 20.000 62.475 ;
        RECT  11.380 63.475 20.000 66.975 ;
        RECT  11.380 67.975 20.000 71.475 ;
        RECT  11.380 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  11.380 83.670 20.000 87.170 ;
        RECT  11.380 88.020 20.000 91.520 ;
        RECT  11.380 92.370 20.000 95.870 ;
        RECT  11.380 96.720 20.000 100.220 ;
        RECT  11.380 101.070 20.000 104.570 ;
        RECT  11.380 105.420 20.000 108.920 ;
        RECT  11.380 109.770 20.000 113.270 ;
        RECT  11.380 114.010 20.000 117.510 ;
        RECT  8.620 1.250 11.380 39.290 ;
        RECT  8.620 40.975 11.380 75.975 ;
        RECT  8.620 83.670 11.380 117.510 ;
        RECT  0.000 1.250 8.620 5.750 ;
        RECT  0.000 7.250 8.620 11.750 ;
        RECT  0.000 13.250 8.620 17.750 ;
        RECT  0.000 19.250 8.620 23.750 ;
        RECT  0.000 25.250 8.620 29.750 ;
        RECT  0.000 31.250 8.620 35.750 ;
        RECT  0.000 36.750 8.620 39.290 ;
        RECT  0.000 40.975 8.620 44.475 ;
        RECT  0.000 45.475 8.620 48.975 ;
        RECT  0.000 49.975 8.620 53.475 ;
        RECT  0.000 54.475 8.620 57.975 ;
        RECT  0.000 58.975 8.620 62.475 ;
        RECT  0.000 63.475 8.620 66.975 ;
        RECT  0.000 67.975 8.620 71.475 ;
        RECT  0.000 72.475 8.620 75.975 ;
        RECT  0.000 83.670 8.620 87.170 ;
        RECT  0.000 88.020 8.620 91.520 ;
        RECT  0.000 92.370 8.620 95.870 ;
        RECT  0.000 96.720 8.620 100.220 ;
        RECT  0.000 101.070 8.620 104.570 ;
        RECT  0.000 105.420 8.620 108.920 ;
        RECT  0.000 109.770 8.620 113.270 ;
        RECT  0.000 114.010 8.620 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 20.000 120.000 ;
    END
END PFILLER20A_G

MACRO PFILLER20_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER20_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 4.750 18.000 4.750 18.000 5.750
                 20.000 5.750 20.000 9.250 18.000 9.250 18.000 10.250 20.000 10.250
                 20.000 13.750 18.000 13.750 18.000 14.750 20.000 14.750 20.000 18.250
                 18.000 18.250 18.000 19.250 20.000 19.250 20.000 22.750 18.000 22.750
                 18.000 23.750 20.000 23.750 20.000 27.250 18.000 27.250 18.000 28.250
                 20.000 28.250 20.000 31.750 18.000 31.750 18.000 33.080 20.000 33.080
                 20.000 37.580 17.000 37.580 17.000 4.750 13.000 4.750 13.000 5.750
                 17.000 5.750 17.000 9.250 13.000 9.250 13.000 10.250 17.000 10.250
                 17.000 13.750 13.000 13.750 13.000 14.750 17.000 14.750 17.000 18.250
                 13.000 18.250 13.000 19.250 17.000 19.250 17.000 22.750 13.000 22.750
                 13.000 23.750 17.000 23.750 17.000 27.250 13.000 27.250 13.000 28.250
                 17.000 28.250 17.000 31.750 13.000 31.750 13.000 33.080 17.000 33.080
                 17.000 37.580 12.000 37.580 12.000 4.750 8.000 4.750 8.000 5.750
                 12.000 5.750 12.000 9.250 8.000 9.250 8.000 10.250 12.000 10.250
                 12.000 13.750 8.000 13.750 8.000 14.750 12.000 14.750 12.000 18.250
                 8.000 18.250 8.000 19.250 12.000 19.250 12.000 22.750 8.000 22.750
                 8.000 23.750 12.000 23.750 12.000 27.250 8.000 27.250 8.000 28.250
                 12.000 28.250 12.000 31.750 8.000 31.750 8.000 33.080 12.000 33.080
                 12.000 37.580 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750
                 7.000 9.250 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750
                 3.000 13.750 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250
                 3.000 19.250 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750
                 7.000 23.750 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250
                 7.000 31.750 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 4.750 18.000 4.750 18.000 5.750
                 20.000 5.750 20.000 9.250 18.000 9.250 18.000 10.250 20.000 10.250
                 20.000 13.750 18.000 13.750 18.000 14.750 20.000 14.750 20.000 18.250
                 18.000 18.250 18.000 19.250 20.000 19.250 20.000 22.750 18.000 22.750
                 18.000 23.750 20.000 23.750 20.000 27.250 18.000 27.250 18.000 28.250
                 20.000 28.250 20.000 31.750 18.000 31.750 18.000 33.080 20.000 33.080
                 20.000 37.580 17.000 37.580 17.000 4.750 13.000 4.750 13.000 5.750
                 17.000 5.750 17.000 9.250 13.000 9.250 13.000 10.250 17.000 10.250
                 17.000 13.750 13.000 13.750 13.000 14.750 17.000 14.750 17.000 18.250
                 13.000 18.250 13.000 19.250 17.000 19.250 17.000 22.750 13.000 22.750
                 13.000 23.750 17.000 23.750 17.000 27.250 13.000 27.250 13.000 28.250
                 17.000 28.250 17.000 31.750 13.000 31.750 13.000 33.080 17.000 33.080
                 17.000 37.580 12.000 37.580 12.000 4.750 8.000 4.750 8.000 5.750
                 12.000 5.750 12.000 9.250 8.000 9.250 8.000 10.250 12.000 10.250
                 12.000 13.750 8.000 13.750 8.000 14.750 12.000 14.750 12.000 18.250
                 8.000 18.250 8.000 19.250 12.000 19.250 12.000 22.750 8.000 22.750
                 8.000 23.750 12.000 23.750 12.000 27.250 8.000 27.250 8.000 28.250
                 12.000 28.250 12.000 31.750 8.000 31.750 8.000 33.080 12.000 33.080
                 12.000 37.580 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750
                 7.000 9.250 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750
                 3.000 13.750 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250
                 3.000 19.250 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750
                 7.000 23.750 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250
                 7.000 31.750 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 4.750 18.000 4.750 18.000 5.750
                 20.000 5.750 20.000 9.250 18.000 9.250 18.000 10.250 20.000 10.250
                 20.000 13.750 18.000 13.750 18.000 14.750 20.000 14.750 20.000 18.250
                 18.000 18.250 18.000 19.250 20.000 19.250 20.000 22.750 18.000 22.750
                 18.000 23.750 20.000 23.750 20.000 27.250 18.000 27.250 18.000 28.250
                 20.000 28.250 20.000 31.750 18.000 31.750 18.000 33.080 20.000 33.080
                 20.000 37.580 17.000 37.580 17.000 4.750 13.000 4.750 13.000 5.750
                 17.000 5.750 17.000 9.250 13.000 9.250 13.000 10.250 17.000 10.250
                 17.000 13.750 13.000 13.750 13.000 14.750 17.000 14.750 17.000 18.250
                 13.000 18.250 13.000 19.250 17.000 19.250 17.000 22.750 13.000 22.750
                 13.000 23.750 17.000 23.750 17.000 27.250 13.000 27.250 13.000 28.250
                 17.000 28.250 17.000 31.750 13.000 31.750 13.000 33.080 17.000 33.080
                 17.000 37.580 12.000 37.580 12.000 4.750 8.000 4.750 8.000 5.750
                 12.000 5.750 12.000 9.250 8.000 9.250 8.000 10.250 12.000 10.250
                 12.000 13.750 8.000 13.750 8.000 14.750 12.000 14.750 12.000 18.250
                 8.000 18.250 8.000 19.250 12.000 19.250 12.000 22.750 8.000 22.750
                 8.000 23.750 12.000 23.750 12.000 27.250 8.000 27.250 8.000 28.250
                 12.000 28.250 12.000 31.750 8.000 31.750 8.000 33.080 12.000 33.080
                 12.000 37.580 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750
                 7.000 9.250 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750
                 3.000 13.750 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250
                 3.000 19.250 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750
                 7.000 23.750 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250
                 7.000 31.750 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 4.750 18.000 4.750 18.000 5.750
                 20.000 5.750 20.000 9.250 18.000 9.250 18.000 10.250 20.000 10.250
                 20.000 13.750 18.000 13.750 18.000 14.750 20.000 14.750 20.000 18.250
                 18.000 18.250 18.000 19.250 20.000 19.250 20.000 22.750 18.000 22.750
                 18.000 23.750 20.000 23.750 20.000 27.250 18.000 27.250 18.000 28.250
                 20.000 28.250 20.000 31.750 18.000 31.750 18.000 33.080 20.000 33.080
                 20.000 37.580 17.000 37.580 17.000 4.750 13.000 4.750 13.000 5.750
                 17.000 5.750 17.000 9.250 13.000 9.250 13.000 10.250 17.000 10.250
                 17.000 13.750 13.000 13.750 13.000 14.750 17.000 14.750 17.000 18.250
                 13.000 18.250 13.000 19.250 17.000 19.250 17.000 22.750 13.000 22.750
                 13.000 23.750 17.000 23.750 17.000 27.250 13.000 27.250 13.000 28.250
                 17.000 28.250 17.000 31.750 13.000 31.750 13.000 33.080 17.000 33.080
                 17.000 37.580 12.000 37.580 12.000 4.750 8.000 4.750 8.000 5.750
                 12.000 5.750 12.000 9.250 8.000 9.250 8.000 10.250 12.000 10.250
                 12.000 13.750 8.000 13.750 8.000 14.750 12.000 14.750 12.000 18.250
                 8.000 18.250 8.000 19.250 12.000 19.250 12.000 22.750 8.000 22.750
                 8.000 23.750 12.000 23.750 12.000 27.250 8.000 27.250 8.000 28.250
                 12.000 28.250 12.000 31.750 8.000 31.750 8.000 33.080 12.000 33.080
                 12.000 37.580 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750
                 7.000 9.250 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750
                 3.000 13.750 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250
                 3.000 19.250 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750
                 7.000 23.750 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250
                 7.000 31.750 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 20.000 1.250 20.000 4.750 18.000 4.750 18.000 5.750
                 20.000 5.750 20.000 9.250 18.000 9.250 18.000 10.250 20.000 10.250
                 20.000 13.750 18.000 13.750 18.000 14.750 20.000 14.750 20.000 18.250
                 18.000 18.250 18.000 19.250 20.000 19.250 20.000 22.750 18.000 22.750
                 18.000 23.750 20.000 23.750 20.000 27.250 18.000 27.250 18.000 28.250
                 20.000 28.250 20.000 31.750 18.000 31.750 18.000 33.080 20.000 33.080
                 20.000 37.580 17.000 37.580 17.000 4.750 13.000 4.750 13.000 5.750
                 17.000 5.750 17.000 9.250 13.000 9.250 13.000 10.250 17.000 10.250
                 17.000 13.750 13.000 13.750 13.000 14.750 17.000 14.750 17.000 18.250
                 13.000 18.250 13.000 19.250 17.000 19.250 17.000 22.750 13.000 22.750
                 13.000 23.750 17.000 23.750 17.000 27.250 13.000 27.250 13.000 28.250
                 17.000 28.250 17.000 31.750 13.000 31.750 13.000 33.080 17.000 33.080
                 17.000 37.580 12.000 37.580 12.000 4.750 8.000 4.750 8.000 5.750
                 12.000 5.750 12.000 9.250 8.000 9.250 8.000 10.250 12.000 10.250
                 12.000 13.750 8.000 13.750 8.000 14.750 12.000 14.750 12.000 18.250
                 8.000 18.250 8.000 19.250 12.000 19.250 12.000 22.750 8.000 22.750
                 8.000 23.750 12.000 23.750 12.000 27.250 8.000 27.250 8.000 28.250
                 12.000 28.250 12.000 31.750 8.000 31.750 8.000 33.080 12.000 33.080
                 12.000 37.580 7.000 37.580 7.000 4.750 3.000 4.750 3.000 5.750 7.000 5.750
                 7.000 9.250 3.000 9.250 3.000 10.250 7.000 10.250 7.000 13.750
                 3.000 13.750 3.000 14.750 7.000 14.750 7.000 18.250 3.000 18.250
                 3.000 19.250 7.000 19.250 7.000 22.750 3.000 22.750 3.000 23.750
                 7.000 23.750 7.000 27.250 3.000 27.250 3.000 28.250 7.000 28.250
                 7.000 31.750 3.000 31.750 3.000 33.080 7.000 33.080 7.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 18.000 87.170 18.000 88.020
                 20.000 88.020 20.000 91.520 18.000 91.520 18.000 92.370 20.000 92.370
                 20.000 95.870 18.000 95.870 18.000 96.720 20.000 96.720 20.000 100.220
                 18.000 100.220 18.000 101.070 20.000 101.070 20.000 104.570
                 18.000 104.570 18.000 105.420 20.000 105.420 20.000 108.920
                 18.000 108.920 18.000 109.770 20.000 109.770 20.000 113.270
                 18.000 113.270 18.000 114.010 20.000 114.010 20.000 117.510
                 17.000 117.510 17.000 87.170 13.000 87.170 13.000 88.020 17.000 88.020
                 17.000 91.520 13.000 91.520 13.000 92.370 17.000 92.370 17.000 95.870
                 13.000 95.870 13.000 96.720 17.000 96.720 17.000 100.220 13.000 100.220
                 13.000 101.070 17.000 101.070 17.000 104.570 13.000 104.570
                 13.000 105.420 17.000 105.420 17.000 108.920 13.000 108.920
                 13.000 109.770 17.000 109.770 17.000 113.270 13.000 113.270
                 13.000 114.010 17.000 114.010 17.000 117.510 12.000 117.510
                 12.000 87.170 8.000 87.170 8.000 88.020 12.000 88.020 12.000 91.520
                 8.000 91.520 8.000 92.370 12.000 92.370 12.000 95.870 8.000 95.870
                 8.000 96.720 12.000 96.720 12.000 100.220 8.000 100.220 8.000 101.070
                 12.000 101.070 12.000 104.570 8.000 104.570 8.000 105.420 12.000 105.420
                 12.000 108.920 8.000 108.920 8.000 109.770 12.000 109.770 12.000 113.270
                 8.000 113.270 8.000 114.010 12.000 114.010 12.000 117.510 7.000 117.510
                 7.000 87.170 3.000 87.170 3.000 88.020 7.000 88.020 7.000 91.520
                 3.000 91.520 3.000 92.370 7.000 92.370 7.000 95.870 3.000 95.870
                 3.000 96.720 7.000 96.720 7.000 100.220 3.000 100.220 3.000 101.070
                 7.000 101.070 7.000 104.570 3.000 104.570 3.000 105.420 7.000 105.420
                 7.000 108.920 3.000 108.920 3.000 109.770 7.000 109.770 7.000 113.270
                 3.000 113.270 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510
                 0.000 114.010 2.000 114.010 2.000 113.270 0.000 113.270 0.000 109.770
                 2.000 109.770 2.000 108.920 0.000 108.920 0.000 105.420 2.000 105.420
                 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070 2.000 100.220
                 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870 0.000 95.870
                 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520 0.000 88.020
                 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 18.000 87.170 18.000 88.020
                 20.000 88.020 20.000 91.520 18.000 91.520 18.000 92.370 20.000 92.370
                 20.000 95.870 18.000 95.870 18.000 96.720 20.000 96.720 20.000 100.220
                 18.000 100.220 18.000 101.070 20.000 101.070 20.000 104.570
                 18.000 104.570 18.000 105.420 20.000 105.420 20.000 108.920
                 18.000 108.920 18.000 109.770 20.000 109.770 20.000 113.270
                 18.000 113.270 18.000 114.010 20.000 114.010 20.000 117.510
                 17.000 117.510 17.000 87.170 13.000 87.170 13.000 88.020 17.000 88.020
                 17.000 91.520 13.000 91.520 13.000 92.370 17.000 92.370 17.000 95.870
                 13.000 95.870 13.000 96.720 17.000 96.720 17.000 100.220 13.000 100.220
                 13.000 101.070 17.000 101.070 17.000 104.570 13.000 104.570
                 13.000 105.420 17.000 105.420 17.000 108.920 13.000 108.920
                 13.000 109.770 17.000 109.770 17.000 113.270 13.000 113.270
                 13.000 114.010 17.000 114.010 17.000 117.510 12.000 117.510
                 12.000 87.170 8.000 87.170 8.000 88.020 12.000 88.020 12.000 91.520
                 8.000 91.520 8.000 92.370 12.000 92.370 12.000 95.870 8.000 95.870
                 8.000 96.720 12.000 96.720 12.000 100.220 8.000 100.220 8.000 101.070
                 12.000 101.070 12.000 104.570 8.000 104.570 8.000 105.420 12.000 105.420
                 12.000 108.920 8.000 108.920 8.000 109.770 12.000 109.770 12.000 113.270
                 8.000 113.270 8.000 114.010 12.000 114.010 12.000 117.510 7.000 117.510
                 7.000 87.170 3.000 87.170 3.000 88.020 7.000 88.020 7.000 91.520
                 3.000 91.520 3.000 92.370 7.000 92.370 7.000 95.870 3.000 95.870
                 3.000 96.720 7.000 96.720 7.000 100.220 3.000 100.220 3.000 101.070
                 7.000 101.070 7.000 104.570 3.000 104.570 3.000 105.420 7.000 105.420
                 7.000 108.920 3.000 108.920 3.000 109.770 7.000 109.770 7.000 113.270
                 3.000 113.270 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510
                 0.000 114.010 2.000 114.010 2.000 113.270 0.000 113.270 0.000 109.770
                 2.000 109.770 2.000 108.920 0.000 108.920 0.000 105.420 2.000 105.420
                 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070 2.000 100.220
                 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870 0.000 95.870
                 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520 0.000 88.020
                 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 18.000 87.170 18.000 88.020
                 20.000 88.020 20.000 91.520 18.000 91.520 18.000 92.370 20.000 92.370
                 20.000 95.870 18.000 95.870 18.000 96.720 20.000 96.720 20.000 100.220
                 18.000 100.220 18.000 101.070 20.000 101.070 20.000 104.570
                 18.000 104.570 18.000 105.420 20.000 105.420 20.000 108.920
                 18.000 108.920 18.000 109.770 20.000 109.770 20.000 113.270
                 18.000 113.270 18.000 114.010 20.000 114.010 20.000 117.510
                 17.000 117.510 17.000 87.170 13.000 87.170 13.000 88.020 17.000 88.020
                 17.000 91.520 13.000 91.520 13.000 92.370 17.000 92.370 17.000 95.870
                 13.000 95.870 13.000 96.720 17.000 96.720 17.000 100.220 13.000 100.220
                 13.000 101.070 17.000 101.070 17.000 104.570 13.000 104.570
                 13.000 105.420 17.000 105.420 17.000 108.920 13.000 108.920
                 13.000 109.770 17.000 109.770 17.000 113.270 13.000 113.270
                 13.000 114.010 17.000 114.010 17.000 117.510 12.000 117.510
                 12.000 87.170 8.000 87.170 8.000 88.020 12.000 88.020 12.000 91.520
                 8.000 91.520 8.000 92.370 12.000 92.370 12.000 95.870 8.000 95.870
                 8.000 96.720 12.000 96.720 12.000 100.220 8.000 100.220 8.000 101.070
                 12.000 101.070 12.000 104.570 8.000 104.570 8.000 105.420 12.000 105.420
                 12.000 108.920 8.000 108.920 8.000 109.770 12.000 109.770 12.000 113.270
                 8.000 113.270 8.000 114.010 12.000 114.010 12.000 117.510 7.000 117.510
                 7.000 87.170 3.000 87.170 3.000 88.020 7.000 88.020 7.000 91.520
                 3.000 91.520 3.000 92.370 7.000 92.370 7.000 95.870 3.000 95.870
                 3.000 96.720 7.000 96.720 7.000 100.220 3.000 100.220 3.000 101.070
                 7.000 101.070 7.000 104.570 3.000 104.570 3.000 105.420 7.000 105.420
                 7.000 108.920 3.000 108.920 3.000 109.770 7.000 109.770 7.000 113.270
                 3.000 113.270 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510
                 0.000 114.010 2.000 114.010 2.000 113.270 0.000 113.270 0.000 109.770
                 2.000 109.770 2.000 108.920 0.000 108.920 0.000 105.420 2.000 105.420
                 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070 2.000 100.220
                 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870 0.000 95.870
                 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520 0.000 88.020
                 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 18.000 87.170 18.000 88.020
                 20.000 88.020 20.000 91.520 18.000 91.520 18.000 92.370 20.000 92.370
                 20.000 95.870 18.000 95.870 18.000 96.720 20.000 96.720 20.000 100.220
                 18.000 100.220 18.000 101.070 20.000 101.070 20.000 104.570
                 18.000 104.570 18.000 105.420 20.000 105.420 20.000 108.920
                 18.000 108.920 18.000 109.770 20.000 109.770 20.000 113.270
                 18.000 113.270 18.000 114.010 20.000 114.010 20.000 117.510
                 17.000 117.510 17.000 87.170 13.000 87.170 13.000 88.020 17.000 88.020
                 17.000 91.520 13.000 91.520 13.000 92.370 17.000 92.370 17.000 95.870
                 13.000 95.870 13.000 96.720 17.000 96.720 17.000 100.220 13.000 100.220
                 13.000 101.070 17.000 101.070 17.000 104.570 13.000 104.570
                 13.000 105.420 17.000 105.420 17.000 108.920 13.000 108.920
                 13.000 109.770 17.000 109.770 17.000 113.270 13.000 113.270
                 13.000 114.010 17.000 114.010 17.000 117.510 12.000 117.510
                 12.000 87.170 8.000 87.170 8.000 88.020 12.000 88.020 12.000 91.520
                 8.000 91.520 8.000 92.370 12.000 92.370 12.000 95.870 8.000 95.870
                 8.000 96.720 12.000 96.720 12.000 100.220 8.000 100.220 8.000 101.070
                 12.000 101.070 12.000 104.570 8.000 104.570 8.000 105.420 12.000 105.420
                 12.000 108.920 8.000 108.920 8.000 109.770 12.000 109.770 12.000 113.270
                 8.000 113.270 8.000 114.010 12.000 114.010 12.000 117.510 7.000 117.510
                 7.000 87.170 3.000 87.170 3.000 88.020 7.000 88.020 7.000 91.520
                 3.000 91.520 3.000 92.370 7.000 92.370 7.000 95.870 3.000 95.870
                 3.000 96.720 7.000 96.720 7.000 100.220 3.000 100.220 3.000 101.070
                 7.000 101.070 7.000 104.570 3.000 104.570 3.000 105.420 7.000 105.420
                 7.000 108.920 3.000 108.920 3.000 109.770 7.000 109.770 7.000 113.270
                 3.000 113.270 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510
                 0.000 114.010 2.000 114.010 2.000 113.270 0.000 113.270 0.000 109.770
                 2.000 109.770 2.000 108.920 0.000 108.920 0.000 105.420 2.000 105.420
                 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070 2.000 100.220
                 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870 0.000 95.870
                 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520 0.000 88.020
                 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 20.000 83.670 20.000 87.170 18.000 87.170 18.000 88.020
                 20.000 88.020 20.000 91.520 18.000 91.520 18.000 92.370 20.000 92.370
                 20.000 95.870 18.000 95.870 18.000 96.720 20.000 96.720 20.000 100.220
                 18.000 100.220 18.000 101.070 20.000 101.070 20.000 104.570
                 18.000 104.570 18.000 105.420 20.000 105.420 20.000 108.920
                 17.000 108.920 17.000 87.170 13.000 87.170 13.000 88.020 17.000 88.020
                 17.000 91.520 13.000 91.520 13.000 92.370 17.000 92.370 17.000 95.870
                 13.000 95.870 13.000 96.720 17.000 96.720 17.000 100.220 13.000 100.220
                 13.000 101.070 17.000 101.070 17.000 104.570 13.000 104.570
                 13.000 105.420 17.000 105.420 17.000 108.920 12.000 108.920
                 12.000 87.170 8.000 87.170 8.000 88.020 12.000 88.020 12.000 91.520
                 8.000 91.520 8.000 92.370 12.000 92.370 12.000 95.870 8.000 95.870
                 8.000 96.720 12.000 96.720 12.000 100.220 8.000 100.220 8.000 101.070
                 12.000 101.070 12.000 104.570 8.000 104.570 8.000 105.420 12.000 105.420
                 12.000 108.920 7.000 108.920 7.000 87.170 3.000 87.170 3.000 88.020
                 7.000 88.020 7.000 91.520 3.000 91.520 3.000 92.370 7.000 92.370
                 7.000 95.870 3.000 95.870 3.000 96.720 7.000 96.720 7.000 100.220
                 3.000 100.220 3.000 101.070 7.000 101.070 7.000 104.570 3.000 104.570
                 3.000 105.420 7.000 105.420 7.000 108.920 0.000 108.920 0.000 105.420
                 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070
                 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870
                 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520
                 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        END
    END VSS
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 20.000 109.770 20.000 113.270 18.000 113.270
                 18.000 114.010 20.000 114.010 20.000 117.510 17.000 117.510
                 17.000 113.270 13.000 113.270 13.000 114.010 17.000 114.010
                 17.000 117.510 12.000 117.510 12.000 113.270 8.000 113.270 8.000 114.010
                 12.000 114.010 12.000 117.510 7.000 117.510 7.000 113.270 3.000 113.270
                 3.000 114.010 7.000 114.010 7.000 117.510 0.000 117.510 0.000 114.010
                 2.000 114.010 2.000 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 20.000 118.500 ;
        END
    END POC
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 18.000 44.475 18.000 45.475
                 20.000 45.475 20.000 48.975 18.000 48.975 18.000 49.975 20.000 49.975
                 20.000 53.475 18.000 53.475 18.000 54.475 20.000 54.475 20.000 57.975
                 18.000 57.975 18.000 58.975 20.000 58.975 20.000 62.475 18.000 62.475
                 18.000 63.475 20.000 63.475 20.000 66.975 18.000 66.975 18.000 67.975
                 20.000 67.975 20.000 71.475 18.000 71.475 18.000 72.475 20.000 72.475
                 20.000 75.975 17.000 75.975 17.000 44.475 13.000 44.475 13.000 45.475
                 17.000 45.475 17.000 48.975 13.000 48.975 13.000 49.975 17.000 49.975
                 17.000 53.475 13.000 53.475 13.000 54.475 17.000 54.475 17.000 57.975
                 13.000 57.975 13.000 58.975 17.000 58.975 17.000 62.475 13.000 62.475
                 13.000 63.475 17.000 63.475 17.000 66.975 13.000 66.975 13.000 67.975
                 17.000 67.975 17.000 71.475 13.000 71.475 13.000 72.475 17.000 72.475
                 17.000 75.975 12.000 75.975 12.000 44.475 8.000 44.475 8.000 45.475
                 12.000 45.475 12.000 48.975 8.000 48.975 8.000 49.975 12.000 49.975
                 12.000 53.475 8.000 53.475 8.000 54.475 12.000 54.475 12.000 57.975
                 8.000 57.975 8.000 58.975 12.000 58.975 12.000 62.475 8.000 62.475
                 8.000 63.475 12.000 63.475 12.000 66.975 8.000 66.975 8.000 67.975
                 12.000 67.975 12.000 71.475 8.000 71.475 8.000 72.475 12.000 72.475
                 12.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 18.000 44.475 18.000 45.475
                 20.000 45.475 20.000 48.975 18.000 48.975 18.000 49.975 20.000 49.975
                 20.000 53.475 18.000 53.475 18.000 54.475 20.000 54.475 20.000 57.975
                 18.000 57.975 18.000 58.975 20.000 58.975 20.000 62.475 18.000 62.475
                 18.000 63.475 20.000 63.475 20.000 66.975 18.000 66.975 18.000 67.975
                 20.000 67.975 20.000 71.475 18.000 71.475 18.000 72.475 20.000 72.475
                 20.000 75.975 17.000 75.975 17.000 44.475 13.000 44.475 13.000 45.475
                 17.000 45.475 17.000 48.975 13.000 48.975 13.000 49.975 17.000 49.975
                 17.000 53.475 13.000 53.475 13.000 54.475 17.000 54.475 17.000 57.975
                 13.000 57.975 13.000 58.975 17.000 58.975 17.000 62.475 13.000 62.475
                 13.000 63.475 17.000 63.475 17.000 66.975 13.000 66.975 13.000 67.975
                 17.000 67.975 17.000 71.475 13.000 71.475 13.000 72.475 17.000 72.475
                 17.000 75.975 12.000 75.975 12.000 44.475 8.000 44.475 8.000 45.475
                 12.000 45.475 12.000 48.975 8.000 48.975 8.000 49.975 12.000 49.975
                 12.000 53.475 8.000 53.475 8.000 54.475 12.000 54.475 12.000 57.975
                 8.000 57.975 8.000 58.975 12.000 58.975 12.000 62.475 8.000 62.475
                 8.000 63.475 12.000 63.475 12.000 66.975 8.000 66.975 8.000 67.975
                 12.000 67.975 12.000 71.475 8.000 71.475 8.000 72.475 12.000 72.475
                 12.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 18.000 44.475 18.000 45.475
                 20.000 45.475 20.000 48.975 18.000 48.975 18.000 49.975 20.000 49.975
                 20.000 53.475 18.000 53.475 18.000 54.475 20.000 54.475 20.000 57.975
                 18.000 57.975 18.000 58.975 20.000 58.975 20.000 62.475 18.000 62.475
                 18.000 63.475 20.000 63.475 20.000 66.975 18.000 66.975 18.000 67.975
                 20.000 67.975 20.000 71.475 18.000 71.475 18.000 72.475 20.000 72.475
                 20.000 75.975 17.000 75.975 17.000 44.475 13.000 44.475 13.000 45.475
                 17.000 45.475 17.000 48.975 13.000 48.975 13.000 49.975 17.000 49.975
                 17.000 53.475 13.000 53.475 13.000 54.475 17.000 54.475 17.000 57.975
                 13.000 57.975 13.000 58.975 17.000 58.975 17.000 62.475 13.000 62.475
                 13.000 63.475 17.000 63.475 17.000 66.975 13.000 66.975 13.000 67.975
                 17.000 67.975 17.000 71.475 13.000 71.475 13.000 72.475 17.000 72.475
                 17.000 75.975 12.000 75.975 12.000 44.475 8.000 44.475 8.000 45.475
                 12.000 45.475 12.000 48.975 8.000 48.975 8.000 49.975 12.000 49.975
                 12.000 53.475 8.000 53.475 8.000 54.475 12.000 54.475 12.000 57.975
                 8.000 57.975 8.000 58.975 12.000 58.975 12.000 62.475 8.000 62.475
                 8.000 63.475 12.000 63.475 12.000 66.975 8.000 66.975 8.000 67.975
                 12.000 67.975 12.000 71.475 8.000 71.475 8.000 72.475 12.000 72.475
                 12.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 18.000 44.475 18.000 45.475
                 20.000 45.475 20.000 48.975 18.000 48.975 18.000 49.975 20.000 49.975
                 20.000 53.475 18.000 53.475 18.000 54.475 20.000 54.475 20.000 57.975
                 18.000 57.975 18.000 58.975 20.000 58.975 20.000 62.475 18.000 62.475
                 18.000 63.475 20.000 63.475 20.000 66.975 18.000 66.975 18.000 67.975
                 20.000 67.975 20.000 71.475 18.000 71.475 18.000 72.475 20.000 72.475
                 20.000 75.975 17.000 75.975 17.000 44.475 13.000 44.475 13.000 45.475
                 17.000 45.475 17.000 48.975 13.000 48.975 13.000 49.975 17.000 49.975
                 17.000 53.475 13.000 53.475 13.000 54.475 17.000 54.475 17.000 57.975
                 13.000 57.975 13.000 58.975 17.000 58.975 17.000 62.475 13.000 62.475
                 13.000 63.475 17.000 63.475 17.000 66.975 13.000 66.975 13.000 67.975
                 17.000 67.975 17.000 71.475 13.000 71.475 13.000 72.475 17.000 72.475
                 17.000 75.975 12.000 75.975 12.000 44.475 8.000 44.475 8.000 45.475
                 12.000 45.475 12.000 48.975 8.000 48.975 8.000 49.975 12.000 49.975
                 12.000 53.475 8.000 53.475 8.000 54.475 12.000 54.475 12.000 57.975
                 8.000 57.975 8.000 58.975 12.000 58.975 12.000 62.475 8.000 62.475
                 8.000 63.475 12.000 63.475 12.000 66.975 8.000 66.975 8.000 67.975
                 12.000 67.975 12.000 71.475 8.000 71.475 8.000 72.475 12.000 72.475
                 12.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 20.000 82.975 ;
                POLYGON  0.000 40.975 20.000 40.975 20.000 44.475 18.000 44.475 18.000 45.475
                 20.000 45.475 20.000 48.975 18.000 48.975 18.000 49.975 20.000 49.975
                 20.000 53.475 18.000 53.475 18.000 54.475 20.000 54.475 20.000 57.975
                 18.000 57.975 18.000 58.975 20.000 58.975 20.000 62.475 18.000 62.475
                 18.000 63.475 20.000 63.475 20.000 66.975 18.000 66.975 18.000 67.975
                 20.000 67.975 20.000 71.475 18.000 71.475 18.000 72.475 20.000 72.475
                 20.000 75.975 17.000 75.975 17.000 44.475 13.000 44.475 13.000 45.475
                 17.000 45.475 17.000 48.975 13.000 48.975 13.000 49.975 17.000 49.975
                 17.000 53.475 13.000 53.475 13.000 54.475 17.000 54.475 17.000 57.975
                 13.000 57.975 13.000 58.975 17.000 58.975 17.000 62.475 13.000 62.475
                 13.000 63.475 17.000 63.475 17.000 66.975 13.000 66.975 13.000 67.975
                 17.000 67.975 17.000 71.475 13.000 71.475 13.000 72.475 17.000 72.475
                 17.000 75.975 12.000 75.975 12.000 44.475 8.000 44.475 8.000 45.475
                 12.000 45.475 12.000 48.975 8.000 48.975 8.000 49.975 12.000 49.975
                 12.000 53.475 8.000 53.475 8.000 54.475 12.000 54.475 12.000 57.975
                 8.000 57.975 8.000 58.975 12.000 58.975 12.000 62.475 8.000 62.475
                 8.000 63.475 12.000 63.475 12.000 66.975 8.000 66.975 8.000 67.975
                 12.000 67.975 12.000 71.475 8.000 71.475 8.000 72.475 12.000 72.475
                 12.000 75.975 7.000 75.975 7.000 44.475 3.000 44.475 3.000 45.475
                 7.000 45.475 7.000 48.975 3.000 48.975 3.000 49.975 7.000 49.975
                 7.000 53.475 3.000 53.475 3.000 54.475 7.000 54.475 7.000 57.975
                 3.000 57.975 3.000 58.975 7.000 58.975 7.000 62.475 3.000 62.475
                 3.000 63.475 7.000 63.475 7.000 66.975 3.000 66.975 3.000 67.975
                 7.000 67.975 7.000 71.475 3.000 71.475 3.000 72.475 7.000 72.475
                 7.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        END
    END VDDPST
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA2 ;
        RECT  18.000 1.250 20.000 4.750 ;
        RECT  18.000 5.750 20.000 9.250 ;
        RECT  18.000 10.250 20.000 13.750 ;
        RECT  18.000 14.750 20.000 18.250 ;
        RECT  18.000 19.250 20.000 22.750 ;
        RECT  18.000 23.750 20.000 27.250 ;
        RECT  18.000 28.250 20.000 31.750 ;
        RECT  18.000 33.080 20.000 37.580 ;
        RECT  18.000 40.975 20.000 44.475 ;
        RECT  18.000 45.475 20.000 48.975 ;
        RECT  18.000 49.975 20.000 53.475 ;
        RECT  18.000 54.475 20.000 57.975 ;
        RECT  18.000 58.975 20.000 62.475 ;
        RECT  18.000 63.475 20.000 66.975 ;
        RECT  18.000 67.975 20.000 71.475 ;
        RECT  18.000 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  18.000 83.670 20.000 87.170 ;
        RECT  18.000 88.020 20.000 91.520 ;
        RECT  18.000 92.370 20.000 95.870 ;
        RECT  18.000 96.720 20.000 100.220 ;
        RECT  18.000 101.070 20.000 104.570 ;
        RECT  18.000 105.420 20.000 108.920 ;
        RECT  18.000 109.770 20.000 113.270 ;
        RECT  18.000 114.010 20.000 117.510 ;
        RECT  17.000 1.250 18.000 37.580 ;
        RECT  17.000 40.975 18.000 75.975 ;
        RECT  17.000 83.670 18.000 108.920 ;
        RECT  17.000 109.770 18.000 117.510 ;
        RECT  13.000 1.250 17.000 4.750 ;
        RECT  13.000 5.750 17.000 9.250 ;
        RECT  13.000 10.250 17.000 13.750 ;
        RECT  13.000 14.750 17.000 18.250 ;
        RECT  13.000 19.250 17.000 22.750 ;
        RECT  13.000 23.750 17.000 27.250 ;
        RECT  13.000 28.250 17.000 31.750 ;
        RECT  13.000 33.080 17.000 37.580 ;
        RECT  13.000 40.975 17.000 44.475 ;
        RECT  13.000 45.475 17.000 48.975 ;
        RECT  13.000 49.975 17.000 53.475 ;
        RECT  13.000 54.475 17.000 57.975 ;
        RECT  13.000 58.975 17.000 62.475 ;
        RECT  13.000 63.475 17.000 66.975 ;
        RECT  13.000 67.975 17.000 71.475 ;
        RECT  13.000 72.475 17.000 75.975 ;
        RECT  13.000 83.670 17.000 87.170 ;
        RECT  13.000 88.020 17.000 91.520 ;
        RECT  13.000 92.370 17.000 95.870 ;
        RECT  13.000 96.720 17.000 100.220 ;
        RECT  13.000 101.070 17.000 104.570 ;
        RECT  13.000 105.420 17.000 108.920 ;
        RECT  13.000 109.770 17.000 113.270 ;
        RECT  13.000 114.010 17.000 117.510 ;
        RECT  12.000 1.250 13.000 37.580 ;
        RECT  12.000 40.975 13.000 75.975 ;
        RECT  12.000 83.670 13.000 108.920 ;
        RECT  12.000 109.770 13.000 117.510 ;
        RECT  8.000 1.250 12.000 4.750 ;
        RECT  8.000 5.750 12.000 9.250 ;
        RECT  8.000 10.250 12.000 13.750 ;
        RECT  8.000 14.750 12.000 18.250 ;
        RECT  8.000 19.250 12.000 22.750 ;
        RECT  8.000 23.750 12.000 27.250 ;
        RECT  8.000 28.250 12.000 31.750 ;
        RECT  8.000 33.080 12.000 37.580 ;
        RECT  8.000 40.975 12.000 44.475 ;
        RECT  8.000 45.475 12.000 48.975 ;
        RECT  8.000 49.975 12.000 53.475 ;
        RECT  8.000 54.475 12.000 57.975 ;
        RECT  8.000 58.975 12.000 62.475 ;
        RECT  8.000 63.475 12.000 66.975 ;
        RECT  8.000 67.975 12.000 71.475 ;
        RECT  8.000 72.475 12.000 75.975 ;
        RECT  8.000 83.670 12.000 87.170 ;
        RECT  8.000 88.020 12.000 91.520 ;
        RECT  8.000 92.370 12.000 95.870 ;
        RECT  8.000 96.720 12.000 100.220 ;
        RECT  8.000 101.070 12.000 104.570 ;
        RECT  8.000 105.420 12.000 108.920 ;
        RECT  8.000 109.770 12.000 113.270 ;
        RECT  8.000 114.010 12.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 108.920 ;
        RECT  7.000 109.770 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 108.920 ;
        RECT  2.000 109.770 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA3 ;
        RECT  18.000 1.250 20.000 4.750 ;
        RECT  18.000 5.750 20.000 9.250 ;
        RECT  18.000 10.250 20.000 13.750 ;
        RECT  18.000 14.750 20.000 18.250 ;
        RECT  18.000 19.250 20.000 22.750 ;
        RECT  18.000 23.750 20.000 27.250 ;
        RECT  18.000 28.250 20.000 31.750 ;
        RECT  18.000 33.080 20.000 37.580 ;
        RECT  18.000 40.975 20.000 44.475 ;
        RECT  18.000 45.475 20.000 48.975 ;
        RECT  18.000 49.975 20.000 53.475 ;
        RECT  18.000 54.475 20.000 57.975 ;
        RECT  18.000 58.975 20.000 62.475 ;
        RECT  18.000 63.475 20.000 66.975 ;
        RECT  18.000 67.975 20.000 71.475 ;
        RECT  18.000 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  18.000 83.670 20.000 87.170 ;
        RECT  18.000 88.020 20.000 91.520 ;
        RECT  18.000 92.370 20.000 95.870 ;
        RECT  18.000 96.720 20.000 100.220 ;
        RECT  18.000 101.070 20.000 104.570 ;
        RECT  18.000 105.420 20.000 108.920 ;
        RECT  18.000 109.770 20.000 113.270 ;
        RECT  18.000 114.010 20.000 117.510 ;
        RECT  17.000 1.250 18.000 37.580 ;
        RECT  17.000 40.975 18.000 75.975 ;
        RECT  17.000 83.670 18.000 117.510 ;
        RECT  13.000 1.250 17.000 4.750 ;
        RECT  13.000 5.750 17.000 9.250 ;
        RECT  13.000 10.250 17.000 13.750 ;
        RECT  13.000 14.750 17.000 18.250 ;
        RECT  13.000 19.250 17.000 22.750 ;
        RECT  13.000 23.750 17.000 27.250 ;
        RECT  13.000 28.250 17.000 31.750 ;
        RECT  13.000 33.080 17.000 37.580 ;
        RECT  13.000 40.975 17.000 44.475 ;
        RECT  13.000 45.475 17.000 48.975 ;
        RECT  13.000 49.975 17.000 53.475 ;
        RECT  13.000 54.475 17.000 57.975 ;
        RECT  13.000 58.975 17.000 62.475 ;
        RECT  13.000 63.475 17.000 66.975 ;
        RECT  13.000 67.975 17.000 71.475 ;
        RECT  13.000 72.475 17.000 75.975 ;
        RECT  13.000 83.670 17.000 87.170 ;
        RECT  13.000 88.020 17.000 91.520 ;
        RECT  13.000 92.370 17.000 95.870 ;
        RECT  13.000 96.720 17.000 100.220 ;
        RECT  13.000 101.070 17.000 104.570 ;
        RECT  13.000 105.420 17.000 108.920 ;
        RECT  13.000 109.770 17.000 113.270 ;
        RECT  13.000 114.010 17.000 117.510 ;
        RECT  12.000 1.250 13.000 37.580 ;
        RECT  12.000 40.975 13.000 75.975 ;
        RECT  12.000 83.670 13.000 117.510 ;
        RECT  8.000 1.250 12.000 4.750 ;
        RECT  8.000 5.750 12.000 9.250 ;
        RECT  8.000 10.250 12.000 13.750 ;
        RECT  8.000 14.750 12.000 18.250 ;
        RECT  8.000 19.250 12.000 22.750 ;
        RECT  8.000 23.750 12.000 27.250 ;
        RECT  8.000 28.250 12.000 31.750 ;
        RECT  8.000 33.080 12.000 37.580 ;
        RECT  8.000 40.975 12.000 44.475 ;
        RECT  8.000 45.475 12.000 48.975 ;
        RECT  8.000 49.975 12.000 53.475 ;
        RECT  8.000 54.475 12.000 57.975 ;
        RECT  8.000 58.975 12.000 62.475 ;
        RECT  8.000 63.475 12.000 66.975 ;
        RECT  8.000 67.975 12.000 71.475 ;
        RECT  8.000 72.475 12.000 75.975 ;
        RECT  8.000 83.670 12.000 87.170 ;
        RECT  8.000 88.020 12.000 91.520 ;
        RECT  8.000 92.370 12.000 95.870 ;
        RECT  8.000 96.720 12.000 100.220 ;
        RECT  8.000 101.070 12.000 104.570 ;
        RECT  8.000 105.420 12.000 108.920 ;
        RECT  8.000 109.770 12.000 113.270 ;
        RECT  8.000 114.010 12.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA4 ;
        RECT  18.000 1.250 20.000 4.750 ;
        RECT  18.000 5.750 20.000 9.250 ;
        RECT  18.000 10.250 20.000 13.750 ;
        RECT  18.000 14.750 20.000 18.250 ;
        RECT  18.000 19.250 20.000 22.750 ;
        RECT  18.000 23.750 20.000 27.250 ;
        RECT  18.000 28.250 20.000 31.750 ;
        RECT  18.000 33.080 20.000 37.580 ;
        RECT  18.000 40.975 20.000 44.475 ;
        RECT  18.000 45.475 20.000 48.975 ;
        RECT  18.000 49.975 20.000 53.475 ;
        RECT  18.000 54.475 20.000 57.975 ;
        RECT  18.000 58.975 20.000 62.475 ;
        RECT  18.000 63.475 20.000 66.975 ;
        RECT  18.000 67.975 20.000 71.475 ;
        RECT  18.000 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  18.000 83.670 20.000 87.170 ;
        RECT  18.000 88.020 20.000 91.520 ;
        RECT  18.000 92.370 20.000 95.870 ;
        RECT  18.000 96.720 20.000 100.220 ;
        RECT  18.000 101.070 20.000 104.570 ;
        RECT  18.000 105.420 20.000 108.920 ;
        RECT  18.000 109.770 20.000 113.270 ;
        RECT  18.000 114.010 20.000 117.510 ;
        RECT  17.000 1.250 18.000 37.580 ;
        RECT  17.000 40.975 18.000 75.975 ;
        RECT  17.000 83.670 18.000 117.510 ;
        RECT  13.000 1.250 17.000 4.750 ;
        RECT  13.000 5.750 17.000 9.250 ;
        RECT  13.000 10.250 17.000 13.750 ;
        RECT  13.000 14.750 17.000 18.250 ;
        RECT  13.000 19.250 17.000 22.750 ;
        RECT  13.000 23.750 17.000 27.250 ;
        RECT  13.000 28.250 17.000 31.750 ;
        RECT  13.000 33.080 17.000 37.580 ;
        RECT  13.000 40.975 17.000 44.475 ;
        RECT  13.000 45.475 17.000 48.975 ;
        RECT  13.000 49.975 17.000 53.475 ;
        RECT  13.000 54.475 17.000 57.975 ;
        RECT  13.000 58.975 17.000 62.475 ;
        RECT  13.000 63.475 17.000 66.975 ;
        RECT  13.000 67.975 17.000 71.475 ;
        RECT  13.000 72.475 17.000 75.975 ;
        RECT  13.000 83.670 17.000 87.170 ;
        RECT  13.000 88.020 17.000 91.520 ;
        RECT  13.000 92.370 17.000 95.870 ;
        RECT  13.000 96.720 17.000 100.220 ;
        RECT  13.000 101.070 17.000 104.570 ;
        RECT  13.000 105.420 17.000 108.920 ;
        RECT  13.000 109.770 17.000 113.270 ;
        RECT  13.000 114.010 17.000 117.510 ;
        RECT  12.000 1.250 13.000 37.580 ;
        RECT  12.000 40.975 13.000 75.975 ;
        RECT  12.000 83.670 13.000 117.510 ;
        RECT  8.000 1.250 12.000 4.750 ;
        RECT  8.000 5.750 12.000 9.250 ;
        RECT  8.000 10.250 12.000 13.750 ;
        RECT  8.000 14.750 12.000 18.250 ;
        RECT  8.000 19.250 12.000 22.750 ;
        RECT  8.000 23.750 12.000 27.250 ;
        RECT  8.000 28.250 12.000 31.750 ;
        RECT  8.000 33.080 12.000 37.580 ;
        RECT  8.000 40.975 12.000 44.475 ;
        RECT  8.000 45.475 12.000 48.975 ;
        RECT  8.000 49.975 12.000 53.475 ;
        RECT  8.000 54.475 12.000 57.975 ;
        RECT  8.000 58.975 12.000 62.475 ;
        RECT  8.000 63.475 12.000 66.975 ;
        RECT  8.000 67.975 12.000 71.475 ;
        RECT  8.000 72.475 12.000 75.975 ;
        RECT  8.000 83.670 12.000 87.170 ;
        RECT  8.000 88.020 12.000 91.520 ;
        RECT  8.000 92.370 12.000 95.870 ;
        RECT  8.000 96.720 12.000 100.220 ;
        RECT  8.000 101.070 12.000 104.570 ;
        RECT  8.000 105.420 12.000 108.920 ;
        RECT  8.000 109.770 12.000 113.270 ;
        RECT  8.000 114.010 12.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA5 ;
        RECT  18.000 1.250 20.000 4.750 ;
        RECT  18.000 5.750 20.000 9.250 ;
        RECT  18.000 10.250 20.000 13.750 ;
        RECT  18.000 14.750 20.000 18.250 ;
        RECT  18.000 19.250 20.000 22.750 ;
        RECT  18.000 23.750 20.000 27.250 ;
        RECT  18.000 28.250 20.000 31.750 ;
        RECT  18.000 33.080 20.000 37.580 ;
        RECT  18.000 40.975 20.000 44.475 ;
        RECT  18.000 45.475 20.000 48.975 ;
        RECT  18.000 49.975 20.000 53.475 ;
        RECT  18.000 54.475 20.000 57.975 ;
        RECT  18.000 58.975 20.000 62.475 ;
        RECT  18.000 63.475 20.000 66.975 ;
        RECT  18.000 67.975 20.000 71.475 ;
        RECT  18.000 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  18.000 83.670 20.000 87.170 ;
        RECT  18.000 88.020 20.000 91.520 ;
        RECT  18.000 92.370 20.000 95.870 ;
        RECT  18.000 96.720 20.000 100.220 ;
        RECT  18.000 101.070 20.000 104.570 ;
        RECT  18.000 105.420 20.000 108.920 ;
        RECT  18.000 109.770 20.000 113.270 ;
        RECT  18.000 114.010 20.000 117.510 ;
        RECT  17.000 1.250 18.000 37.580 ;
        RECT  17.000 40.975 18.000 75.975 ;
        RECT  17.000 83.670 18.000 117.510 ;
        RECT  13.000 1.250 17.000 4.750 ;
        RECT  13.000 5.750 17.000 9.250 ;
        RECT  13.000 10.250 17.000 13.750 ;
        RECT  13.000 14.750 17.000 18.250 ;
        RECT  13.000 19.250 17.000 22.750 ;
        RECT  13.000 23.750 17.000 27.250 ;
        RECT  13.000 28.250 17.000 31.750 ;
        RECT  13.000 33.080 17.000 37.580 ;
        RECT  13.000 40.975 17.000 44.475 ;
        RECT  13.000 45.475 17.000 48.975 ;
        RECT  13.000 49.975 17.000 53.475 ;
        RECT  13.000 54.475 17.000 57.975 ;
        RECT  13.000 58.975 17.000 62.475 ;
        RECT  13.000 63.475 17.000 66.975 ;
        RECT  13.000 67.975 17.000 71.475 ;
        RECT  13.000 72.475 17.000 75.975 ;
        RECT  13.000 83.670 17.000 87.170 ;
        RECT  13.000 88.020 17.000 91.520 ;
        RECT  13.000 92.370 17.000 95.870 ;
        RECT  13.000 96.720 17.000 100.220 ;
        RECT  13.000 101.070 17.000 104.570 ;
        RECT  13.000 105.420 17.000 108.920 ;
        RECT  13.000 109.770 17.000 113.270 ;
        RECT  13.000 114.010 17.000 117.510 ;
        RECT  12.000 1.250 13.000 37.580 ;
        RECT  12.000 40.975 13.000 75.975 ;
        RECT  12.000 83.670 13.000 117.510 ;
        RECT  8.000 1.250 12.000 4.750 ;
        RECT  8.000 5.750 12.000 9.250 ;
        RECT  8.000 10.250 12.000 13.750 ;
        RECT  8.000 14.750 12.000 18.250 ;
        RECT  8.000 19.250 12.000 22.750 ;
        RECT  8.000 23.750 12.000 27.250 ;
        RECT  8.000 28.250 12.000 31.750 ;
        RECT  8.000 33.080 12.000 37.580 ;
        RECT  8.000 40.975 12.000 44.475 ;
        RECT  8.000 45.475 12.000 48.975 ;
        RECT  8.000 49.975 12.000 53.475 ;
        RECT  8.000 54.475 12.000 57.975 ;
        RECT  8.000 58.975 12.000 62.475 ;
        RECT  8.000 63.475 12.000 66.975 ;
        RECT  8.000 67.975 12.000 71.475 ;
        RECT  8.000 72.475 12.000 75.975 ;
        RECT  8.000 83.670 12.000 87.170 ;
        RECT  8.000 88.020 12.000 91.520 ;
        RECT  8.000 92.370 12.000 95.870 ;
        RECT  8.000 96.720 12.000 100.220 ;
        RECT  8.000 101.070 12.000 104.570 ;
        RECT  8.000 105.420 12.000 108.920 ;
        RECT  8.000 109.770 12.000 113.270 ;
        RECT  8.000 114.010 12.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 20.000 120.000 ;
        LAYER VIA6 ;
        RECT  18.000 1.250 20.000 4.750 ;
        RECT  18.000 5.750 20.000 9.250 ;
        RECT  18.000 10.250 20.000 13.750 ;
        RECT  18.000 14.750 20.000 18.250 ;
        RECT  18.000 19.250 20.000 22.750 ;
        RECT  18.000 23.750 20.000 27.250 ;
        RECT  18.000 28.250 20.000 31.750 ;
        RECT  18.000 33.080 20.000 37.580 ;
        RECT  18.000 40.975 20.000 44.475 ;
        RECT  18.000 45.475 20.000 48.975 ;
        RECT  18.000 49.975 20.000 53.475 ;
        RECT  18.000 54.475 20.000 57.975 ;
        RECT  18.000 58.975 20.000 62.475 ;
        RECT  18.000 63.475 20.000 66.975 ;
        RECT  18.000 67.975 20.000 71.475 ;
        RECT  18.000 72.475 20.000 75.975 ;
        RECT  0.000 79.975 20.000 82.975 ;
        RECT  18.000 83.670 20.000 87.170 ;
        RECT  18.000 88.020 20.000 91.520 ;
        RECT  18.000 92.370 20.000 95.870 ;
        RECT  18.000 96.720 20.000 100.220 ;
        RECT  18.000 101.070 20.000 104.570 ;
        RECT  18.000 105.420 20.000 108.920 ;
        RECT  18.000 109.770 20.000 113.270 ;
        RECT  18.000 114.010 20.000 117.510 ;
        RECT  17.000 1.250 18.000 37.580 ;
        RECT  17.000 40.975 18.000 75.975 ;
        RECT  17.000 83.670 18.000 117.510 ;
        RECT  13.000 1.250 17.000 4.750 ;
        RECT  13.000 5.750 17.000 9.250 ;
        RECT  13.000 10.250 17.000 13.750 ;
        RECT  13.000 14.750 17.000 18.250 ;
        RECT  13.000 19.250 17.000 22.750 ;
        RECT  13.000 23.750 17.000 27.250 ;
        RECT  13.000 28.250 17.000 31.750 ;
        RECT  13.000 33.080 17.000 37.580 ;
        RECT  13.000 40.975 17.000 44.475 ;
        RECT  13.000 45.475 17.000 48.975 ;
        RECT  13.000 49.975 17.000 53.475 ;
        RECT  13.000 54.475 17.000 57.975 ;
        RECT  13.000 58.975 17.000 62.475 ;
        RECT  13.000 63.475 17.000 66.975 ;
        RECT  13.000 67.975 17.000 71.475 ;
        RECT  13.000 72.475 17.000 75.975 ;
        RECT  13.000 83.670 17.000 87.170 ;
        RECT  13.000 88.020 17.000 91.520 ;
        RECT  13.000 92.370 17.000 95.870 ;
        RECT  13.000 96.720 17.000 100.220 ;
        RECT  13.000 101.070 17.000 104.570 ;
        RECT  13.000 105.420 17.000 108.920 ;
        RECT  13.000 109.770 17.000 113.270 ;
        RECT  13.000 114.010 17.000 117.510 ;
        RECT  12.000 1.250 13.000 37.580 ;
        RECT  12.000 40.975 13.000 75.975 ;
        RECT  12.000 83.670 13.000 117.510 ;
        RECT  8.000 1.250 12.000 4.750 ;
        RECT  8.000 5.750 12.000 9.250 ;
        RECT  8.000 10.250 12.000 13.750 ;
        RECT  8.000 14.750 12.000 18.250 ;
        RECT  8.000 19.250 12.000 22.750 ;
        RECT  8.000 23.750 12.000 27.250 ;
        RECT  8.000 28.250 12.000 31.750 ;
        RECT  8.000 33.080 12.000 37.580 ;
        RECT  8.000 40.975 12.000 44.475 ;
        RECT  8.000 45.475 12.000 48.975 ;
        RECT  8.000 49.975 12.000 53.475 ;
        RECT  8.000 54.475 12.000 57.975 ;
        RECT  8.000 58.975 12.000 62.475 ;
        RECT  8.000 63.475 12.000 66.975 ;
        RECT  8.000 67.975 12.000 71.475 ;
        RECT  8.000 72.475 12.000 75.975 ;
        RECT  8.000 83.670 12.000 87.170 ;
        RECT  8.000 88.020 12.000 91.520 ;
        RECT  8.000 92.370 12.000 95.870 ;
        RECT  8.000 96.720 12.000 100.220 ;
        RECT  8.000 101.070 12.000 104.570 ;
        RECT  8.000 105.420 12.000 108.920 ;
        RECT  8.000 109.770 12.000 113.270 ;
        RECT  8.000 114.010 12.000 117.510 ;
        RECT  7.000 1.250 8.000 37.580 ;
        RECT  7.000 40.975 8.000 75.975 ;
        RECT  7.000 83.670 8.000 117.510 ;
        RECT  3.000 1.250 7.000 4.750 ;
        RECT  3.000 5.750 7.000 9.250 ;
        RECT  3.000 10.250 7.000 13.750 ;
        RECT  3.000 14.750 7.000 18.250 ;
        RECT  3.000 19.250 7.000 22.750 ;
        RECT  3.000 23.750 7.000 27.250 ;
        RECT  3.000 28.250 7.000 31.750 ;
        RECT  3.000 33.080 7.000 37.580 ;
        RECT  3.000 40.975 7.000 44.475 ;
        RECT  3.000 45.475 7.000 48.975 ;
        RECT  3.000 49.975 7.000 53.475 ;
        RECT  3.000 54.475 7.000 57.975 ;
        RECT  3.000 58.975 7.000 62.475 ;
        RECT  3.000 63.475 7.000 66.975 ;
        RECT  3.000 67.975 7.000 71.475 ;
        RECT  3.000 72.475 7.000 75.975 ;
        RECT  3.000 83.670 7.000 87.170 ;
        RECT  3.000 88.020 7.000 91.520 ;
        RECT  3.000 92.370 7.000 95.870 ;
        RECT  3.000 96.720 7.000 100.220 ;
        RECT  3.000 101.070 7.000 104.570 ;
        RECT  3.000 105.420 7.000 108.920 ;
        RECT  3.000 109.770 7.000 113.270 ;
        RECT  3.000 114.010 7.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 20.000 120.000 ;
    END
END PFILLER20_G

MACRO PFILLER5A_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER5A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        LAYER M6 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        LAYER M5 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        LAYER M4 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        LAYER M3 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        LAYER M6 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        LAYER M5 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        LAYER M4 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        LAYER M3 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 1.250 5.000 5.750 ;
        RECT  0.000 7.250 5.000 11.750 ;
        RECT  0.000 13.250 5.000 17.750 ;
        RECT  0.000 19.250 5.000 23.750 ;
        RECT  0.000 25.250 5.000 29.750 ;
        RECT  0.000 31.250 5.000 35.750 ;
        RECT  0.000 36.750 5.000 39.290 ;
        RECT  0.000 40.975 5.000 44.475 ;
        RECT  0.000 45.475 5.000 48.975 ;
        RECT  0.000 49.975 5.000 53.475 ;
        RECT  0.000 54.475 5.000 57.975 ;
        RECT  0.000 58.975 5.000 62.475 ;
        RECT  0.000 63.475 5.000 66.975 ;
        RECT  0.000 67.975 5.000 71.475 ;
        RECT  0.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  0.000 83.670 5.000 87.170 ;
        RECT  0.000 88.020 5.000 91.520 ;
        RECT  0.000 92.370 5.000 95.870 ;
        RECT  0.000 96.720 5.000 100.220 ;
        RECT  0.000 101.070 5.000 104.570 ;
        RECT  0.000 105.420 5.000 108.920 ;
        RECT  0.000 109.770 5.000 113.270 ;
        RECT  0.000 114.010 5.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 5.000 120.000 ;
    END
END PFILLER5A_G

MACRO PFILLER5_G
    CLASS PAD SPACER ;
    FOREIGN PFILLER5_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 5.000 1.250 5.000 4.750 3.000 4.750 3.000 5.750 5.000 5.750
                 5.000 9.250 3.000 9.250 3.000 10.250 5.000 10.250 5.000 13.750
                 3.000 13.750 3.000 14.750 5.000 14.750 5.000 18.250 3.000 18.250
                 3.000 19.250 5.000 19.250 5.000 22.750 3.000 22.750 3.000 23.750
                 5.000 23.750 5.000 27.250 3.000 27.250 3.000 28.250 5.000 28.250
                 5.000 31.750 3.000 31.750 3.000 33.080 5.000 33.080 5.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 5.000 1.250 5.000 4.750 3.000 4.750 3.000 5.750 5.000 5.750
                 5.000 9.250 3.000 9.250 3.000 10.250 5.000 10.250 5.000 13.750
                 3.000 13.750 3.000 14.750 5.000 14.750 5.000 18.250 3.000 18.250
                 3.000 19.250 5.000 19.250 5.000 22.750 3.000 22.750 3.000 23.750
                 5.000 23.750 5.000 27.250 3.000 27.250 3.000 28.250 5.000 28.250
                 5.000 31.750 3.000 31.750 3.000 33.080 5.000 33.080 5.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 5.000 1.250 5.000 4.750 3.000 4.750 3.000 5.750 5.000 5.750
                 5.000 9.250 3.000 9.250 3.000 10.250 5.000 10.250 5.000 13.750
                 3.000 13.750 3.000 14.750 5.000 14.750 5.000 18.250 3.000 18.250
                 3.000 19.250 5.000 19.250 5.000 22.750 3.000 22.750 3.000 23.750
                 5.000 23.750 5.000 27.250 3.000 27.250 3.000 28.250 5.000 28.250
                 5.000 31.750 3.000 31.750 3.000 33.080 5.000 33.080 5.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 5.000 1.250 5.000 4.750 3.000 4.750 3.000 5.750 5.000 5.750
                 5.000 9.250 3.000 9.250 3.000 10.250 5.000 10.250 5.000 13.750
                 3.000 13.750 3.000 14.750 5.000 14.750 5.000 18.250 3.000 18.250
                 3.000 19.250 5.000 19.250 5.000 22.750 3.000 22.750 3.000 23.750
                 5.000 23.750 5.000 27.250 3.000 27.250 3.000 28.250 5.000 28.250
                 5.000 31.750 3.000 31.750 3.000 33.080 5.000 33.080 5.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 5.000 1.250 5.000 4.750 3.000 4.750 3.000 5.750 5.000 5.750
                 5.000 9.250 3.000 9.250 3.000 10.250 5.000 10.250 5.000 13.750
                 3.000 13.750 3.000 14.750 5.000 14.750 5.000 18.250 3.000 18.250
                 3.000 19.250 5.000 19.250 5.000 22.750 3.000 22.750 3.000 23.750
                 5.000 23.750 5.000 27.250 3.000 27.250 3.000 28.250 5.000 28.250
                 5.000 31.750 3.000 31.750 3.000 33.080 5.000 33.080 5.000 37.580
                 0.000 37.580 0.000 33.080 2.000 33.080 2.000 31.750 0.000 31.750
                 0.000 28.250 2.000 28.250 2.000 27.250 0.000 27.250 0.000 23.750
                 2.000 23.750 2.000 22.750 0.000 22.750 0.000 19.250 2.000 19.250
                 2.000 18.250 0.000 18.250 0.000 14.750 2.000 14.750 2.000 13.750
                 0.000 13.750 0.000 10.250 2.000 10.250 2.000 9.250 0.000 9.250 0.000 5.750
                 2.000 5.750 2.000 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 5.000 83.670 5.000 87.170 3.000 87.170 3.000 88.020
                 5.000 88.020 5.000 91.520 3.000 91.520 3.000 92.370 5.000 92.370
                 5.000 95.870 3.000 95.870 3.000 96.720 5.000 96.720 5.000 100.220
                 3.000 100.220 3.000 101.070 5.000 101.070 5.000 104.570 3.000 104.570
                 3.000 105.420 5.000 105.420 5.000 108.920 3.000 108.920 3.000 109.770
                 5.000 109.770 5.000 113.270 3.000 113.270 3.000 114.010 5.000 114.010
                 5.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 5.000 83.670 5.000 87.170 3.000 87.170 3.000 88.020
                 5.000 88.020 5.000 91.520 3.000 91.520 3.000 92.370 5.000 92.370
                 5.000 95.870 3.000 95.870 3.000 96.720 5.000 96.720 5.000 100.220
                 3.000 100.220 3.000 101.070 5.000 101.070 5.000 104.570 3.000 104.570
                 3.000 105.420 5.000 105.420 5.000 108.920 3.000 108.920 3.000 109.770
                 5.000 109.770 5.000 113.270 3.000 113.270 3.000 114.010 5.000 114.010
                 5.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 5.000 83.670 5.000 87.170 3.000 87.170 3.000 88.020
                 5.000 88.020 5.000 91.520 3.000 91.520 3.000 92.370 5.000 92.370
                 5.000 95.870 3.000 95.870 3.000 96.720 5.000 96.720 5.000 100.220
                 3.000 100.220 3.000 101.070 5.000 101.070 5.000 104.570 3.000 104.570
                 3.000 105.420 5.000 105.420 5.000 108.920 3.000 108.920 3.000 109.770
                 5.000 109.770 5.000 113.270 3.000 113.270 3.000 114.010 5.000 114.010
                 5.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 5.000 83.670 5.000 87.170 3.000 87.170 3.000 88.020
                 5.000 88.020 5.000 91.520 3.000 91.520 3.000 92.370 5.000 92.370
                 5.000 95.870 3.000 95.870 3.000 96.720 5.000 96.720 5.000 100.220
                 3.000 100.220 3.000 101.070 5.000 101.070 5.000 104.570 3.000 104.570
                 3.000 105.420 5.000 105.420 5.000 108.920 3.000 108.920 3.000 109.770
                 5.000 109.770 5.000 113.270 3.000 113.270 3.000 114.010 5.000 114.010
                 5.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010 2.000 113.270
                 0.000 113.270 0.000 109.770 2.000 109.770 2.000 108.920 0.000 108.920
                 0.000 105.420 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070
                 2.000 101.070 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720
                 2.000 95.870 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520
                 0.000 91.520 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 5.000 83.670 5.000 87.170 3.000 87.170 3.000 88.020
                 5.000 88.020 5.000 91.520 3.000 91.520 3.000 92.370 5.000 92.370
                 5.000 95.870 3.000 95.870 3.000 96.720 5.000 96.720 5.000 100.220
                 3.000 100.220 3.000 101.070 5.000 101.070 5.000 104.570 3.000 104.570
                 3.000 105.420 5.000 105.420 5.000 108.920 0.000 108.920 0.000 105.420
                 2.000 105.420 2.000 104.570 0.000 104.570 0.000 101.070 2.000 101.070
                 2.000 100.220 0.000 100.220 0.000 96.720 2.000 96.720 2.000 95.870
                 0.000 95.870 0.000 92.370 2.000 92.370 2.000 91.520 0.000 91.520
                 0.000 88.020 2.000 88.020 2.000 87.170 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 5.000 82.975 ;
                POLYGON  0.000 40.975 5.000 40.975 5.000 44.475 3.000 44.475 3.000 45.475
                 5.000 45.475 5.000 48.975 3.000 48.975 3.000 49.975 5.000 49.975
                 5.000 53.475 3.000 53.475 3.000 54.475 5.000 54.475 5.000 57.975
                 3.000 57.975 3.000 58.975 5.000 58.975 5.000 62.475 3.000 62.475
                 3.000 63.475 5.000 63.475 5.000 66.975 3.000 66.975 3.000 67.975
                 5.000 67.975 5.000 71.475 3.000 71.475 3.000 72.475 5.000 72.475
                 5.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 5.000 82.975 ;
                POLYGON  0.000 40.975 5.000 40.975 5.000 44.475 3.000 44.475 3.000 45.475
                 5.000 45.475 5.000 48.975 3.000 48.975 3.000 49.975 5.000 49.975
                 5.000 53.475 3.000 53.475 3.000 54.475 5.000 54.475 5.000 57.975
                 3.000 57.975 3.000 58.975 5.000 58.975 5.000 62.475 3.000 62.475
                 3.000 63.475 5.000 63.475 5.000 66.975 3.000 66.975 3.000 67.975
                 5.000 67.975 5.000 71.475 3.000 71.475 3.000 72.475 5.000 72.475
                 5.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 5.000 82.975 ;
                POLYGON  0.000 40.975 5.000 40.975 5.000 44.475 3.000 44.475 3.000 45.475
                 5.000 45.475 5.000 48.975 3.000 48.975 3.000 49.975 5.000 49.975
                 5.000 53.475 3.000 53.475 3.000 54.475 5.000 54.475 5.000 57.975
                 3.000 57.975 3.000 58.975 5.000 58.975 5.000 62.475 3.000 62.475
                 3.000 63.475 5.000 63.475 5.000 66.975 3.000 66.975 3.000 67.975
                 5.000 67.975 5.000 71.475 3.000 71.475 3.000 72.475 5.000 72.475
                 5.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 5.000 82.975 ;
                POLYGON  0.000 40.975 5.000 40.975 5.000 44.475 3.000 44.475 3.000 45.475
                 5.000 45.475 5.000 48.975 3.000 48.975 3.000 49.975 5.000 49.975
                 5.000 53.475 3.000 53.475 3.000 54.475 5.000 54.475 5.000 57.975
                 3.000 57.975 3.000 58.975 5.000 58.975 5.000 62.475 3.000 62.475
                 3.000 63.475 5.000 63.475 5.000 66.975 3.000 66.975 3.000 67.975
                 5.000 67.975 5.000 71.475 3.000 71.475 3.000 72.475 5.000 72.475
                 5.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 5.000 82.975 ;
                POLYGON  0.000 40.975 5.000 40.975 5.000 44.475 3.000 44.475 3.000 45.475
                 5.000 45.475 5.000 48.975 3.000 48.975 3.000 49.975 5.000 49.975
                 5.000 53.475 3.000 53.475 3.000 54.475 5.000 54.475 5.000 57.975
                 3.000 57.975 3.000 58.975 5.000 58.975 5.000 62.475 3.000 62.475
                 3.000 63.475 5.000 63.475 5.000 66.975 3.000 66.975 3.000 67.975
                 5.000 67.975 5.000 71.475 3.000 71.475 3.000 72.475 5.000 72.475
                 5.000 75.975 0.000 75.975 0.000 72.475 2.000 72.475 2.000 71.475
                 0.000 71.475 0.000 67.975 2.000 67.975 2.000 66.975 0.000 66.975
                 0.000 63.475 2.000 63.475 2.000 62.475 0.000 62.475 0.000 58.975
                 2.000 58.975 2.000 57.975 0.000 57.975 0.000 54.475 2.000 54.475
                 2.000 53.475 0.000 53.475 0.000 49.975 2.000 49.975 2.000 48.975
                 0.000 48.975 0.000 45.475 2.000 45.475 2.000 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 5.000 109.770 5.000 113.270 3.000 113.270 3.000 114.010
                 5.000 114.010 5.000 117.510 0.000 117.510 0.000 114.010 2.000 114.010
                 2.000 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 5.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA2 ;
        RECT  3.000 1.250 5.000 4.750 ;
        RECT  3.000 5.750 5.000 9.250 ;
        RECT  3.000 10.250 5.000 13.750 ;
        RECT  3.000 14.750 5.000 18.250 ;
        RECT  3.000 19.250 5.000 22.750 ;
        RECT  3.000 23.750 5.000 27.250 ;
        RECT  3.000 28.250 5.000 31.750 ;
        RECT  3.000 33.080 5.000 37.580 ;
        RECT  3.000 40.975 5.000 44.475 ;
        RECT  3.000 45.475 5.000 48.975 ;
        RECT  3.000 49.975 5.000 53.475 ;
        RECT  3.000 54.475 5.000 57.975 ;
        RECT  3.000 58.975 5.000 62.475 ;
        RECT  3.000 63.475 5.000 66.975 ;
        RECT  3.000 67.975 5.000 71.475 ;
        RECT  3.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  3.000 83.670 5.000 87.170 ;
        RECT  3.000 88.020 5.000 91.520 ;
        RECT  3.000 92.370 5.000 95.870 ;
        RECT  3.000 96.720 5.000 100.220 ;
        RECT  3.000 101.070 5.000 104.570 ;
        RECT  3.000 105.420 5.000 108.920 ;
        RECT  3.000 109.770 5.000 113.270 ;
        RECT  3.000 114.010 5.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 108.920 ;
        RECT  2.000 109.770 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA3 ;
        RECT  3.000 1.250 5.000 4.750 ;
        RECT  3.000 5.750 5.000 9.250 ;
        RECT  3.000 10.250 5.000 13.750 ;
        RECT  3.000 14.750 5.000 18.250 ;
        RECT  3.000 19.250 5.000 22.750 ;
        RECT  3.000 23.750 5.000 27.250 ;
        RECT  3.000 28.250 5.000 31.750 ;
        RECT  3.000 33.080 5.000 37.580 ;
        RECT  3.000 40.975 5.000 44.475 ;
        RECT  3.000 45.475 5.000 48.975 ;
        RECT  3.000 49.975 5.000 53.475 ;
        RECT  3.000 54.475 5.000 57.975 ;
        RECT  3.000 58.975 5.000 62.475 ;
        RECT  3.000 63.475 5.000 66.975 ;
        RECT  3.000 67.975 5.000 71.475 ;
        RECT  3.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  3.000 83.670 5.000 87.170 ;
        RECT  3.000 88.020 5.000 91.520 ;
        RECT  3.000 92.370 5.000 95.870 ;
        RECT  3.000 96.720 5.000 100.220 ;
        RECT  3.000 101.070 5.000 104.570 ;
        RECT  3.000 105.420 5.000 108.920 ;
        RECT  3.000 109.770 5.000 113.270 ;
        RECT  3.000 114.010 5.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA4 ;
        RECT  3.000 1.250 5.000 4.750 ;
        RECT  3.000 5.750 5.000 9.250 ;
        RECT  3.000 10.250 5.000 13.750 ;
        RECT  3.000 14.750 5.000 18.250 ;
        RECT  3.000 19.250 5.000 22.750 ;
        RECT  3.000 23.750 5.000 27.250 ;
        RECT  3.000 28.250 5.000 31.750 ;
        RECT  3.000 33.080 5.000 37.580 ;
        RECT  3.000 40.975 5.000 44.475 ;
        RECT  3.000 45.475 5.000 48.975 ;
        RECT  3.000 49.975 5.000 53.475 ;
        RECT  3.000 54.475 5.000 57.975 ;
        RECT  3.000 58.975 5.000 62.475 ;
        RECT  3.000 63.475 5.000 66.975 ;
        RECT  3.000 67.975 5.000 71.475 ;
        RECT  3.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  3.000 83.670 5.000 87.170 ;
        RECT  3.000 88.020 5.000 91.520 ;
        RECT  3.000 92.370 5.000 95.870 ;
        RECT  3.000 96.720 5.000 100.220 ;
        RECT  3.000 101.070 5.000 104.570 ;
        RECT  3.000 105.420 5.000 108.920 ;
        RECT  3.000 109.770 5.000 113.270 ;
        RECT  3.000 114.010 5.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA5 ;
        RECT  3.000 1.250 5.000 4.750 ;
        RECT  3.000 5.750 5.000 9.250 ;
        RECT  3.000 10.250 5.000 13.750 ;
        RECT  3.000 14.750 5.000 18.250 ;
        RECT  3.000 19.250 5.000 22.750 ;
        RECT  3.000 23.750 5.000 27.250 ;
        RECT  3.000 28.250 5.000 31.750 ;
        RECT  3.000 33.080 5.000 37.580 ;
        RECT  3.000 40.975 5.000 44.475 ;
        RECT  3.000 45.475 5.000 48.975 ;
        RECT  3.000 49.975 5.000 53.475 ;
        RECT  3.000 54.475 5.000 57.975 ;
        RECT  3.000 58.975 5.000 62.475 ;
        RECT  3.000 63.475 5.000 66.975 ;
        RECT  3.000 67.975 5.000 71.475 ;
        RECT  3.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  3.000 83.670 5.000 87.170 ;
        RECT  3.000 88.020 5.000 91.520 ;
        RECT  3.000 92.370 5.000 95.870 ;
        RECT  3.000 96.720 5.000 100.220 ;
        RECT  3.000 101.070 5.000 104.570 ;
        RECT  3.000 105.420 5.000 108.920 ;
        RECT  3.000 109.770 5.000 113.270 ;
        RECT  3.000 114.010 5.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 5.000 120.000 ;
        LAYER VIA6 ;
        RECT  3.000 1.250 5.000 4.750 ;
        RECT  3.000 5.750 5.000 9.250 ;
        RECT  3.000 10.250 5.000 13.750 ;
        RECT  3.000 14.750 5.000 18.250 ;
        RECT  3.000 19.250 5.000 22.750 ;
        RECT  3.000 23.750 5.000 27.250 ;
        RECT  3.000 28.250 5.000 31.750 ;
        RECT  3.000 33.080 5.000 37.580 ;
        RECT  3.000 40.975 5.000 44.475 ;
        RECT  3.000 45.475 5.000 48.975 ;
        RECT  3.000 49.975 5.000 53.475 ;
        RECT  3.000 54.475 5.000 57.975 ;
        RECT  3.000 58.975 5.000 62.475 ;
        RECT  3.000 63.475 5.000 66.975 ;
        RECT  3.000 67.975 5.000 71.475 ;
        RECT  3.000 72.475 5.000 75.975 ;
        RECT  0.000 79.975 5.000 82.975 ;
        RECT  3.000 83.670 5.000 87.170 ;
        RECT  3.000 88.020 5.000 91.520 ;
        RECT  3.000 92.370 5.000 95.870 ;
        RECT  3.000 96.720 5.000 100.220 ;
        RECT  3.000 101.070 5.000 104.570 ;
        RECT  3.000 105.420 5.000 108.920 ;
        RECT  3.000 109.770 5.000 113.270 ;
        RECT  3.000 114.010 5.000 117.510 ;
        RECT  2.000 1.250 3.000 37.580 ;
        RECT  2.000 40.975 3.000 75.975 ;
        RECT  2.000 83.670 3.000 117.510 ;
        RECT  0.000 1.250 2.000 4.750 ;
        RECT  0.000 5.750 2.000 9.250 ;
        RECT  0.000 10.250 2.000 13.750 ;
        RECT  0.000 14.750 2.000 18.250 ;
        RECT  0.000 19.250 2.000 22.750 ;
        RECT  0.000 23.750 2.000 27.250 ;
        RECT  0.000 28.250 2.000 31.750 ;
        RECT  0.000 33.080 2.000 37.580 ;
        RECT  0.000 40.975 2.000 44.475 ;
        RECT  0.000 45.475 2.000 48.975 ;
        RECT  0.000 49.975 2.000 53.475 ;
        RECT  0.000 54.475 2.000 57.975 ;
        RECT  0.000 58.975 2.000 62.475 ;
        RECT  0.000 63.475 2.000 66.975 ;
        RECT  0.000 67.975 2.000 71.475 ;
        RECT  0.000 72.475 2.000 75.975 ;
        RECT  0.000 83.670 2.000 87.170 ;
        RECT  0.000 88.020 2.000 91.520 ;
        RECT  0.000 92.370 2.000 95.870 ;
        RECT  0.000 96.720 2.000 100.220 ;
        RECT  0.000 101.070 2.000 104.570 ;
        RECT  0.000 105.420 2.000 108.920 ;
        RECT  0.000 109.770 2.000 113.270 ;
        RECT  0.000 114.010 2.000 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 5.000 120.000 ;
    END
END PFILLER5_G

MACRO PRCUTA_G
    CLASS PAD ;
    FOREIGN PRCUTA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRCUTA_G

MACRO PRCUT_G
    CLASS PAD ;
    FOREIGN PRCUT_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRCUT_G

MACRO PRDW08DGZ_G
    CLASS PAD ;
    FOREIGN PRDW08DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW08DGZ_G

MACRO PRDW08SDGZ_G
    CLASS PAD ;
    FOREIGN PRDW08SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW08SDGZ_G

MACRO PRDW12DGZ_G
    CLASS PAD ;
    FOREIGN PRDW12DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW12DGZ_G

MACRO PRDW12SDGZ_G
    CLASS PAD ;
    FOREIGN PRDW12SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW12SDGZ_G

MACRO PRDW16DGZ_G
    CLASS PAD ;
    FOREIGN PRDW16DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW16DGZ_G

MACRO PRDW16SDGZ_G
    CLASS PAD ;
    FOREIGN PRDW16SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRDW16SDGZ_G

MACRO PRUW08DGZ_G
    CLASS PAD ;
    FOREIGN PRUW08DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW08DGZ_G

MACRO PRUW08SDGZ_G
    CLASS PAD ;
    FOREIGN PRUW08SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW08SDGZ_G

MACRO PRUW12DGZ_G
    CLASS PAD ;
    FOREIGN PRUW12DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW12DGZ_G

MACRO PRUW12SDGZ_G
    CLASS PAD ;
    FOREIGN PRUW12SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW12SDGZ_G

MACRO PRUW16DGZ_G
    CLASS PAD ;
    FOREIGN PRUW16DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW16DGZ_G

MACRO PRUW16SDGZ_G
    CLASS PAD ;
    FOREIGN PRUW16SDGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN REN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M6 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M5 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M4 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M3 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M2 ;
        RECT  15.550 119.000 18.440 120.000 ;
        LAYER M1 ;
        RECT  15.550 119.000 18.440 120.000 ;
        END
        ANTENNAGATEAREA 8.1200 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.3072 LAYER M1 ;
        ANTENNAMAXAREACAR 11.9554 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5586 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 8.1200 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 3.3258 LAYER M2 ;
        ANTENNAMAXAREACAR 12.3649 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3485 LAYER VIA2 ;
        ANTENNAGATEAREA 8.1200 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.7208 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4137 LAYER VIA3 ;
        ANTENNAGATEAREA 8.1200 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 13.0768 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.4789 LAYER VIA4 ;
        ANTENNAGATEAREA 8.1200 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4327 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.5440 LAYER VIA5 ;
        ANTENNAGATEAREA 8.1200 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.7886 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.6092 LAYER VIA6 ;
        ANTENNAGATEAREA 8.1200 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.1445 LAYER M7 ;
    END REN
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        END
        ANTENNADIFFAREA 928.8100 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA3 ;
        ANTENNADIFFAREA 928.8100 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA4 ;
        ANTENNADIFFAREA 928.8100 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA5 ;
        ANTENNADIFFAREA 928.8100 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 11.1132 LAYER VIA6 ;
        ANTENNADIFFAREA 928.8100 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 60.6900 LAYER M7 ;
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M6 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M5 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M4 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M3 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M2 ;
        RECT  11.590 119.000 14.480 120.000 ;
        LAYER M1 ;
        RECT  11.590 119.000 14.480 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 7.4753 LAYER M1 ;
        ANTENNAMAXAREACAR 17.1963 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.6174 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.7967 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 5.2982 LAYER M2 ;
        ANTENNAMAXAREACAR 18.0677 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.8837 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 18.5431 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.9707 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 19.0184 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 2.0578 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 19.4937 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 2.1448 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 19.9691 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 2.2319 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 20.4444 LAYER M7 ;
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M4 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M3 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M1 ;
        RECT  0.995 119.000 3.885 120.000 ;
        END
        ANTENNAGATEAREA 6.0800 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 6.9162 LAYER M1 ;
        ANTENNAMAXAREACAR 11.1877 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5978 LAYER VIA1 ;
        ANTENNAMAXAREACAR 1.2833 LAYER VIA1 ;
        ANTENNAGATEAREA 6.0800 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 4.8677 LAYER M2 ;
        ANTENNAMAXAREACAR 11.9883 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNAMAXAREACAR 1.3704 LAYER VIA2 ;
        ANTENNAGATEAREA 6.0800 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAMAXAREACAR 12.4637 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNAMAXAREACAR 1.4574 LAYER VIA3 ;
        ANTENNAGATEAREA 6.0800 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAMAXAREACAR 12.9390 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNAMAXAREACAR 1.5445 LAYER VIA4 ;
        ANTENNAGATEAREA 6.0800 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAMAXAREACAR 13.4143 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNAMAXAREACAR 1.6315 LAYER VIA5 ;
        ANTENNAGATEAREA 6.0800 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAMAXAREACAR 13.8897 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNAMAXAREACAR 1.7185 LAYER VIA6 ;
        ANTENNAGATEAREA 6.0800 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
        ANTENNAMAXAREACAR 14.3650 LAYER M7 ;
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M6 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M5 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M4 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M3 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M2 ;
        RECT  21.230 119.000 24.120 120.000 ;
        LAYER M1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        END
        ANTENNADIFFAREA 1.0700 LAYER M1 ;
        ANTENNAPARTIALMETALAREA 5.2015 LAYER M1 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA1 ;
        ANTENNADIFFAREA 1.0700 LAYER M2 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M2 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA2 ;
        ANTENNADIFFAREA 1.0700 LAYER M3 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M3 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA3 ;
        ANTENNADIFFAREA 1.0700 LAYER M4 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M4 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA4 ;
        ANTENNADIFFAREA 1.0700 LAYER M5 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M5 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA5 ;
        ANTENNADIFFAREA 1.0700 LAYER M6 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M6 ;
        ANTENNAPARTIALCUTAREA 0.5292 LAYER VIA6 ;
        ANTENNADIFFAREA 1.0700 LAYER M7 ;
        ANTENNAPARTIALMETALAREA 2.8900 LAYER M7 ;
    END C
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 24.085 37.580 24.085 40.710 23.755 40.710 23.755 37.580
                 20.445 37.580 20.445 40.230 19.955 40.230 19.955 37.580 14.285 37.580
                 14.285 40.230 13.795 40.230 13.795 37.580 8.125 37.580 8.125 40.230
                 7.635 40.230 7.635 37.580 1.435 37.580 1.435 40.710 0.945 40.710
                 0.945 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.585 40.975 1.585 39.450 1.915 39.450 1.915 40.975
                 4.555 40.975 4.555 39.450 5.045 39.450 5.045 40.975 10.715 40.975
                 10.715 39.450 11.205 39.450 11.205 40.975 16.875 40.975 16.875 39.450
                 17.365 39.450 17.365 40.975 23.115 40.975 23.115 39.450 23.605 39.450
                 23.605 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  24.085 33.080 25.000 37.580 ;
        RECT  23.605 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  23.755 33.080 24.085 40.710 ;
        RECT  20.445 33.080 23.755 37.580 ;
        RECT  23.115 39.450 23.605 44.475 ;
        RECT  17.365 40.975 23.115 44.475 ;
        RECT  19.955 33.080 20.445 40.230 ;
        RECT  14.285 33.080 19.955 37.580 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  16.875 39.450 17.365 44.475 ;
        RECT  13.880 40.975 16.875 44.475 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  13.880 33.080 14.285 40.230 ;
        RECT  13.795 1.250 13.880 40.230 ;
        RECT  11.205 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.120 1.250 13.795 37.580 ;
        RECT  11.120 39.450 11.205 75.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  8.125 33.080 11.120 37.580 ;
        RECT  10.715 39.450 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  5.045 40.975 10.715 44.475 ;
        RECT  7.635 33.080 8.125 40.230 ;
        RECT  1.435 33.080 7.635 37.580 ;
        RECT  4.555 39.450 5.045 44.475 ;
        RECT  1.915 40.975 4.555 44.475 ;
        RECT  0.995 119.000 3.885 120.000 ;
        RECT  1.585 39.450 1.915 44.475 ;
        RECT  0.000 40.975 1.585 44.475 ;
        RECT  0.945 33.080 1.435 40.710 ;
        RECT  0.000 33.080 0.945 37.580 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  21.230 119.000 24.120 120.000 ;
        RECT  15.550 119.000 18.440 120.000 ;
        RECT  11.590 119.000 14.480 120.000 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  0.995 119.000 3.885 120.000 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PRUW16SDGZ_G

MACRO PVBUS_G
    CLASS PAD ;
    FOREIGN PVBUS_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VBUS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  2.38 118.2 4.14 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  7 118.2 8.76 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.62 118.2 13.38 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  16.24 118.2 18 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  20.86 118.2 22.62 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  2.285 118.2 4.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.905 118.2 8.855 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.525 118.2 13.475 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  16.145 118.2 18.095 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  20.765 118.2 22.715 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.285 76.475 22.715 79.475 ;
        LAYER M2 ;
        RECT  20.765 118.200 22.715 120.000 ;
        RECT  16.145 118.200 18.095 120.000 ;
        RECT  11.525 118.200 13.475 120.000 ;
        RECT  6.905 118.200 8.855 120.000 ;
        RECT  2.285 118.200 4.235 120.000 ;
        LAYER M1 ;
        RECT  20.860 118.200 22.620 120.000 ;
        RECT  16.240 118.200 18.000 120.000 ;
        RECT  11.620 118.200 13.380 120.000 ;
        RECT  7.000 118.200 8.760 120.000 ;
        RECT  2.380 118.200 4.140 120.000 ;
        END
    END VBUS
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  20.765 118.200 22.715 120.000 ;
        RECT  16.145 118.200 18.095 120.000 ;
        RECT  11.525 118.200 13.475 120.000 ;
        RECT  6.905 118.200 8.855 120.000 ;
        RECT  2.285 118.200 4.235 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVBUS_G

MACRO PVDD1ANA_G
    CLASS PAD ;
    FOREIGN PVDD1ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    PIN AVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  2.525 118.5 3.095 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  3.545 118.5 4.115 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  4.565 118.5 5.135 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.585 118.5 6.155 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  6.605 118.5 7.175 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  7.625 118.5 8.195 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.645 118.5 9.215 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  9.665 118.5 10.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  10.685 118.5 11.255 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.705 118.5 12.275 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  12.725 118.5 13.295 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  13.745 118.5 14.315 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.765 118.5 15.335 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.785 118.5 16.355 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  16.805 118.5 17.375 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  17.825 118.5 18.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  18.845 118.5 19.415 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  19.865 118.5 20.435 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  20.885 118.5 21.455 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.905 118.5 22.475 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  2.525 118.5 3.095 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  3.545 118.5 4.115 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  4.565 118.5 5.135 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.585 118.5 6.155 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.605 118.5 7.175 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  7.625 118.5 8.195 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.645 118.5 9.215 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  9.665 118.5 10.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  10.685 118.5 11.255 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.705 118.5 12.275 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  12.725 118.5 13.295 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  13.745 118.5 14.315 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.765 118.5 15.335 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  15.785 118.5 16.355 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  16.805 118.5 17.375 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  17.825 118.5 18.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  18.845 118.5 19.415 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  19.865 118.5 20.435 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  20.885 118.5 21.455 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.905 118.5 22.475 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M2 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        LAYER M1 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD1ANA_G

MACRO PVDD1DGZ_G
    CLASS PAD ;
    FOREIGN PVDD1DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  2.525 118.5 3.095 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  3.545 118.5 4.115 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  4.565 118.5 5.135 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.585 118.5 6.155 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  6.605 118.5 7.175 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  7.625 118.5 8.195 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.645 118.5 9.215 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  9.665 118.5 10.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  10.685 118.5 11.255 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.705 118.5 12.275 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  12.725 118.5 13.295 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  13.745 118.5 14.315 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.765 118.5 15.335 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.785 118.5 16.355 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  16.805 118.5 17.375 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  17.825 118.5 18.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  18.845 118.5 19.415 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  19.865 118.5 20.435 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  20.885 118.5 21.455 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.905 118.5 22.475 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  2.525 118.5 3.095 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  3.545 118.5 4.115 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  4.565 118.5 5.135 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.585 118.5 6.155 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.605 118.5 7.175 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  7.625 118.5 8.195 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.645 118.5 9.215 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  9.665 118.5 10.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  10.685 118.5 11.255 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.705 118.5 12.275 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  12.725 118.5 13.295 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  13.745 118.5 14.315 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.765 118.5 15.335 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  15.785 118.5 16.355 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  16.805 118.5 17.375 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  17.825 118.5 18.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  18.845 118.5 19.415 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  19.865 118.5 20.435 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  20.885 118.5 21.455 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.905 118.5 22.475 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        LAYER M2 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        LAYER M1 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.905 118.500 22.475 120.000 ;
        RECT  20.885 118.500 21.455 120.000 ;
        RECT  19.865 118.500 20.435 120.000 ;
        RECT  18.845 118.500 19.415 120.000 ;
        RECT  17.825 118.500 18.395 120.000 ;
        RECT  16.805 118.500 17.375 120.000 ;
        RECT  15.785 118.500 16.355 120.000 ;
        RECT  14.765 118.500 15.335 120.000 ;
        RECT  13.745 118.500 14.315 120.000 ;
        RECT  12.725 118.500 13.295 120.000 ;
        RECT  11.705 118.500 12.275 120.000 ;
        RECT  10.685 118.500 11.255 120.000 ;
        RECT  9.665 118.500 10.235 120.000 ;
        RECT  8.645 118.500 9.215 120.000 ;
        RECT  7.625 118.500 8.195 120.000 ;
        RECT  6.605 118.500 7.175 120.000 ;
        RECT  5.585 118.500 6.155 120.000 ;
        RECT  4.565 118.500 5.135 120.000 ;
        RECT  3.545 118.500 4.115 120.000 ;
        RECT  2.525 118.500 3.095 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD1DGZ_G

MACRO PVDD2ANA_G
    CLASS PAD ;
    FOREIGN PVDD2ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 1.120 40.975 1.120 39.450 1.450 39.450 1.450 40.975
                 23.550 40.975 23.550 39.450 23.880 39.450 23.880 40.975 25.000 40.975
                 25.000 44.475 13.880 44.475 13.880 45.475 25.000 45.475 25.000 48.975
                 13.880 48.975 13.880 49.975 25.000 49.975 25.000 53.475 13.880 53.475
                 13.880 54.475 25.000 54.475 25.000 57.975 13.880 57.975 13.880 58.975
                 25.000 58.975 25.000 62.475 13.880 62.475 13.880 63.475 25.000 63.475
                 25.000 66.975 13.880 66.975 13.880 67.975 25.000 67.975 25.000 71.475
                 13.880 71.475 13.880 72.475 25.000 72.475 25.000 75.975 0.000 75.975
                 0.000 72.475 11.120 72.475 11.120 71.475 0.000 71.475 0.000 67.975
                 11.120 67.975 11.120 66.975 0.000 66.975 0.000 63.475 11.120 63.475
                 11.120 62.475 0.000 62.475 0.000 58.975 11.120 58.975 11.120 57.975
                 0.000 57.975 0.000 54.475 11.120 54.475 11.120 53.475 0.000 53.475
                 0.000 49.975 11.120 49.975 11.120 48.975 0.000 48.975 0.000 45.475
                 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    PIN AVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  3.15 118.5 5.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  7.15 118.5 9.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.15 118.5 13.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.15 118.5 17.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  19.15 118.5 21.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  3.15 118.5 5.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  7.15 118.5 9.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.15 118.5 13.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  15.15 118.5 17.85 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  19.15 118.5 21.85 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  2.310 76.475 22.690 79.475 ;
        LAYER M2 ;
        RECT  19.150 118.500 21.850 120.000 ;
        RECT  15.150 118.500 17.850 120.000 ;
        RECT  11.150 118.500 13.850 120.000 ;
        RECT  7.150 118.500 9.850 120.000 ;
        RECT  3.150 118.500 5.850 120.000 ;
        LAYER M1 ;
        RECT  19.150 118.500 21.850 120.000 ;
        RECT  15.150 118.500 17.850 120.000 ;
        RECT  11.150 118.500 13.850 120.000 ;
        RECT  7.150 118.500 9.850 120.000 ;
        RECT  3.150 118.500 5.850 120.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  19.150 118.500 21.850 120.000 ;
        RECT  15.150 118.500 17.850 120.000 ;
        RECT  11.150 118.500 13.850 120.000 ;
        RECT  7.150 118.500 9.850 120.000 ;
        RECT  3.150 118.500 5.850 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  23.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  23.550 39.450 23.880 44.475 ;
        RECT  13.880 40.975 23.550 44.475 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.450 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  1.120 39.450 1.450 44.475 ;
        RECT  0.000 40.975 1.120 44.475 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  23.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  23.550 39.450 23.880 44.475 ;
        RECT  13.880 40.975 23.550 44.475 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.450 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  1.120 39.450 1.450 44.475 ;
        RECT  0.000 40.975 1.120 44.475 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD2ANA_G

MACRO PVDD2DGZ_G
    CLASS PAD ;
    FOREIGN PVDD2DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
                POLYGON  0.000 40.975 0.915 40.975 0.915 39.450 1.245 39.450 1.245 40.975
                 23.755 40.975 23.755 39.450 24.085 39.450 24.085 40.975 25.000 40.975
                 25.000 44.475 13.880 44.475 13.880 45.475 25.000 45.475 25.000 48.975
                 13.880 48.975 13.880 49.975 25.000 49.975 25.000 53.475 13.880 53.475
                 13.880 54.475 25.000 54.475 25.000 57.975 13.880 57.975 13.880 58.975
                 25.000 58.975 25.000 62.475 13.880 62.475 13.880 63.475 25.000 63.475
                 25.000 66.975 13.880 66.975 13.880 67.975 25.000 67.975 25.000 71.475
                 13.880 71.475 13.880 72.475 25.000 72.475 25.000 75.975 23.135 75.975
                 23.135 79.975 25.000 79.975 25.000 82.975 21.885 82.975 21.885 75.975
                 21.315 75.975 21.315 76.475 21.885 76.475 21.885 79.475 21.315 79.475
                 21.315 79.975 21.885 79.975 21.885 82.975 20.065 82.975 20.065 75.975
                 19.495 75.975 19.495 76.475 20.065 76.475 20.065 79.475 19.495 79.475
                 19.495 79.975 20.065 79.975 20.065 82.975 18.245 82.975 18.245 75.975
                 17.675 75.975 17.675 76.475 18.245 76.475 18.245 79.475 17.675 79.475
                 17.675 79.975 18.245 79.975 18.245 82.975 16.425 82.975 16.425 75.975
                 15.855 75.975 15.855 76.475 16.425 76.475 16.425 79.475 15.855 79.475
                 15.855 79.975 16.425 79.975 16.425 82.975 14.605 82.975 14.605 75.975
                 14.035 75.975 14.035 76.475 14.605 76.475 14.605 79.475 14.035 79.475
                 14.035 79.975 14.605 79.975 14.605 82.975 12.785 82.975 12.785 75.975
                 12.215 75.975 12.215 76.475 12.785 76.475 12.785 79.475 12.215 79.475
                 12.215 79.975 12.785 79.975 12.785 82.975 10.965 82.975 10.965 75.975
                 10.395 75.975 10.395 76.475 10.965 76.475 10.965 79.475 10.395 79.475
                 10.395 79.975 10.965 79.975 10.965 82.975 9.145 82.975 9.145 75.975
                 8.575 75.975 8.575 76.475 9.145 76.475 9.145 79.475 8.575 79.475
                 8.575 79.975 9.145 79.975 9.145 82.975 7.325 82.975 7.325 75.975
                 6.755 75.975 6.755 76.475 7.325 76.475 7.325 79.475 6.755 79.475
                 6.755 79.975 7.325 79.975 7.325 82.975 5.505 82.975 5.505 75.975
                 4.935 75.975 4.935 76.475 5.505 76.475 5.505 79.475 4.935 79.475
                 4.935 79.975 5.505 79.975 5.505 82.975 3.685 82.975 3.685 75.975
                 3.115 75.975 3.115 76.475 3.685 76.475 3.685 79.475 3.115 79.475
                 3.115 79.975 3.685 79.975 3.685 82.975 0.000 82.975 0.000 79.975
                 1.865 79.975 1.865 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  24.085 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.135 72.475 25.000 75.975 ;
        RECT  23.135 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  23.755 39.450 24.085 44.475 ;
        RECT  13.880 40.975 23.755 44.475 ;
        RECT  21.885 72.475 23.135 82.975 ;
        RECT  21.315 72.475 21.885 75.975 ;
        RECT  21.315 76.475 21.885 79.475 ;
        RECT  21.315 79.975 21.885 82.975 ;
        RECT  20.065 72.475 21.315 82.975 ;
        RECT  19.495 72.475 20.065 75.975 ;
        RECT  19.495 76.475 20.065 79.475 ;
        RECT  19.495 79.975 20.065 82.975 ;
        RECT  18.245 72.475 19.495 82.975 ;
        RECT  17.675 72.475 18.245 75.975 ;
        RECT  17.675 76.475 18.245 79.475 ;
        RECT  17.675 79.975 18.245 82.975 ;
        RECT  16.425 72.475 17.675 82.975 ;
        RECT  15.855 72.475 16.425 75.975 ;
        RECT  15.855 76.475 16.425 79.475 ;
        RECT  15.855 79.975 16.425 82.975 ;
        RECT  14.605 72.475 15.855 82.975 ;
        RECT  14.035 72.475 14.605 75.975 ;
        RECT  14.035 76.475 14.605 79.475 ;
        RECT  14.035 79.975 14.605 82.975 ;
        RECT  13.880 72.475 14.035 82.975 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  12.785 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  12.215 40.975 12.785 75.975 ;
        RECT  12.215 76.475 12.785 79.475 ;
        RECT  12.215 79.975 12.785 82.975 ;
        RECT  11.120 40.975 12.215 82.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.245 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.965 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.395 72.475 10.965 75.975 ;
        RECT  10.395 76.475 10.965 79.475 ;
        RECT  10.395 79.975 10.965 82.975 ;
        RECT  9.145 72.475 10.395 82.975 ;
        RECT  8.575 72.475 9.145 75.975 ;
        RECT  8.575 76.475 9.145 79.475 ;
        RECT  8.575 79.975 9.145 82.975 ;
        RECT  7.325 72.475 8.575 82.975 ;
        RECT  6.755 72.475 7.325 75.975 ;
        RECT  6.755 76.475 7.325 79.475 ;
        RECT  6.755 79.975 7.325 82.975 ;
        RECT  5.505 72.475 6.755 82.975 ;
        RECT  4.935 72.475 5.505 75.975 ;
        RECT  4.935 76.475 5.505 79.475 ;
        RECT  4.935 79.975 5.505 82.975 ;
        RECT  3.685 72.475 4.935 82.975 ;
        RECT  3.115 72.475 3.685 75.975 ;
        RECT  3.115 76.475 3.685 79.475 ;
        RECT  3.115 79.975 3.685 82.975 ;
        RECT  1.865 72.475 3.115 82.975 ;
        RECT  0.000 72.475 1.865 75.975 ;
        RECT  0.000 79.975 1.865 82.975 ;
        RECT  0.915 39.450 1.245 44.475 ;
        RECT  0.000 40.975 0.915 44.475 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  24.085 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.135 72.475 25.000 75.975 ;
        RECT  23.135 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  23.755 39.450 24.085 44.475 ;
        RECT  13.880 40.975 23.755 44.475 ;
        RECT  21.885 72.475 23.135 82.975 ;
        RECT  21.315 72.475 21.885 75.975 ;
        RECT  21.315 76.475 21.885 79.475 ;
        RECT  21.315 79.975 21.885 82.975 ;
        RECT  20.065 72.475 21.315 82.975 ;
        RECT  19.495 72.475 20.065 75.975 ;
        RECT  19.495 76.475 20.065 79.475 ;
        RECT  19.495 79.975 20.065 82.975 ;
        RECT  18.245 72.475 19.495 82.975 ;
        RECT  17.675 72.475 18.245 75.975 ;
        RECT  17.675 76.475 18.245 79.475 ;
        RECT  17.675 79.975 18.245 82.975 ;
        RECT  16.425 72.475 17.675 82.975 ;
        RECT  15.855 72.475 16.425 75.975 ;
        RECT  15.855 76.475 16.425 79.475 ;
        RECT  15.855 79.975 16.425 82.975 ;
        RECT  14.605 72.475 15.855 82.975 ;
        RECT  14.035 72.475 14.605 75.975 ;
        RECT  14.035 76.475 14.605 79.475 ;
        RECT  14.035 79.975 14.605 82.975 ;
        RECT  13.880 72.475 14.035 82.975 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  12.785 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  12.215 40.975 12.785 75.975 ;
        RECT  12.215 76.475 12.785 79.475 ;
        RECT  12.215 79.975 12.785 82.975 ;
        RECT  11.120 40.975 12.215 82.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.245 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.965 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.395 72.475 10.965 75.975 ;
        RECT  10.395 76.475 10.965 79.475 ;
        RECT  10.395 79.975 10.965 82.975 ;
        RECT  9.145 72.475 10.395 82.975 ;
        RECT  8.575 72.475 9.145 75.975 ;
        RECT  8.575 76.475 9.145 79.475 ;
        RECT  8.575 79.975 9.145 82.975 ;
        RECT  7.325 72.475 8.575 82.975 ;
        RECT  6.755 72.475 7.325 75.975 ;
        RECT  6.755 76.475 7.325 79.475 ;
        RECT  6.755 79.975 7.325 82.975 ;
        RECT  5.505 72.475 6.755 82.975 ;
        RECT  4.935 72.475 5.505 75.975 ;
        RECT  4.935 76.475 5.505 79.475 ;
        RECT  4.935 79.975 5.505 82.975 ;
        RECT  3.685 72.475 4.935 82.975 ;
        RECT  3.115 72.475 3.685 75.975 ;
        RECT  3.115 76.475 3.685 79.475 ;
        RECT  3.115 79.975 3.685 82.975 ;
        RECT  1.865 72.475 3.115 82.975 ;
        RECT  0.000 72.475 1.865 75.975 ;
        RECT  0.000 79.975 1.865 82.975 ;
        RECT  0.915 39.450 1.245 44.475 ;
        RECT  0.000 40.975 0.915 44.475 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD2DGZ_G

MACRO PVDD2POC_G
    CLASS PAD ;
    FOREIGN PVDD2POC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
                POLYGON  0.000 40.975 0.915 40.975 0.915 39.450 1.245 39.450 1.245 40.975
                 23.755 40.975 23.755 39.450 24.085 39.450 24.085 40.975 25.000 40.975
                 25.000 44.475 13.880 44.475 13.880 45.475 25.000 45.475 25.000 48.975
                 13.880 48.975 13.880 49.975 25.000 49.975 25.000 53.475 13.880 53.475
                 13.880 54.475 25.000 54.475 25.000 57.975 13.880 57.975 13.880 58.975
                 25.000 58.975 25.000 62.475 13.880 62.475 13.880 63.475 25.000 63.475
                 25.000 66.975 13.880 66.975 13.880 67.975 25.000 67.975 25.000 71.475
                 13.880 71.475 13.880 72.475 25.000 72.475 25.000 75.975 23.135 75.975
                 23.135 79.975 25.000 79.975 25.000 82.975 21.885 82.975 21.885 75.975
                 21.315 75.975 21.315 76.475 21.885 76.475 21.885 79.475 21.315 79.475
                 21.315 79.975 21.885 79.975 21.885 82.975 20.065 82.975 20.065 75.975
                 19.495 75.975 19.495 76.475 20.065 76.475 20.065 79.475 19.495 79.475
                 19.495 79.975 20.065 79.975 20.065 82.975 18.245 82.975 18.245 75.975
                 17.675 75.975 17.675 76.475 18.245 76.475 18.245 79.475 17.675 79.475
                 17.675 79.975 18.245 79.975 18.245 82.975 16.425 82.975 16.425 75.975
                 15.855 75.975 15.855 76.475 16.425 76.475 16.425 79.475 15.855 79.475
                 15.855 79.975 16.425 79.975 16.425 82.975 14.605 82.975 14.605 75.975
                 14.035 75.975 14.035 76.475 14.605 76.475 14.605 79.475 14.035 79.475
                 14.035 79.975 14.605 79.975 14.605 82.975 12.785 82.975 12.785 75.975
                 12.215 75.975 12.215 76.475 12.785 76.475 12.785 79.475 12.215 79.475
                 12.215 79.975 12.785 79.975 12.785 82.975 10.965 82.975 10.965 75.975
                 10.395 75.975 10.395 76.475 10.965 76.475 10.965 79.475 10.395 79.475
                 10.395 79.975 10.965 79.975 10.965 82.975 9.145 82.975 9.145 75.975
                 8.575 75.975 8.575 76.475 9.145 76.475 9.145 79.475 8.575 79.475
                 8.575 79.975 9.145 79.975 9.145 82.975 7.325 82.975 7.325 75.975
                 6.755 75.975 6.755 76.475 7.325 76.475 7.325 79.475 6.755 79.475
                 6.755 79.975 7.325 79.975 7.325 82.975 5.505 82.975 5.505 75.975
                 4.935 75.975 4.935 76.475 5.505 76.475 5.505 79.475 4.935 79.475
                 4.935 79.975 5.505 79.975 5.505 82.975 3.685 82.975 3.685 75.975
                 3.115 75.975 3.115 76.475 3.685 76.475 3.685 79.475 3.115 79.475
                 3.115 79.975 3.685 79.975 3.685 82.975 0.000 82.975 0.000 79.975
                 1.865 79.975 1.865 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  24.085 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.135 72.475 25.000 75.975 ;
        RECT  23.135 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  0.000 118.010 25.000 118.500 ;
        RECT  23.755 39.450 24.085 44.475 ;
        RECT  13.880 40.975 23.755 44.475 ;
        RECT  21.885 72.475 23.135 82.975 ;
        RECT  21.315 72.475 21.885 75.975 ;
        RECT  21.315 76.475 21.885 79.475 ;
        RECT  21.315 79.975 21.885 82.975 ;
        RECT  20.065 72.475 21.315 82.975 ;
        RECT  19.495 72.475 20.065 75.975 ;
        RECT  19.495 76.475 20.065 79.475 ;
        RECT  19.495 79.975 20.065 82.975 ;
        RECT  18.245 72.475 19.495 82.975 ;
        RECT  17.675 72.475 18.245 75.975 ;
        RECT  17.675 76.475 18.245 79.475 ;
        RECT  17.675 79.975 18.245 82.975 ;
        RECT  16.425 72.475 17.675 82.975 ;
        RECT  15.855 72.475 16.425 75.975 ;
        RECT  15.855 76.475 16.425 79.475 ;
        RECT  15.855 79.975 16.425 82.975 ;
        RECT  14.605 72.475 15.855 82.975 ;
        RECT  14.035 72.475 14.605 75.975 ;
        RECT  14.035 76.475 14.605 79.475 ;
        RECT  14.035 79.975 14.605 82.975 ;
        RECT  13.880 72.475 14.035 82.975 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  12.785 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  12.215 40.975 12.785 75.975 ;
        RECT  12.215 76.475 12.785 79.475 ;
        RECT  12.215 79.975 12.785 82.975 ;
        RECT  11.120 40.975 12.215 82.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.245 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.965 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.395 72.475 10.965 75.975 ;
        RECT  10.395 76.475 10.965 79.475 ;
        RECT  10.395 79.975 10.965 82.975 ;
        RECT  9.145 72.475 10.395 82.975 ;
        RECT  8.575 72.475 9.145 75.975 ;
        RECT  8.575 76.475 9.145 79.475 ;
        RECT  8.575 79.975 9.145 82.975 ;
        RECT  7.325 72.475 8.575 82.975 ;
        RECT  6.755 72.475 7.325 75.975 ;
        RECT  6.755 76.475 7.325 79.475 ;
        RECT  6.755 79.975 7.325 82.975 ;
        RECT  5.505 72.475 6.755 82.975 ;
        RECT  4.935 72.475 5.505 75.975 ;
        RECT  4.935 76.475 5.505 79.475 ;
        RECT  4.935 79.975 5.505 82.975 ;
        RECT  3.685 72.475 4.935 82.975 ;
        RECT  3.115 72.475 3.685 75.975 ;
        RECT  3.115 76.475 3.685 79.475 ;
        RECT  3.115 79.975 3.685 82.975 ;
        RECT  1.865 72.475 3.115 82.975 ;
        RECT  0.000 72.475 1.865 75.975 ;
        RECT  0.000 79.975 1.865 82.975 ;
        RECT  0.915 39.450 1.245 44.475 ;
        RECT  0.000 40.975 0.915 44.475 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  24.085 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.135 72.475 25.000 75.975 ;
        RECT  23.135 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  23.755 39.450 24.085 44.475 ;
        RECT  13.880 40.975 23.755 44.475 ;
        RECT  21.885 72.475 23.135 82.975 ;
        RECT  21.315 72.475 21.885 75.975 ;
        RECT  21.315 76.475 21.885 79.475 ;
        RECT  21.315 79.975 21.885 82.975 ;
        RECT  20.065 72.475 21.315 82.975 ;
        RECT  19.495 72.475 20.065 75.975 ;
        RECT  19.495 76.475 20.065 79.475 ;
        RECT  19.495 79.975 20.065 82.975 ;
        RECT  18.245 72.475 19.495 82.975 ;
        RECT  17.675 72.475 18.245 75.975 ;
        RECT  17.675 76.475 18.245 79.475 ;
        RECT  17.675 79.975 18.245 82.975 ;
        RECT  16.425 72.475 17.675 82.975 ;
        RECT  15.855 72.475 16.425 75.975 ;
        RECT  15.855 76.475 16.425 79.475 ;
        RECT  15.855 79.975 16.425 82.975 ;
        RECT  14.605 72.475 15.855 82.975 ;
        RECT  14.035 72.475 14.605 75.975 ;
        RECT  14.035 76.475 14.605 79.475 ;
        RECT  14.035 79.975 14.605 82.975 ;
        RECT  13.880 72.475 14.035 82.975 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  12.785 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  12.215 40.975 12.785 75.975 ;
        RECT  12.215 76.475 12.785 79.475 ;
        RECT  12.215 79.975 12.785 82.975 ;
        RECT  11.120 40.975 12.215 82.975 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  1.245 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.965 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.395 72.475 10.965 75.975 ;
        RECT  10.395 76.475 10.965 79.475 ;
        RECT  10.395 79.975 10.965 82.975 ;
        RECT  9.145 72.475 10.395 82.975 ;
        RECT  8.575 72.475 9.145 75.975 ;
        RECT  8.575 76.475 9.145 79.475 ;
        RECT  8.575 79.975 9.145 82.975 ;
        RECT  7.325 72.475 8.575 82.975 ;
        RECT  6.755 72.475 7.325 75.975 ;
        RECT  6.755 76.475 7.325 79.475 ;
        RECT  6.755 79.975 7.325 82.975 ;
        RECT  5.505 72.475 6.755 82.975 ;
        RECT  4.935 72.475 5.505 75.975 ;
        RECT  4.935 76.475 5.505 79.475 ;
        RECT  4.935 79.975 5.505 82.975 ;
        RECT  3.685 72.475 4.935 82.975 ;
        RECT  3.115 72.475 3.685 75.975 ;
        RECT  3.115 76.475 3.685 79.475 ;
        RECT  3.115 79.975 3.685 82.975 ;
        RECT  1.865 72.475 3.115 82.975 ;
        RECT  0.000 72.475 1.865 75.975 ;
        RECT  0.000 79.975 1.865 82.975 ;
        RECT  0.915 39.450 1.245 44.475 ;
        RECT  0.000 40.975 0.915 44.475 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD2POC_G

MACRO PVDD3AC_G
    CLASS PAD ;
    FOREIGN PVDD3AC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TACVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TACVSS
    PIN TACVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M6 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M5 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M4 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M3 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 23.035 75.975 23.035 79.975 25.000 79.975 25.000 82.975
                 22.485 82.975 22.485 75.975 21.955 75.975 21.955 76.475 22.485 76.475
                 22.485 79.475 21.955 79.475 21.955 79.975 22.485 79.975 22.485 82.975
                 21.405 82.975 21.405 75.975 20.875 75.975 20.875 76.475 21.405 76.475
                 21.405 79.475 20.875 79.475 20.875 79.975 21.405 79.975 21.405 82.975
                 20.325 82.975 20.325 75.975 19.795 75.975 19.795 76.475 20.325 76.475
                 20.325 79.475 19.795 79.475 19.795 79.975 20.325 79.975 20.325 82.975
                 19.245 82.975 19.245 75.975 18.715 75.975 18.715 76.475 19.245 76.475
                 19.245 79.475 18.715 79.475 18.715 79.975 19.245 79.975 19.245 82.975
                 18.165 82.975 18.165 75.975 17.635 75.975 17.635 76.475 18.165 76.475
                 18.165 79.475 17.635 79.475 17.635 79.975 18.165 79.975 18.165 82.975
                 17.085 82.975 17.085 75.975 16.555 75.975 16.555 76.475 17.085 76.475
                 17.085 79.475 16.555 79.475 16.555 79.975 17.085 79.975 17.085 82.975
                 16.005 82.975 16.005 75.975 15.475 75.975 15.475 76.475 16.005 76.475
                 16.005 79.475 15.475 79.475 15.475 79.975 16.005 79.975 16.005 82.975
                 14.925 82.975 14.925 75.975 14.395 75.975 14.395 76.475 14.925 76.475
                 14.925 79.475 14.395 79.475 14.395 79.975 14.925 79.975 14.925 82.975
                 13.845 82.975 13.845 75.975 13.315 75.975 13.315 76.475 13.845 76.475
                 13.845 79.475 13.315 79.475 13.315 79.975 13.845 79.975 13.845 82.975
                 12.765 82.975 12.765 75.975 12.235 75.975 12.235 76.475 12.765 76.475
                 12.765 79.475 12.235 79.475 12.235 79.975 12.765 79.975 12.765 82.975
                 11.685 82.975 11.685 75.975 11.155 75.975 11.155 76.475 11.685 76.475
                 11.685 79.475 11.155 79.475 11.155 79.975 11.685 79.975 11.685 82.975
                 10.605 82.975 10.605 75.975 10.075 75.975 10.075 76.475 10.605 76.475
                 10.605 79.475 10.075 79.475 10.075 79.975 10.605 79.975 10.605 82.975
                 9.525 82.975 9.525 75.975 8.995 75.975 8.995 76.475 9.525 76.475
                 9.525 79.475 8.995 79.475 8.995 79.975 9.525 79.975 9.525 82.975
                 8.445 82.975 8.445 75.975 7.915 75.975 7.915 76.475 8.445 76.475
                 8.445 79.475 7.915 79.475 7.915 79.975 8.445 79.975 8.445 82.975
                 7.365 82.975 7.365 75.975 6.835 75.975 6.835 76.475 7.365 76.475
                 7.365 79.475 6.835 79.475 6.835 79.975 7.365 79.975 7.365 82.975
                 6.285 82.975 6.285 75.975 5.755 75.975 5.755 76.475 6.285 76.475
                 6.285 79.475 5.755 79.475 5.755 79.975 6.285 79.975 6.285 82.975
                 5.205 82.975 5.205 75.975 4.675 75.975 4.675 76.475 5.205 76.475
                 5.205 79.475 4.675 79.475 4.675 79.975 5.205 79.975 5.205 82.975
                 4.125 82.975 4.125 75.975 3.595 75.975 3.595 76.475 4.125 76.475
                 4.125 79.475 3.595 79.475 3.595 79.975 4.125 79.975 4.125 82.975
                 3.045 82.975 3.045 75.975 2.515 75.975 2.515 76.475 3.045 76.475
                 3.045 79.475 2.515 79.475 2.515 79.975 3.045 79.975 3.045 82.975
                 0.000 82.975 0.000 79.975 1.965 79.975 1.965 75.975 0.000 75.975
                 0.000 72.475 11.120 72.475 11.120 71.475 0.000 71.475 0.000 67.975
                 11.120 67.975 11.120 66.975 0.000 66.975 0.000 63.475 11.120 63.475
                 11.120 62.475 0.000 62.475 0.000 58.975 11.120 58.975 11.120 57.975
                 0.000 57.975 0.000 54.475 11.120 54.475 11.120 53.475 0.000 53.475
                 0.000 49.975 11.120 49.975 11.120 48.975 0.000 48.975 0.000 45.475
                 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TACVDD
    PIN AVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.965 118.255 3.595 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  4.125 118.255 5.755 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  6.285 118.255 7.915 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.445 118.255 10.075 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  10.605 118.255 12.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  12.765 118.255 14.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.925 118.255 16.555 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  17.085 118.255 18.715 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  19.245 118.255 20.875 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.405 118.255 23.035 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.965 118.255 3.595 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  4.125 118.255 5.755 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.285 118.255 7.915 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.445 118.255 10.075 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  10.605 118.255 12.235 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  12.765 118.255 14.395 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.925 118.255 16.555 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  17.085 118.255 18.715 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  19.245 118.255 20.875 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.405 118.255 23.035 120 ;
        END
        PORT
        LAYER M2 ;
        RECT  21.405 118.255 23.035 120.000 ;
        RECT  19.245 118.255 20.875 120.000 ;
        RECT  17.085 118.255 18.715 120.000 ;
        RECT  14.925 118.255 16.555 120.000 ;
        RECT  12.765 118.255 14.395 120.000 ;
        RECT  10.605 118.255 12.235 120.000 ;
        RECT  8.445 118.255 10.075 120.000 ;
        RECT  6.285 118.255 7.915 120.000 ;
        RECT  4.125 118.255 5.755 120.000 ;
        RECT  1.965 118.255 3.595 120.000 ;
        LAYER M1 ;
        RECT  21.405 118.255 23.035 120.000 ;
        RECT  19.245 118.255 20.875 120.000 ;
        RECT  17.085 118.255 18.715 120.000 ;
        RECT  14.925 118.255 16.555 120.000 ;
        RECT  12.765 118.255 14.395 120.000 ;
        RECT  10.605 118.255 12.235 120.000 ;
        RECT  8.445 118.255 10.075 120.000 ;
        RECT  6.285 118.255 7.915 120.000 ;
        RECT  4.125 118.255 5.755 120.000 ;
        RECT  1.965 118.255 3.595 120.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.405 118.255 23.035 120.000 ;
        RECT  19.245 118.255 20.875 120.000 ;
        RECT  17.085 118.255 18.715 120.000 ;
        RECT  14.925 118.255 16.555 120.000 ;
        RECT  12.765 118.255 14.395 120.000 ;
        RECT  10.605 118.255 12.235 120.000 ;
        RECT  8.445 118.255 10.075 120.000 ;
        RECT  6.285 118.255 7.915 120.000 ;
        RECT  4.125 118.255 5.755 120.000 ;
        RECT  1.965 118.255 3.595 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.035 72.475 25.000 75.975 ;
        RECT  23.035 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.485 72.475 23.035 82.975 ;
        RECT  21.955 72.475 22.485 75.975 ;
        RECT  21.955 76.475 22.485 79.475 ;
        RECT  21.955 79.975 22.485 82.975 ;
        RECT  21.405 72.475 21.955 82.975 ;
        RECT  20.875 72.475 21.405 75.975 ;
        RECT  20.875 76.475 21.405 79.475 ;
        RECT  20.875 79.975 21.405 82.975 ;
        RECT  20.325 72.475 20.875 82.975 ;
        RECT  19.795 72.475 20.325 75.975 ;
        RECT  19.795 76.475 20.325 79.475 ;
        RECT  19.795 79.975 20.325 82.975 ;
        RECT  19.245 72.475 19.795 82.975 ;
        RECT  18.715 72.475 19.245 75.975 ;
        RECT  18.715 76.475 19.245 79.475 ;
        RECT  18.715 79.975 19.245 82.975 ;
        RECT  18.165 72.475 18.715 82.975 ;
        RECT  17.635 72.475 18.165 75.975 ;
        RECT  17.635 76.475 18.165 79.475 ;
        RECT  17.635 79.975 18.165 82.975 ;
        RECT  17.085 72.475 17.635 82.975 ;
        RECT  16.555 72.475 17.085 75.975 ;
        RECT  16.555 76.475 17.085 79.475 ;
        RECT  16.555 79.975 17.085 82.975 ;
        RECT  16.005 72.475 16.555 82.975 ;
        RECT  15.475 72.475 16.005 75.975 ;
        RECT  15.475 76.475 16.005 79.475 ;
        RECT  15.475 79.975 16.005 82.975 ;
        RECT  14.925 72.475 15.475 82.975 ;
        RECT  14.395 72.475 14.925 75.975 ;
        RECT  14.395 76.475 14.925 79.475 ;
        RECT  14.395 79.975 14.925 82.975 ;
        RECT  13.880 72.475 14.395 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.845 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  13.315 40.975 13.845 75.975 ;
        RECT  13.315 76.475 13.845 79.475 ;
        RECT  13.315 79.975 13.845 82.975 ;
        RECT  12.765 40.975 13.315 82.975 ;
        RECT  12.235 40.975 12.765 75.975 ;
        RECT  12.235 76.475 12.765 79.475 ;
        RECT  12.235 79.975 12.765 82.975 ;
        RECT  11.685 40.975 12.235 82.975 ;
        RECT  11.155 40.975 11.685 75.975 ;
        RECT  11.155 76.475 11.685 79.475 ;
        RECT  11.155 79.975 11.685 82.975 ;
        RECT  11.120 40.975 11.155 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.605 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.075 72.475 10.605 75.975 ;
        RECT  10.075 76.475 10.605 79.475 ;
        RECT  10.075 79.975 10.605 82.975 ;
        RECT  9.525 72.475 10.075 82.975 ;
        RECT  8.995 72.475 9.525 75.975 ;
        RECT  8.995 76.475 9.525 79.475 ;
        RECT  8.995 79.975 9.525 82.975 ;
        RECT  8.445 72.475 8.995 82.975 ;
        RECT  7.915 72.475 8.445 75.975 ;
        RECT  7.915 76.475 8.445 79.475 ;
        RECT  7.915 79.975 8.445 82.975 ;
        RECT  7.365 72.475 7.915 82.975 ;
        RECT  6.835 72.475 7.365 75.975 ;
        RECT  6.835 76.475 7.365 79.475 ;
        RECT  6.835 79.975 7.365 82.975 ;
        RECT  6.285 72.475 6.835 82.975 ;
        RECT  5.755 72.475 6.285 75.975 ;
        RECT  5.755 76.475 6.285 79.475 ;
        RECT  5.755 79.975 6.285 82.975 ;
        RECT  5.205 72.475 5.755 82.975 ;
        RECT  4.675 72.475 5.205 75.975 ;
        RECT  4.675 76.475 5.205 79.475 ;
        RECT  4.675 79.975 5.205 82.975 ;
        RECT  4.125 72.475 4.675 82.975 ;
        RECT  3.595 72.475 4.125 75.975 ;
        RECT  3.595 76.475 4.125 79.475 ;
        RECT  3.595 79.975 4.125 82.975 ;
        RECT  3.045 72.475 3.595 82.975 ;
        RECT  2.515 72.475 3.045 75.975 ;
        RECT  2.515 76.475 3.045 79.475 ;
        RECT  2.515 79.975 3.045 82.975 ;
        RECT  1.965 72.475 2.515 82.975 ;
        RECT  0.000 72.475 1.965 75.975 ;
        RECT  0.000 79.975 1.965 82.975 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.035 72.475 25.000 75.975 ;
        RECT  23.035 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.485 72.475 23.035 82.975 ;
        RECT  22.265 72.475 22.485 75.975 ;
        RECT  22.265 76.475 22.485 79.475 ;
        RECT  22.265 79.975 22.485 82.975 ;
        RECT  20.325 72.475 22.265 82.975 ;
        RECT  19.795 72.475 20.325 75.975 ;
        RECT  19.795 76.475 20.325 79.475 ;
        RECT  19.795 79.975 20.325 82.975 ;
        RECT  17.765 72.475 19.795 82.975 ;
        RECT  17.635 72.475 17.765 75.975 ;
        RECT  17.635 76.475 17.765 79.475 ;
        RECT  17.635 79.975 17.765 82.975 ;
        RECT  17.085 72.475 17.635 82.975 ;
        RECT  16.555 72.475 17.085 75.975 ;
        RECT  16.555 76.475 17.085 79.475 ;
        RECT  16.555 79.975 17.085 82.975 ;
        RECT  14.765 72.475 16.555 82.975 ;
        RECT  14.395 72.475 14.765 75.975 ;
        RECT  14.395 76.475 14.765 79.475 ;
        RECT  14.395 79.975 14.765 82.975 ;
        RECT  13.880 72.475 14.395 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.845 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  13.315 40.975 13.845 75.975 ;
        RECT  13.315 76.475 13.845 79.475 ;
        RECT  13.315 79.975 13.845 82.975 ;
        RECT  11.685 40.975 13.315 82.975 ;
        RECT  11.155 40.975 11.685 75.975 ;
        RECT  11.155 76.475 11.685 79.475 ;
        RECT  11.155 79.975 11.685 82.975 ;
        RECT  11.120 40.975 11.155 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.605 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.265 72.475 10.605 75.975 ;
        RECT  10.265 76.475 10.605 79.475 ;
        RECT  10.265 79.975 10.605 82.975 ;
        RECT  8.445 72.475 10.265 82.975 ;
        RECT  7.915 72.475 8.445 75.975 ;
        RECT  7.915 76.475 8.445 79.475 ;
        RECT  7.915 79.975 8.445 82.975 ;
        RECT  7.365 72.475 7.915 82.975 ;
        RECT  7.265 72.475 7.365 75.975 ;
        RECT  7.265 76.475 7.365 79.475 ;
        RECT  7.265 79.975 7.365 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  5.755 72.475 5.765 75.975 ;
        RECT  5.755 76.475 5.765 79.475 ;
        RECT  5.755 79.975 5.765 82.975 ;
        RECT  5.205 72.475 5.755 82.975 ;
        RECT  4.675 72.475 5.205 75.975 ;
        RECT  4.675 76.475 5.205 79.475 ;
        RECT  4.675 79.975 5.205 82.975 ;
        RECT  2.765 72.475 4.675 82.975 ;
        RECT  2.515 72.475 2.765 75.975 ;
        RECT  2.515 76.475 2.765 79.475 ;
        RECT  2.515 79.975 2.765 82.975 ;
        RECT  1.965 72.475 2.515 82.975 ;
        RECT  0.000 72.475 1.965 75.975 ;
        RECT  0.000 79.975 1.965 82.975 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD3AC_G

MACRO PVDD3A_G
    CLASS PAD ;
    FOREIGN PVDD3A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M6 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M5 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M4 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 22.265 75.975 22.265 76.475 22.615 76.475 22.615 79.475
                 22.265 79.475 22.265 79.975 25.000 79.975 25.000 82.975 20.765 82.975
                 20.765 75.975 19.265 75.975 19.265 76.475 20.765 76.475 20.765 79.475
                 19.265 79.475 19.265 79.975 20.765 79.975 20.765 82.975 17.765 82.975
                 17.765 75.975 16.265 75.975 16.265 76.475 17.765 76.475 17.765 79.475
                 16.265 79.475 16.265 79.975 17.765 79.975 17.765 82.975 14.765 82.975
                 14.765 75.975 13.265 75.975 13.265 76.475 14.765 76.475 14.765 79.475
                 13.265 79.475 13.265 79.975 14.765 79.975 14.765 82.975 11.765 82.975
                 11.765 75.975 10.265 75.975 10.265 76.475 11.765 76.475 11.765 79.475
                 10.265 79.475 10.265 79.975 11.765 79.975 11.765 82.975 8.765 82.975
                 8.765 75.975 7.265 75.975 7.265 76.475 8.765 76.475 8.765 79.475
                 7.265 79.475 7.265 79.975 8.765 79.975 8.765 82.975 5.765 82.975
                 5.765 75.975 4.265 75.975 4.265 76.475 5.765 76.475 5.765 79.475
                 4.265 79.475 4.265 79.975 5.765 79.975 5.765 82.975 0.000 82.975
                 0.000 79.975 2.765 79.975 2.765 79.475 2.385 79.475 2.385 76.475
                 2.765 76.475 2.765 75.975 0.000 75.975 0.000 72.475 11.120 72.475
                 11.120 71.475 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975
                 0.000 66.975 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475
                 0.000 58.975 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475
                 11.120 54.475 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975
                 11.120 48.975 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475
                 0.000 44.475 ;
        LAYER M3 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 23.120 75.975 23.120 79.975 25.000 79.975 25.000 82.975
                 22.120 82.975 22.120 75.975 21.280 75.975 21.280 76.475 22.120 76.475
                 22.120 79.475 21.280 79.475 21.280 79.975 22.120 79.975 22.120 82.975
                 20.280 82.975 20.280 75.975 19.440 75.975 19.440 76.475 20.280 76.475
                 20.280 79.475 19.440 79.475 19.440 79.975 20.280 79.975 20.280 82.975
                 18.440 82.975 18.440 75.975 17.600 75.975 17.600 76.475 18.440 76.475
                 18.440 79.475 17.600 79.475 17.600 79.975 18.440 79.975 18.440 82.975
                 16.600 82.975 16.600 75.975 15.760 75.975 15.760 76.475 16.600 76.475
                 16.600 79.475 15.760 79.475 15.760 79.975 16.600 79.975 16.600 82.975
                 14.760 82.975 14.760 75.975 13.920 75.975 13.920 76.475 14.760 76.475
                 14.760 79.475 13.920 79.475 13.920 79.975 14.760 79.975 14.760 82.975
                 12.920 82.975 12.920 75.975 12.080 75.975 12.080 76.475 12.920 76.475
                 12.920 79.475 12.080 79.475 12.080 79.975 12.920 79.975 12.920 82.975
                 11.080 82.975 11.080 75.975 10.240 75.975 10.240 76.475 11.080 76.475
                 11.080 79.475 10.240 79.475 10.240 79.975 11.080 79.975 11.080 82.975
                 9.240 82.975 9.240 75.975 8.400 75.975 8.400 76.475 9.240 76.475
                 9.240 79.475 8.400 79.475 8.400 79.975 9.240 79.975 9.240 82.975
                 7.400 82.975 7.400 75.975 6.560 75.975 6.560 76.475 7.400 76.475
                 7.400 79.475 6.560 79.475 6.560 79.975 7.400 79.975 7.400 82.975
                 5.560 82.975 5.560 75.975 4.720 75.975 4.720 76.475 5.560 76.475
                 5.560 79.475 4.720 79.475 4.720 79.975 5.560 79.975 5.560 82.975
                 3.720 82.975 3.720 75.975 2.880 75.975 2.880 76.475 3.720 76.475
                 3.720 79.475 2.880 79.475 2.880 79.975 3.720 79.975 3.720 82.975
                 0.000 82.975 0.000 79.975 1.880 79.975 1.880 75.975 0.000 75.975
                 0.000 72.475 11.120 72.475 11.120 71.475 0.000 71.475 0.000 67.975
                 11.120 67.975 11.120 66.975 0.000 66.975 0.000 63.475 11.120 63.475
                 11.120 62.475 0.000 62.475 0.000 58.975 11.120 58.975 11.120 57.975
                 0.000 57.975 0.000 54.475 11.120 54.475 11.120 53.475 0.000 53.475
                 0.000 49.975 11.120 49.975 11.120 48.975 0.000 48.975 0.000 45.475
                 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TAVDD
    PIN AVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.91 118.255 3.41 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.19 118.255 6.69 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.47 118.255 9.97 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.75 118.255 13.25 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.03 118.255 16.53 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  18.31 118.255 19.81 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.59 118.255 23.09 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.73 118.255 3.59 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.01 118.255 6.87 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.29 118.255 10.15 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.57 118.255 13.43 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.85 118.255 16.71 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  18.13 118.255 19.99 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.41 118.255 23.27 120 ;
        END
        PORT
        LAYER M2 ;
        RECT  21.410 118.255 23.270 120.000 ;
        RECT  18.130 118.255 19.990 120.000 ;
        RECT  14.850 118.255 16.710 120.000 ;
        RECT  11.570 118.255 13.430 120.000 ;
        RECT  8.290 118.255 10.150 120.000 ;
        RECT  5.010 118.255 6.870 120.000 ;
        RECT  1.730 118.255 3.590 120.000 ;
        LAYER M1 ;
        RECT  21.590 118.255 23.090 120.000 ;
        RECT  18.310 118.255 19.810 120.000 ;
        RECT  15.030 118.255 16.530 120.000 ;
        RECT  11.750 118.255 13.250 120.000 ;
        RECT  8.470 118.255 9.970 120.000 ;
        RECT  5.190 118.255 6.690 120.000 ;
        RECT  1.910 118.255 3.410 120.000 ;
        END
    END AVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.410 118.255 23.270 120.000 ;
        RECT  18.130 118.255 19.990 120.000 ;
        RECT  14.850 118.255 16.710 120.000 ;
        RECT  11.570 118.255 13.430 120.000 ;
        RECT  8.290 118.255 10.150 120.000 ;
        RECT  5.010 118.255 6.870 120.000 ;
        RECT  1.730 118.255 3.590 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.120 72.475 25.000 75.975 ;
        RECT  23.120 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.120 72.475 23.120 82.975 ;
        RECT  21.280 72.475 22.120 75.975 ;
        RECT  21.280 76.475 22.120 79.475 ;
        RECT  21.280 79.975 22.120 82.975 ;
        RECT  20.280 72.475 21.280 82.975 ;
        RECT  19.440 72.475 20.280 75.975 ;
        RECT  19.440 76.475 20.280 79.475 ;
        RECT  19.440 79.975 20.280 82.975 ;
        RECT  18.440 72.475 19.440 82.975 ;
        RECT  17.600 72.475 18.440 75.975 ;
        RECT  17.600 76.475 18.440 79.475 ;
        RECT  17.600 79.975 18.440 82.975 ;
        RECT  16.600 72.475 17.600 82.975 ;
        RECT  15.760 72.475 16.600 75.975 ;
        RECT  15.760 76.475 16.600 79.475 ;
        RECT  15.760 79.975 16.600 82.975 ;
        RECT  14.760 72.475 15.760 82.975 ;
        RECT  13.920 72.475 14.760 75.975 ;
        RECT  13.920 76.475 14.760 79.475 ;
        RECT  13.920 79.975 14.760 82.975 ;
        RECT  13.880 72.475 13.920 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  12.920 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  12.080 40.975 12.920 75.975 ;
        RECT  12.080 76.475 12.920 79.475 ;
        RECT  12.080 79.975 12.920 82.975 ;
        RECT  11.120 40.975 12.080 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  11.080 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.240 72.475 11.080 75.975 ;
        RECT  10.240 76.475 11.080 79.475 ;
        RECT  10.240 79.975 11.080 82.975 ;
        RECT  9.240 72.475 10.240 82.975 ;
        RECT  8.400 72.475 9.240 75.975 ;
        RECT  8.400 76.475 9.240 79.475 ;
        RECT  8.400 79.975 9.240 82.975 ;
        RECT  7.400 72.475 8.400 82.975 ;
        RECT  6.560 72.475 7.400 75.975 ;
        RECT  6.560 76.475 7.400 79.475 ;
        RECT  6.560 79.975 7.400 82.975 ;
        RECT  5.560 72.475 6.560 82.975 ;
        RECT  4.720 72.475 5.560 75.975 ;
        RECT  4.720 76.475 5.560 79.475 ;
        RECT  4.720 79.975 5.560 82.975 ;
        RECT  3.720 72.475 4.720 82.975 ;
        RECT  2.880 72.475 3.720 75.975 ;
        RECT  2.880 76.475 3.720 79.475 ;
        RECT  2.880 79.975 3.720 82.975 ;
        RECT  1.880 72.475 2.880 82.975 ;
        RECT  0.000 72.475 1.880 75.975 ;
        RECT  0.000 79.975 1.880 82.975 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  23.120 72.475 25.000 75.975 ;
        RECT  23.120 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  20.280 72.475 23.120 82.975 ;
        RECT  19.440 72.475 20.280 75.975 ;
        RECT  19.440 76.475 20.280 79.475 ;
        RECT  19.440 79.975 20.280 82.975 ;
        RECT  17.765 72.475 19.440 82.975 ;
        RECT  17.600 72.475 17.765 75.975 ;
        RECT  17.600 76.475 17.765 79.475 ;
        RECT  17.600 79.975 17.765 82.975 ;
        RECT  16.600 72.475 17.600 82.975 ;
        RECT  16.265 72.475 16.600 75.975 ;
        RECT  16.265 76.475 16.600 79.475 ;
        RECT  16.265 79.975 16.600 82.975 ;
        RECT  14.760 72.475 16.265 82.975 ;
        RECT  13.920 72.475 14.760 75.975 ;
        RECT  13.920 76.475 14.760 79.475 ;
        RECT  13.920 79.975 14.760 82.975 ;
        RECT  13.880 72.475 13.920 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 82.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  11.080 72.475 11.120 82.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  10.265 72.475 11.080 75.975 ;
        RECT  10.265 76.475 11.080 79.475 ;
        RECT  10.265 79.975 11.080 82.975 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  8.400 72.475 8.765 75.975 ;
        RECT  8.400 76.475 8.765 79.475 ;
        RECT  8.400 79.975 8.765 82.975 ;
        RECT  7.400 72.475 8.400 82.975 ;
        RECT  7.265 72.475 7.400 75.975 ;
        RECT  7.265 76.475 7.400 79.475 ;
        RECT  7.265 79.975 7.400 82.975 ;
        RECT  5.560 72.475 7.265 82.975 ;
        RECT  4.720 72.475 5.560 75.975 ;
        RECT  4.720 76.475 5.560 79.475 ;
        RECT  4.720 79.975 5.560 82.975 ;
        RECT  1.880 72.475 4.720 82.975 ;
        RECT  0.000 72.475 1.880 75.975 ;
        RECT  0.000 79.975 1.880 82.975 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  22.265 72.475 25.000 75.975 ;
        RECT  22.265 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  22.265 76.475 22.615 79.475 ;
        RECT  20.765 72.475 22.265 82.975 ;
        RECT  19.265 72.475 20.765 75.975 ;
        RECT  19.265 76.475 20.765 79.475 ;
        RECT  19.265 79.975 20.765 82.975 ;
        RECT  17.765 72.475 19.265 82.975 ;
        RECT  16.265 72.475 17.765 75.975 ;
        RECT  16.265 76.475 17.765 79.475 ;
        RECT  16.265 79.975 17.765 82.975 ;
        RECT  14.765 72.475 16.265 82.975 ;
        RECT  13.880 72.475 14.765 75.975 ;
        RECT  13.265 76.475 14.765 79.475 ;
        RECT  13.265 79.975 14.765 82.975 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  13.265 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  11.765 40.975 13.265 82.975 ;
        RECT  11.120 40.975 11.765 75.975 ;
        RECT  10.265 76.475 11.765 79.475 ;
        RECT  10.265 79.975 11.765 82.975 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  10.265 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        RECT  8.765 72.475 10.265 82.975 ;
        RECT  7.265 72.475 8.765 75.975 ;
        RECT  7.265 76.475 8.765 79.475 ;
        RECT  7.265 79.975 8.765 82.975 ;
        RECT  5.765 72.475 7.265 82.975 ;
        RECT  4.265 72.475 5.765 75.975 ;
        RECT  4.265 76.475 5.765 79.475 ;
        RECT  4.265 79.975 5.765 82.975 ;
        RECT  2.765 72.475 4.265 82.975 ;
        RECT  0.000 72.475 2.765 75.975 ;
        RECT  2.385 76.475 2.765 79.475 ;
        RECT  0.000 79.975 2.765 82.975 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVDD3A_G

MACRO PVSS1ANA_G
    CLASS PAD ;
    FOREIGN PVSS1ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    PIN AVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.97 118.5 3.77 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.18 118.5 6.98 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.39 118.5 10.19 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.6 118.5 13.4 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.81 118.5 16.61 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  18.02 118.5 19.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.23 118.5 23.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.97 118.5 3.77 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.18 118.5 6.98 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.39 118.5 10.19 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.6 118.5 13.4 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.81 118.5 16.61 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  18.02 118.5 19.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.23 118.5 23.03 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  1.920 76.475 23.080 79.475 ;
        LAYER M2 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        LAYER M1 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS1ANA_G

MACRO PVSS1DGZ_G
    CLASS PAD ;
    FOREIGN PVSS1DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.92 118.5 3.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.13 118.5 7.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.34 118.5 10.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.55 118.5 13.45 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.76 118.5 16.66 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  17.97 118.5 19.87 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.18 118.5 23.08 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.92 118.5 3.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.13 118.5 7.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.34 118.5 10.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.55 118.5 13.45 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.76 118.5 16.66 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  17.97 118.5 19.87 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.18 118.5 23.08 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
        RECT  1.920 76.475 23.080 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        LAYER M2 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        LAYER M1 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS1DGZ_G

MACRO PVSS2AC_G
    CLASS PAD ;
    FOREIGN PVSS2AC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TACVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TACVSS
    PIN TACVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TACVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS2AC_G

MACRO PVSS2A_G
    CLASS PAD ;
    FOREIGN PVSS2A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TAVDD
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS2A_G

MACRO PVSS2ANA_G
    CLASS PAD ;
    FOREIGN PVSS2ANA_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    PIN AVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.97 118.5 3.77 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.18 118.5 6.98 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.39 118.5 10.19 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.6 118.5 13.4 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.81 118.5 16.61 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  18.02 118.5 19.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.23 118.5 23.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.97 118.5 3.77 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.18 118.5 6.98 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.39 118.5 10.19 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.6 118.5 13.4 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.81 118.5 16.61 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  18.02 118.5 19.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.23 118.5 23.03 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
        LAYER M3 ;
        RECT  1.920 76.475 23.080 79.475 ;
        LAYER M2 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        LAYER M1 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.230 118.500 23.030 120.000 ;
        RECT  18.020 118.500 19.820 120.000 ;
        RECT  14.810 118.500 16.610 120.000 ;
        RECT  11.600 118.500 13.400 120.000 ;
        RECT  8.390 118.500 10.190 120.000 ;
        RECT  5.180 118.500 6.980 120.000 ;
        RECT  1.970 118.500 3.770 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS2ANA_G

MACRO PVSS2DGZ_G
    CLASS PAD ;
    FOREIGN PVSS2DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSSPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        LAYER M3 ;
        RECT  1.920 76.475 23.080 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
        END
    END VSSPST
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS2DGZ_G

MACRO PVSS3AC_G
    CLASS PAD ;
    FOREIGN PVSS3AC_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TACVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TACVSS
    PIN TACVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TACVDD
    PIN AVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  2.38 117.83 4.78 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  6.84 117.83 9.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.3 117.83 13.7 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.76 117.83 18.16 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  20.22 117.83 22.62 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  2.38 117.83 4.78 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.84 117.83 9.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.3 117.83 13.7 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  15.76 117.83 18.16 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  20.22 117.83 22.62 120 ;
        END
        PORT
        LAYER M2 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        LAYER M1 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS3AC_G

MACRO PVSS3A_G
    CLASS PAD ;
    FOREIGN PVSS3A_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        END
    END VSS
    PIN TAVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        LAYER M3 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 5.750 13.880 5.750 13.880 7.250
                 25.000 7.250 25.000 11.750 13.880 11.750 13.880 13.250 25.000 13.250
                 25.000 17.750 13.880 17.750 13.880 19.250 25.000 19.250 25.000 23.750
                 13.880 23.750 13.880 25.250 25.000 25.250 25.000 29.750 13.880 29.750
                 13.880 31.250 25.000 31.250 25.000 35.750 13.880 35.750 13.880 36.750
                 25.000 36.750 25.000 39.290 0.000 39.290 0.000 36.750 11.120 36.750
                 11.120 35.750 0.000 35.750 0.000 31.250 11.120 31.250 11.120 29.750
                 0.000 29.750 0.000 25.250 11.120 25.250 11.120 23.750 0.000 23.750
                 0.000 19.250 11.120 19.250 11.120 17.750 0.000 17.750 0.000 13.250
                 11.120 13.250 11.120 11.750 0.000 11.750 0.000 7.250 11.120 7.250
                 11.120 5.750 0.000 5.750 ;
        END
    END TAVSS
    PIN TAVDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END TAVDD
    PIN AVSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  2.38 117.83 4.78 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  6.84 117.83 9.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.3 117.83 13.7 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  15.76 117.83 18.16 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  20.22 117.83 22.62 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  2.38 117.83 4.78 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  6.84 117.83 9.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.3 117.83 13.7 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  15.76 117.83 18.16 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  20.22 117.83 22.62 120 ;
        END
        PORT
        LAYER M2 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        LAYER M1 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        END
    END AVSS
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  20.220 117.830 22.620 120.000 ;
        RECT  15.760 117.830 18.160 120.000 ;
        RECT  11.300 117.830 13.700 120.000 ;
        RECT  6.840 117.830 9.240 120.000 ;
        RECT  2.380 117.830 4.780 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 5.750 ;
        RECT  13.880 7.250 25.000 11.750 ;
        RECT  13.880 13.250 25.000 17.750 ;
        RECT  13.880 19.250 25.000 23.750 ;
        RECT  13.880 25.250 25.000 29.750 ;
        RECT  13.880 31.250 25.000 35.750 ;
        RECT  13.880 36.750 25.000 39.290 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 39.290 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 5.750 ;
        RECT  0.000 7.250 11.120 11.750 ;
        RECT  0.000 13.250 11.120 17.750 ;
        RECT  0.000 19.250 11.120 23.750 ;
        RECT  0.000 25.250 11.120 29.750 ;
        RECT  0.000 31.250 11.120 35.750 ;
        RECT  0.000 36.750 11.120 39.290 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS3A_G

MACRO PVSS3DGZ_G
    CLASS PAD ;
    FOREIGN PVSS3DGZ_G 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 120.000 ;
    SYMMETRY X Y R90 ;
    SITE pad ;
    PIN VSS
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  1.92 118.5 3.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  5.13 118.5 7.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  8.34 118.5 10.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  11.55 118.5 13.45 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  14.76 118.5 16.66 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  17.97 118.5 19.87 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M1 ;
        RECT  21.18 118.5 23.08 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  1.92 118.5 3.82 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  5.13 118.5 7.03 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  8.34 118.5 10.24 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  11.55 118.5 13.45 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  14.76 118.5 16.66 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  17.97 118.5 19.87 120 ;
        END
        PORT
        CLASS CORE ;
        LAYER M2 ;
        RECT  21.18 118.5 23.08 120 ;
        END
        PORT
        LAYER M7 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M6 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M5 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M4 ;
        RECT  2.385 76.475 22.615 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 13.880 108.920 13.880 109.770 25.000 109.770 25.000 113.270
                 13.880 113.270 13.880 114.010 25.000 114.010 25.000 117.510
                 0.000 117.510 0.000 114.010 11.120 114.010 11.120 113.270 0.000 113.270
                 0.000 109.770 11.120 109.770 11.120 108.920 0.000 108.920 0.000 105.420
                 11.120 105.420 11.120 104.570 0.000 104.570 0.000 101.070 11.120 101.070
                 11.120 100.220 0.000 100.220 0.000 96.720 11.120 96.720 11.120 95.870
                 0.000 95.870 0.000 92.370 11.120 92.370 11.120 91.520 0.000 91.520
                 0.000 88.020 11.120 88.020 11.120 87.170 0.000 87.170 ;
        LAYER M3 ;
        RECT  1.920 76.475 23.080 79.475 ;
                POLYGON  0.000 1.250 25.000 1.250 25.000 4.750 13.880 4.750 13.880 5.750
                 25.000 5.750 25.000 9.250 13.880 9.250 13.880 10.250 25.000 10.250
                 25.000 13.750 13.880 13.750 13.880 14.750 25.000 14.750 25.000 18.250
                 13.880 18.250 13.880 19.250 25.000 19.250 25.000 22.750 13.880 22.750
                 13.880 23.750 25.000 23.750 25.000 27.250 13.880 27.250 13.880 28.250
                 25.000 28.250 25.000 31.750 13.880 31.750 13.880 33.080 25.000 33.080
                 25.000 37.580 0.000 37.580 0.000 33.080 11.120 33.080 11.120 31.750
                 0.000 31.750 0.000 28.250 11.120 28.250 11.120 27.250 0.000 27.250
                 0.000 23.750 11.120 23.750 11.120 22.750 0.000 22.750 0.000 19.250
                 11.120 19.250 11.120 18.250 0.000 18.250 0.000 14.750 11.120 14.750
                 11.120 13.750 0.000 13.750 0.000 10.250 11.120 10.250 11.120 9.250
                 0.000 9.250 0.000 5.750 11.120 5.750 11.120 4.750 0.000 4.750 ;
                POLYGON  0.000 83.670 25.000 83.670 25.000 87.170 13.880 87.170 13.880 88.020
                 25.000 88.020 25.000 91.520 13.880 91.520 13.880 92.370 25.000 92.370
                 25.000 95.870 13.880 95.870 13.880 96.720 25.000 96.720 25.000 100.220
                 13.880 100.220 13.880 101.070 25.000 101.070 25.000 104.570
                 13.880 104.570 13.880 105.420 25.000 105.420 25.000 108.920
                 0.000 108.920 0.000 105.420 11.120 105.420 11.120 104.570 0.000 104.570
                 0.000 101.070 11.120 101.070 11.120 100.220 0.000 100.220 0.000 96.720
                 11.120 96.720 11.120 95.870 0.000 95.870 0.000 92.370 11.120 92.370
                 11.120 91.520 0.000 91.520 0.000 88.020 11.120 88.020 11.120 87.170
                 0.000 87.170 ;
        LAYER M2 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        LAYER M1 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        END
    END VSS
    PIN VDDPST
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M7 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M6 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M5 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M4 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        LAYER M3 ;
        RECT  0.000 79.975 25.000 82.975 ;
                POLYGON  0.000 40.975 25.000 40.975 25.000 44.475 13.880 44.475 13.880 45.475
                 25.000 45.475 25.000 48.975 13.880 48.975 13.880 49.975 25.000 49.975
                 25.000 53.475 13.880 53.475 13.880 54.475 25.000 54.475 25.000 57.975
                 13.880 57.975 13.880 58.975 25.000 58.975 25.000 62.475 13.880 62.475
                 13.880 63.475 25.000 63.475 25.000 66.975 13.880 66.975 13.880 67.975
                 25.000 67.975 25.000 71.475 13.880 71.475 13.880 72.475 25.000 72.475
                 25.000 75.975 0.000 75.975 0.000 72.475 11.120 72.475 11.120 71.475
                 0.000 71.475 0.000 67.975 11.120 67.975 11.120 66.975 0.000 66.975
                 0.000 63.475 11.120 63.475 11.120 62.475 0.000 62.475 0.000 58.975
                 11.120 58.975 11.120 57.975 0.000 57.975 0.000 54.475 11.120 54.475
                 11.120 53.475 0.000 53.475 0.000 49.975 11.120 49.975 11.120 48.975
                 0.000 48.975 0.000 45.475 11.120 45.475 11.120 44.475 0.000 44.475 ;
        END
    END VDDPST
    PIN VDD
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
                POLYGON  0.000 109.770 25.000 109.770 25.000 113.270 13.880 113.270
                 13.880 114.010 25.000 114.010 25.000 117.510 0.000 117.510 0.000 114.010
                 11.120 114.010 11.120 113.270 0.000 113.270 ;
        END
    END VDD
    PIN POC
        SHAPE FEEDTHRU ;
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M3 ;
        RECT  0.000 118.010 25.000 118.500 ;
        END
    END POC
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA1 ;
        RECT  21.180 118.500 23.080 120.000 ;
        RECT  17.970 118.500 19.870 120.000 ;
        RECT  14.760 118.500 16.660 120.000 ;
        RECT  11.550 118.500 13.450 120.000 ;
        RECT  8.340 118.500 10.240 120.000 ;
        RECT  5.130 118.500 7.030 120.000 ;
        RECT  1.920 118.500 3.820 120.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA2 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 108.920 ;
        RECT  11.120 109.770 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M3 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA3 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M4 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA4 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M5 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA5 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M6 ;
        RECT  0.000 0.000 25.000 120.000 ;
        LAYER VIA6 ;
        RECT  13.880 1.250 25.000 4.750 ;
        RECT  13.880 5.750 25.000 9.250 ;
        RECT  13.880 10.250 25.000 13.750 ;
        RECT  13.880 14.750 25.000 18.250 ;
        RECT  13.880 19.250 25.000 22.750 ;
        RECT  13.880 23.750 25.000 27.250 ;
        RECT  13.880 28.250 25.000 31.750 ;
        RECT  13.880 33.080 25.000 37.580 ;
        RECT  13.880 40.975 25.000 44.475 ;
        RECT  13.880 45.475 25.000 48.975 ;
        RECT  13.880 49.975 25.000 53.475 ;
        RECT  13.880 54.475 25.000 57.975 ;
        RECT  13.880 58.975 25.000 62.475 ;
        RECT  13.880 63.475 25.000 66.975 ;
        RECT  13.880 67.975 25.000 71.475 ;
        RECT  13.880 72.475 25.000 75.975 ;
        RECT  0.000 79.975 25.000 82.975 ;
        RECT  13.880 83.670 25.000 87.170 ;
        RECT  13.880 88.020 25.000 91.520 ;
        RECT  13.880 92.370 25.000 95.870 ;
        RECT  13.880 96.720 25.000 100.220 ;
        RECT  13.880 101.070 25.000 104.570 ;
        RECT  13.880 105.420 25.000 108.920 ;
        RECT  13.880 109.770 25.000 113.270 ;
        RECT  13.880 114.010 25.000 117.510 ;
        RECT  11.120 1.250 13.880 37.580 ;
        RECT  11.120 40.975 13.880 75.975 ;
        RECT  11.120 83.670 13.880 117.510 ;
        RECT  0.000 1.250 11.120 4.750 ;
        RECT  0.000 5.750 11.120 9.250 ;
        RECT  0.000 10.250 11.120 13.750 ;
        RECT  0.000 14.750 11.120 18.250 ;
        RECT  0.000 19.250 11.120 22.750 ;
        RECT  0.000 23.750 11.120 27.250 ;
        RECT  0.000 28.250 11.120 31.750 ;
        RECT  0.000 33.080 11.120 37.580 ;
        RECT  0.000 40.975 11.120 44.475 ;
        RECT  0.000 45.475 11.120 48.975 ;
        RECT  0.000 49.975 11.120 53.475 ;
        RECT  0.000 54.475 11.120 57.975 ;
        RECT  0.000 58.975 11.120 62.475 ;
        RECT  0.000 63.475 11.120 66.975 ;
        RECT  0.000 67.975 11.120 71.475 ;
        RECT  0.000 72.475 11.120 75.975 ;
        RECT  0.000 83.670 11.120 87.170 ;
        RECT  0.000 88.020 11.120 91.520 ;
        RECT  0.000 92.370 11.120 95.870 ;
        RECT  0.000 96.720 11.120 100.220 ;
        RECT  0.000 101.070 11.120 104.570 ;
        RECT  0.000 105.420 11.120 108.920 ;
        RECT  0.000 109.770 11.120 113.270 ;
        RECT  0.000 114.010 11.120 117.510 ;
        LAYER M7 ;
        RECT  0.000 0.000 25.000 120.000 ;
    END
END PVSS3DGZ_G

END LIBRARY
