###############################################################################
#TSMC Library/IP Product
#Filename: tpbn45v_ds_9lm.lef
#Technology: N45
#Product Type: I/O PAD
#Product Name: tpbn45v_ds
#Version: 150a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

MACRO PAD50GAU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD50GAU_DS_SL 0.000 -16.025  ;
    ORIGIN 0.000 16.025 ;
    SIZE 25.000 BY 95.500 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  25.000 -16.025 33.750 73.975 ;
        RECT  0.000 -16.025 25.000 79.475 ;
        RECT  -8.750 -16.025 0.000 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
        LAYER M9 ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  25.000 -16.025 33.750 73.975 ;
        RECT  0.000 -16.025 25.000 79.475 ;
        RECT  -8.750 -16.025 0.000 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
        LAYER AP ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  -8.750 -16.025 33.750 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
    END
END PAD50GAU_DS_SL

MACRO PAD50GU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD50GU_DS_SL 0.000 -16.025  ;
    ORIGIN 0.000 16.025 ;
    SIZE 25.000 BY 95.500 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  25.000 -16.025 33.750 73.975 ;
        RECT  0.000 -16.025 25.000 79.475 ;
        RECT  -8.750 -16.025 0.000 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
        LAYER M9 ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  25.000 -16.025 33.750 73.975 ;
        RECT  0.000 -16.025 25.000 79.475 ;
        RECT  -8.750 -16.025 0.000 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
        LAYER AP ;
        POLYGON  35.500 72.225 33.750 73.975 33.750 -16.025 35.500 -14.275 ;
        RECT  -8.750 -16.025 33.750 73.975 ;
        POLYGON  -8.750 73.975 -10.500 72.225 -10.500 -14.275 -8.750 -16.025 ;
    END
END PAD50GU_DS_SL

MACRO PAD50NAU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD50NAU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 183.975 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  25.000 93.975 33.750 183.975 ;
        RECT  0.000 0.000 25.000 183.975 ;
        RECT  -8.750 93.975 0.000 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
        LAYER M9 ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  25.000 93.975 33.750 183.975 ;
        RECT  0.000 0.000 25.000 183.975 ;
        RECT  -8.750 93.975 0.000 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
        LAYER AP ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  -8.750 93.975 33.750 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
    END
END PAD50NAU_DS_SL

MACRO PAD50NU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD50NU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 183.975 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  25.000 93.975 33.750 183.975 ;
        RECT  0.000 0.000 25.000 183.975 ;
        RECT  -8.750 93.975 0.000 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
        LAYER M9 ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  25.000 93.975 33.750 183.975 ;
        RECT  0.000 0.000 25.000 183.975 ;
        RECT  -8.750 93.975 0.000 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
        LAYER AP ;
        POLYGON  35.500 182.225 33.750 183.975 33.750 93.975 35.500 95.725 ;
        RECT  -8.750 93.975 33.750 183.975 ;
        POLYGON  -8.750 183.975 -10.500 182.225 -10.500 95.725 -8.750 93.975 ;
    END
END PAD50NU_DS_SL

MACRO PAD60GAU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD60GAU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 79.475 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  25.000 5.255 38.750 73.255 ;
        RECT  0.000 0.000 25.000 79.475 ;
        RECT  -13.750 5.255 0.000 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
        LAYER M9 ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  25.000 5.255 38.750 73.255 ;
        RECT  0.000 0.000 25.000 79.475 ;
        RECT  -13.750 5.255 0.000 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
        LAYER AP ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  -13.750 5.255 38.750 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
    END
END PAD60GAU_DS_SL

MACRO PAD60GU_DS
    CLASS BLOCK ;
    FOREIGN PAD60GU_DS 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 86.755 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  43.000 71.505 41.250 73.255 41.250 5.255 43.000 7.005 ;
        RECT  30.000 5.255 41.250 73.255 ;
        RECT  0.000 0.000 30.000 86.755 ;
        RECT  -11.250 5.255 0.000 73.255 ;
        POLYGON  -11.250 73.255 -13.000 71.505 -13.000 7.005 -11.250 5.255 ;
        LAYER M9 ;
        POLYGON  43.000 71.505 41.250 73.255 41.250 5.255 43.000 7.005 ;
        RECT  30.000 5.255 41.250 73.255 ;
        RECT  0.000 0.000 30.000 86.755 ;
        RECT  -11.250 5.255 0.000 73.255 ;
        POLYGON  -11.250 73.255 -13.000 71.505 -13.000 7.005 -11.250 5.255 ;
        LAYER AP ;
        POLYGON  43.000 71.505 41.250 73.255 41.250 5.255 43.000 7.005 ;
        RECT  -11.250 5.255 41.250 73.255 ;
        POLYGON  -11.250 73.255 -13.000 71.505 -13.000 7.005 -11.250 5.255 ;
    END
END PAD60GU_DS

MACRO PAD60GU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD60GU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 79.475 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  25.000 5.255 38.750 73.255 ;
        RECT  0.000 0.000 25.000 79.475 ;
        RECT  -13.750 5.255 0.000 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
        LAYER M9 ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  25.000 5.255 38.750 73.255 ;
        RECT  0.000 0.000 25.000 79.475 ;
        RECT  -13.750 5.255 0.000 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
        LAYER AP ;
        POLYGON  40.500 71.505 38.750 73.255 38.750 5.255 40.500 7.005 ;
        RECT  -13.750 5.255 38.750 73.255 ;
        POLYGON  -13.750 73.255 -15.500 71.505 -15.500 7.005 -13.750 5.255 ;
    END
END PAD60GU_DS_SL

MACRO PAD60NAU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD60NAU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 169.255 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  25.000 101.255 38.750 169.255 ;
        RECT  0.000 0.000 25.000 169.255 ;
        RECT  -13.750 101.255 0.000 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
        LAYER M9 ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  25.000 101.255 38.750 169.255 ;
        RECT  0.000 0.000 25.000 169.255 ;
        RECT  -13.750 101.255 0.000 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
        LAYER AP ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  -13.750 101.255 38.750 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
    END
END PAD60NAU_DS_SL

MACRO PAD60NU_DS
    CLASS BLOCK ;
    FOREIGN PAD60NU_DS 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 169.255 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  43.000 167.505 41.250 169.255 41.250 101.255 43.000 103.005 ;
        RECT  30.000 101.255 41.250 169.255 ;
        RECT  0.000 0.000 30.000 169.255 ;
        RECT  -11.250 101.255 0.000 169.255 ;
        POLYGON  -11.250 169.255 -13.000 167.505 -13.000 103.005 -11.250 101.255 ;
        LAYER M9 ;
        POLYGON  43.000 167.505 41.250 169.255 41.250 101.255 43.000 103.005 ;
        RECT  30.000 101.255 41.250 169.255 ;
        RECT  0.000 0.000 30.000 169.255 ;
        RECT  -11.250 101.255 0.000 169.255 ;
        POLYGON  -11.250 169.255 -13.000 167.505 -13.000 103.005 -11.250 101.255 ;
        LAYER AP ;
        POLYGON  43.000 167.505 41.250 169.255 41.250 101.255 43.000 103.005 ;
        RECT  -11.250 101.255 41.250 169.255 ;
        POLYGON  -11.250 169.255 -13.000 167.505 -13.000 103.005 -11.250 101.255 ;
    END
END PAD60NU_DS

MACRO PAD60NU_DS_SL
    CLASS BLOCK ;
    FOREIGN PAD60NU_DS_SL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.000 BY 169.255 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  25.000 101.255 38.750 169.255 ;
        RECT  0.000 0.000 25.000 169.255 ;
        RECT  -13.750 101.255 0.000 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
        LAYER M9 ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  25.000 101.255 38.750 169.255 ;
        RECT  0.000 0.000 25.000 169.255 ;
        RECT  -13.750 101.255 0.000 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
        LAYER AP ;
        POLYGON  40.500 167.505 38.750 169.255 38.750 101.255 40.500 103.005 ;
        RECT  -13.750 101.255 38.750 169.255 ;
        POLYGON  -13.750 169.255 -15.500 167.505 -15.500 103.005 -13.750 101.255 ;
    END
END PAD60NU_DS_SL

MACRO PAD70GU_DS
    CLASS BLOCK ;
    FOREIGN PAD70GU_DS 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 86.755 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  45.000 71.505 43.250 73.255 43.250 5.255 45.000 7.005 ;
        RECT  30.000 5.255 43.250 73.255 ;
        RECT  0.000 0.000 30.000 86.755 ;
        RECT  -13.250 5.255 0.000 73.255 ;
        POLYGON  -13.250 73.255 -15.000 71.505 -15.000 7.005 -13.250 5.255 ;
        LAYER M9 ;
        POLYGON  45.000 71.505 43.250 73.255 43.250 5.255 45.000 7.005 ;
        RECT  30.000 5.255 43.250 73.255 ;
        RECT  0.000 0.000 30.000 86.755 ;
        RECT  -13.250 5.255 0.000 73.255 ;
        POLYGON  -13.250 73.255 -15.000 71.505 -15.000 7.005 -13.250 5.255 ;
        LAYER AP ;
        POLYGON  45.000 71.505 43.250 73.255 43.250 5.255 45.000 7.005 ;
        RECT  -13.250 5.255 43.250 73.255 ;
        POLYGON  -13.250 73.255 -15.000 71.505 -15.000 7.005 -13.250 5.255 ;
    END
END PAD70GU_DS

MACRO PAD70NU_DS
    CLASS BLOCK ;
    FOREIGN PAD70NU_DS 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 175.255 ;
    SYMMETRY X Y R90 ;
    OBS
        LAYER M8 ;
        POLYGON  45.000 173.505 43.250 175.255 43.250 107.255 45.000 109.005 ;
        RECT  30.000 107.255 43.250 175.255 ;
        RECT  0.000 0.000 30.000 175.255 ;
        RECT  -13.250 107.255 0.000 175.255 ;
        POLYGON  -13.250 175.255 -15.000 173.505 -15.000 109.005 -13.250 107.255 ;
        LAYER M9 ;
        POLYGON  45.000 173.505 43.250 175.255 43.250 107.255 45.000 109.005 ;
        RECT  30.000 107.255 43.250 175.255 ;
        RECT  0.000 0.000 30.000 175.255 ;
        RECT  -13.250 107.255 0.000 175.255 ;
        POLYGON  -13.250 175.255 -15.000 173.505 -15.000 109.005 -13.250 107.255 ;
        LAYER AP ;
        POLYGON  45.000 173.505 43.250 175.255 43.250 107.255 45.000 109.005 ;
        RECT  -13.250 107.255 43.250 175.255 ;
        POLYGON  -13.250 175.255 -15.000 173.505 -15.000 109.005 -13.250 107.255 ;
    END
END PAD70NU_DS

END LIBRARY
