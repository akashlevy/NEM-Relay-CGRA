VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MANUFACTURINGGRID 0.005 ;

MACRO nem_ohmux_invd1_2i_8b
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN nem_ohmux_invd1_2i_8b 0 0 ;
  SIZE 8.84 BY 4.38 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN I0_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.295 2.87 2.465 3.04 ;
    END
  END I0_0
  PIN I0_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.895 2.515 2.065 2.685 ;
    END
  END I0_7
  PIN I0_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.045 2.56 3.215 2.73 ;
    END
  END I0_1
  PIN I0_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 3.195 2.23 3.365 2.4 ;
    END
  END I0_2
  PIN I0_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.95 1.535 3.12 1.705 ;
    END
  END I0_3
  PIN I0_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.575 1.385 2.745 1.555 ;
    END
  END I0_4
  PIN I0_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.84 1.655 2.01 1.825 ;
    END
  END I0_5
  PIN I0_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 1.685 1.995 1.855 2.165 ;
    END
  END I0_6
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 2.365 2.095 2.535 2.265 ;
    END
  END S0
  PIN ZN_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.18 1.265 3.325 1.345 ;
        RECT 3.255 0.515 3.325 1.345 ;
        RECT 3.18 0.515 3.325 0.595 ;
    END
  END ZN_3
  PIN ZN_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.76 1.265 2.905 1.345 ;
        RECT 2.835 0.515 2.905 1.345 ;
        RECT 2.76 0.515 2.905 0.595 ;
    END
  END ZN_6
  PIN ZN_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 1.265 2.485 1.345 ;
        RECT 2.415 0.515 2.485 1.345 ;
        RECT 2.34 0.515 2.485 0.595 ;
    END
  END ZN_4
  PIN ZN_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.92 1.265 2.065 1.345 ;
        RECT 1.995 0.515 2.065 1.345 ;
        RECT 1.92 0.515 2.065 0.595 ;
    END
  END ZN_5
  PIN ZN_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.18 3.785 3.325 3.865 ;
        RECT 3.255 3.035 3.325 3.865 ;
        RECT 3.18 3.035 3.325 3.115 ;
    END
  END ZN_1
  PIN ZN_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.76 3.785 2.905 3.865 ;
        RECT 2.835 3.035 2.905 3.865 ;
        RECT 2.76 3.035 2.905 3.115 ;
    END
  END ZN_2
  PIN ZN_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 3.785 2.485 3.865 ;
        RECT 2.415 3.035 2.485 3.865 ;
        RECT 2.34 3.035 2.485 3.115 ;
    END
  END ZN_0
  PIN ZN_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.92 3.785 2.065 3.865 ;
        RECT 1.995 3.035 2.065 3.865 ;
        RECT 1.92 3.035 2.065 3.115 ;
    END
  END ZN_7
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.145 2.095 6.315 2.265 ;
    END
  END S1
  PIN I1_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.975 2.23 7.145 2.4 ;
    END
  END I1_2
  PIN I1_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.355 1.38 6.525 1.55 ;
    END
  END I1_4
  PIN I1_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.73 1.535 6.9 1.705 ;
    END
  END I1_3
  PIN I1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.825 2.56 6.995 2.73 ;
    END
  END I1_1
  PIN I1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 6.12 2.87 6.29 3.04 ;
    END
  END I1_0
  PIN I1_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.62 1.655 5.79 1.825 ;
    END
  END I1_5
  PIN I1_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.73 2.71 5.9 2.88 ;
    END
  END I1_7
  PIN I1_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 5.465 1.995 5.635 2.165 ;
    END
  END I1_6
  PIN VSNEM
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M8 ;
        RECT 0 0 1.28 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 3.78 0 5.06 4.38 ;
    END
    PORT
      LAYER M8 ;
        RECT 7.56 0 8.84 4.38 ;
    END
  END VSNEM
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.68 2.705 3.36 2.935 ;
        RECT 3.02 2.705 3.1 3.145 ;
        RECT 2.6 2.705 2.68 3.145 ;
        RECT 2.18 2.705 2.26 3.145 ;
        RECT 1.76 2.705 1.84 3.145 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.68 0.185 3.36 0.415 ;
        RECT 3.02 0.185 3.1 0.625 ;
        RECT 2.6 0.185 2.68 0.625 ;
        RECT 2.18 0.185 2.26 0.625 ;
        RECT 1.76 0.185 1.84 0.625 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.68 3.965 3.36 4.195 ;
        RECT 3.02 3.755 3.1 4.195 ;
        RECT 2.6 3.755 2.68 4.195 ;
        RECT 2.18 3.755 2.26 4.195 ;
        RECT 1.76 3.755 1.84 4.195 ;
    END
    PORT
      LAYER M1 ;
        RECT 1.68 1.445 3.36 1.675 ;
        RECT 3.02 1.235 3.1 1.675 ;
        RECT 2.6 1.235 2.68 1.675 ;
        RECT 2.18 1.235 2.26 1.675 ;
        RECT 1.76 1.235 1.84 1.675 ;
    END
  END VDD
  OBS
    LAYER OVERLAP ;
      RECT 0 0 8.84 4.38 ;
    LAYER M1 ;
      RECT 2.975 0.795 3.045 1.065 ;
      RECT 2.975 0.845 3.18 0.915 ;
      RECT 2.975 3.315 3.045 3.585 ;
      RECT 2.975 3.365 3.18 3.435 ;
      RECT 2.555 0.795 2.625 1.065 ;
      RECT 2.555 0.845 2.76 0.915 ;
      RECT 2.555 3.315 2.625 3.585 ;
      RECT 2.555 3.365 2.76 3.435 ;
      RECT 2.135 0.795 2.205 1.065 ;
      RECT 2.135 0.845 2.34 0.915 ;
      RECT 2.135 3.315 2.205 3.585 ;
      RECT 2.135 3.365 2.34 3.435 ;
      RECT 1.715 0.795 1.785 1.065 ;
      RECT 1.715 0.845 1.92 0.915 ;
      RECT 1.715 3.315 1.785 3.585 ;
      RECT 1.715 3.365 1.92 3.435 ;
    LAYER M2 ;
      RECT 2.975 0.675 3.045 1.065 ;
      RECT 2.975 3.195 3.045 3.585 ;
      RECT 2.555 0.675 2.625 1.065 ;
      RECT 2.555 3.195 2.625 3.585 ;
      RECT 2.135 0.675 2.205 1.065 ;
      RECT 2.135 3.195 2.205 3.585 ;
      RECT 1.715 0.675 1.785 1.065 ;
      RECT 1.715 3.195 1.785 3.585 ;
    LAYER M3 ;
      RECT 2.975 0.675 3.045 1.065 ;
      RECT 2.975 3.195 3.045 3.585 ;
      RECT 2.555 0.675 2.625 1.065 ;
      RECT 2.555 3.195 2.625 3.585 ;
      RECT 2.135 0.675 2.205 1.065 ;
      RECT 2.135 3.195 2.205 3.585 ;
      RECT 1.715 0.675 1.785 1.065 ;
      RECT 1.715 3.195 1.785 3.585 ;
    LAYER M4 ;
      RECT 2.975 0.675 3.045 1.065 ;
      RECT 2.975 3.195 3.045 3.585 ;
      RECT 2.555 0.675 2.625 1.065 ;
      RECT 2.555 3.195 2.625 3.585 ;
      RECT 2.135 0.675 2.205 1.065 ;
      RECT 2.135 3.195 2.205 3.585 ;
      RECT 1.715 0.675 1.785 1.065 ;
      RECT 1.715 3.195 1.785 3.585 ;
    LAYER M5 ;
      RECT 2.975 0.675 3.045 1.065 ;
      RECT 2.975 3.195 3.045 3.585 ;
      RECT 2.555 0.675 2.625 1.065 ;
      RECT 2.555 3.195 2.625 3.585 ;
      RECT 2.135 0.675 2.205 1.065 ;
      RECT 2.135 3.195 2.205 3.585 ;
      RECT 1.715 0.675 1.785 1.065 ;
      RECT 1.715 3.195 1.785 3.585 ;
    LAYER M6 ;
      RECT 2.975 0.795 3.045 1.475 ;
      RECT 2.975 2.87 3.045 3.585 ;
      RECT 2.555 0.795 2.625 1.325 ;
      RECT 2.555 2.87 2.625 3.585 ;
      RECT 2.135 0.795 2.205 1.585 ;
      RECT 2.135 2.87 2.205 3.585 ;
      RECT 1.715 0.795 1.785 1.585 ;
      RECT 1.715 2.87 1.785 3.585 ;
    LAYER M7 ;
      RECT 2.945 1.215 3.08 1.455 ;
      RECT 2.97 2.8 3.05 3.14 ;
      RECT 2.455 1.21 2.72 1.315 ;
      RECT 2.555 2.75 2.625 3.14 ;
      RECT 2.13 1.245 2.21 1.585 ;
      RECT 2.135 2.75 2.205 3.14 ;
      RECT 1.71 1.245 1.79 1.585 ;
      RECT 1.715 2.75 1.785 3.14 ;
    LAYER M8 ;
      RECT 7.205 3.335 7.335 3.465 ;
      RECT 7.235 2.15 7.305 3.465 ;
      RECT 7.205 2.15 7.335 2.28 ;
      RECT 7.02 1.37 7.15 1.5 ;
      RECT 7.05 0.505 7.12 1.5 ;
      RECT 7.02 0.505 7.15 0.635 ;
      RECT 6.995 3.735 7.125 3.865 ;
      RECT 7.025 2.885 7.095 3.865 ;
      RECT 6.995 2.885 7.125 3.015 ;
      RECT 5.52 3.535 5.65 3.665 ;
      RECT 5.55 2.87 5.62 3.665 ;
      RECT 5.48 2.87 5.62 3 ;
      RECT 5.49 1.38 5.62 1.51 ;
      RECT 5.52 0.705 5.59 1.51 ;
      RECT 5.49 0.705 5.62 0.835 ;
      RECT 5.275 2.11 5.405 2.24 ;
      RECT 5.305 0.905 5.375 2.24 ;
      RECT 5.275 0.905 5.405 1.035 ;
      RECT 3.425 3.335 3.555 3.465 ;
      RECT 3.455 2.15 3.525 3.465 ;
      RECT 3.425 2.15 3.555 2.28 ;
      RECT 3.24 1.37 3.37 1.5 ;
      RECT 3.27 0.505 3.34 1.5 ;
      RECT 3.24 0.505 3.37 0.635 ;
      RECT 3.215 3.735 3.345 3.865 ;
      RECT 3.245 2.885 3.315 3.865 ;
      RECT 3.215 2.885 3.345 3.015 ;
      RECT 2.975 0.505 3.045 1.465 ;
      RECT 2.945 0.505 3.075 0.635 ;
      RECT 2.945 3.735 3.075 3.865 ;
      RECT 2.975 2.87 3.045 3.865 ;
      RECT 2.555 0.905 2.625 1.315 ;
      RECT 2.525 0.905 2.655 1.035 ;
      RECT 2.525 3.335 2.655 3.465 ;
      RECT 2.555 2.87 2.625 3.465 ;
      RECT 2.135 1.105 2.205 1.515 ;
      RECT 2.105 1.105 2.235 1.235 ;
      RECT 2.105 3.135 2.235 3.265 ;
      RECT 2.135 2.87 2.205 3.265 ;
      RECT 1.685 3.535 1.815 3.665 ;
      RECT 1.715 2.87 1.785 3.665 ;
      RECT 1.715 2.87 1.845 3 ;
      RECT 1.69 1.38 1.82 1.51 ;
      RECT 1.715 0.705 1.785 1.51 ;
      RECT 1.685 0.705 1.815 0.835 ;
      RECT 1.495 2.11 1.625 2.24 ;
      RECT 1.525 0.905 1.595 2.24 ;
      RECT 1.495 0.905 1.625 1.035 ;
      RECT 6.965 2.225 7.135 2.395 ;
      RECT 6.825 2.565 6.995 2.735 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 6.12 2.87 6.29 3.04 ;
      RECT 5.73 2.71 5.9 2.88 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 3.185 2.225 3.355 2.395 ;
      RECT 3.045 2.565 3.215 2.735 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 2.295 2.87 2.465 3.04 ;
      RECT 1.965 2.535 2.09 2.79 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.695 1.99 1.865 2.16 ;
    LAYER M9 ;
      RECT 2.34 2.87 2.51 3.04 ;
      RECT 2.335 2.87 2.51 3 ;
      RECT 8.05 0.165 8.35 0.435 ;
      RECT 8.05 3.945 8.35 4.215 ;
      RECT 7.205 2.15 7.44 2.28 ;
      RECT 1.495 0.505 7.335 0.635 ;
      RECT 1.495 0.705 7.335 0.835 ;
      RECT 1.495 0.905 7.335 1.035 ;
      RECT 1.495 1.105 7.335 1.235 ;
      RECT 1.495 3.135 7.335 3.265 ;
      RECT 1.495 3.335 7.335 3.465 ;
      RECT 1.495 3.535 7.335 3.665 ;
      RECT 1.495 3.735 7.335 3.865 ;
      RECT 7 1.35 7.17 1.52 ;
      RECT 6.975 2.865 7.145 3.035 ;
      RECT 6.965 2.225 7.135 2.395 ;
      RECT 6.825 2.565 6.995 2.735 ;
      RECT 6.73 1.535 6.9 1.705 ;
      RECT 6.34 1.385 6.51 1.555 ;
      RECT 6.145 2.09 6.315 2.26 ;
      RECT 6.12 2.87 6.29 3.04 ;
      RECT 5.73 2.71 5.9 2.88 ;
      RECT 5.62 1.635 5.79 1.805 ;
      RECT 5.475 1.99 5.645 2.16 ;
      RECT 5.47 1.36 5.64 1.53 ;
      RECT 5.46 2.85 5.63 3.02 ;
      RECT 5.19 2.11 5.405 2.24 ;
      RECT 4.27 0.165 4.57 0.435 ;
      RECT 4.27 3.945 4.57 4.215 ;
      RECT 3.425 2.15 3.66 2.28 ;
      RECT 3.22 1.35 3.39 1.52 ;
      RECT 3.195 2.865 3.365 3.035 ;
      RECT 3.185 2.225 3.355 2.395 ;
      RECT 3.045 2.565 3.215 2.735 ;
      RECT 2.95 1.535 3.12 1.705 ;
      RECT 2.56 1.385 2.73 1.555 ;
      RECT 2.365 2.09 2.535 2.26 ;
      RECT 1.955 2.69 2.125 2.86 ;
      RECT 1.84 1.635 2.01 1.805 ;
      RECT 1.695 1.99 1.865 2.16 ;
      RECT 1.695 2.85 1.865 3.02 ;
      RECT 1.67 1.36 1.84 1.53 ;
      RECT 1.41 2.11 1.625 2.24 ;
      RECT 0.49 0.165 0.79 0.435 ;
      RECT 0.49 3.945 0.79 4.215 ;
    LAYER M10 ;
      RECT 4.92 3.375 7.7 3.58 ;
      RECT 7.49 0.8 7.7 3.58 ;
      RECT 6.41 3.075 7.7 3.58 ;
      RECT 7.19 2.335 7.7 3.58 ;
      RECT 4.92 3.07 6.16 3.58 ;
      RECT 4.92 3.07 6.165 3.22 ;
      RECT 6.315 1.57 6.67 3.125 ;
      RECT 4.92 3.07 6.94 3.125 ;
      RECT 6.41 2.785 6.94 3.58 ;
      RECT 4.92 3.065 6.065 3.58 ;
      RECT 5.965 0.8 6.065 3.58 ;
      RECT 5.68 2.91 6.065 3.58 ;
      RECT 4.92 2.295 5.43 3.58 ;
      RECT 5.68 1.845 5.715 3.58 ;
      RECT 6.315 2.785 7.7 2.825 ;
      RECT 7.185 1.555 7.24 2.825 ;
      RECT 5.965 1.26 6.315 2.82 ;
      RECT 4.92 2.295 5.715 2.815 ;
      RECT 7.03 2.435 7.7 2.825 ;
      RECT 5.965 1.715 6.78 2.82 ;
      RECT 4.92 2.295 6.78 2.66 ;
      RECT 5.83 0.8 6.215 2.66 ;
      RECT 4.92 2.435 7.7 2.535 ;
      RECT 5.375 2.2 6.935 2.535 ;
      RECT 5.83 1.715 6.935 2.535 ;
      RECT 4.92 0.8 5.125 3.58 ;
      RECT 5.675 1.845 6.935 2.535 ;
      RECT 5.375 1.565 5.425 3.58 ;
      RECT 6.92 1.555 7.24 2.185 ;
      RECT 7.2 0.8 7.7 2.085 ;
      RECT 4.92 0.8 5.42 2.045 ;
      RECT 4.92 1.845 7.7 1.95 ;
      RECT 4.92 1.565 5.58 1.95 ;
      RECT 5.67 0.8 6.215 1.595 ;
      RECT 6.565 0.8 6.67 3.58 ;
      RECT 4.92 1.565 6.315 1.595 ;
      RECT 6.92 0.8 6.95 2.185 ;
      RECT 6.565 0.8 6.95 1.465 ;
      RECT 5.67 1.26 6.95 1.32 ;
      RECT 4.92 0.8 6.215 1.315 ;
      RECT 6.465 0.8 7.7 1.305 ;
      RECT 6.455 1.16 7.7 1.305 ;
      RECT 4.92 0.8 7.7 1.01 ;
      RECT 1.14 3.375 3.92 3.58 ;
      RECT 3.71 0.8 3.92 3.58 ;
      RECT 2.63 3.075 3.92 3.58 ;
      RECT 3.41 2.335 3.92 3.58 ;
      RECT 1.14 3.07 2.38 3.58 ;
      RECT 1.14 3.07 2.385 3.22 ;
      RECT 2.535 1.57 2.89 3.125 ;
      RECT 1.14 3.07 3.16 3.125 ;
      RECT 2.63 2.785 3.16 3.58 ;
      RECT 1.14 3.065 2.285 3.58 ;
      RECT 2.185 0.8 2.285 3.58 ;
      RECT 1.9 2.91 2.285 3.58 ;
      RECT 1.14 2.295 1.65 3.58 ;
      RECT 1.9 1.845 1.935 3.58 ;
      RECT 2.535 2.785 3.92 2.825 ;
      RECT 3.405 1.555 3.46 2.825 ;
      RECT 2.185 1.26 2.535 2.82 ;
      RECT 1.14 2.295 1.935 2.815 ;
      RECT 3.25 2.435 3.92 2.825 ;
      RECT 2.185 1.715 3 2.82 ;
      RECT 1.14 2.295 3 2.66 ;
      RECT 2.05 0.8 2.435 2.66 ;
      RECT 1.14 2.435 3.92 2.535 ;
      RECT 1.595 2.2 3.155 2.535 ;
      RECT 2.05 1.715 3.155 2.535 ;
      RECT 1.14 0.8 1.345 3.58 ;
      RECT 1.895 1.845 3.155 2.535 ;
      RECT 1.595 1.565 1.645 3.58 ;
      RECT 3.14 1.555 3.46 2.185 ;
      RECT 3.42 0.8 3.92 2.085 ;
      RECT 1.14 0.8 1.64 2.045 ;
      RECT 1.14 1.845 3.92 1.95 ;
      RECT 1.14 1.565 1.8 1.95 ;
      RECT 1.89 0.8 2.435 1.595 ;
      RECT 2.785 0.8 2.89 3.58 ;
      RECT 1.14 1.565 2.535 1.595 ;
      RECT 3.14 0.8 3.17 2.185 ;
      RECT 2.785 0.8 3.17 1.465 ;
      RECT 1.89 1.26 3.17 1.32 ;
      RECT 1.14 0.8 2.435 1.315 ;
      RECT 2.685 0.8 3.92 1.305 ;
      RECT 2.675 1.16 3.92 1.305 ;
      RECT 1.14 0.8 3.92 1.01 ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 7.29 2.135 7.44 2.285 ;
      RECT 7 1.354 7.15 1.504 ;
      RECT 6.991 2.873 7.141 3.023 ;
      RECT 6.985 2.236 7.135 2.386 ;
      RECT 6.832 2.584 6.982 2.734 ;
      RECT 6.718 1.517 6.868 1.667 ;
      RECT 6.366 1.368 6.516 1.518 ;
      RECT 6.264 1.061 6.414 1.211 ;
      RECT 6.211 3.173 6.361 3.323 ;
      RECT 6.115 2.87 6.265 3.02 ;
      RECT 5.764 2.708 5.914 2.858 ;
      RECT 5.63 1.643 5.78 1.793 ;
      RECT 5.478 2.866 5.628 3.016 ;
      RECT 5.477 1.998 5.627 2.148 ;
      RECT 5.47 1.363 5.62 1.513 ;
      RECT 5.173 2.096 5.323 2.246 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 3.51 2.135 3.66 2.285 ;
      RECT 3.22 1.354 3.37 1.504 ;
      RECT 3.211 2.873 3.361 3.023 ;
      RECT 3.205 2.236 3.355 2.386 ;
      RECT 3.052 2.584 3.202 2.734 ;
      RECT 2.938 1.517 3.088 1.667 ;
      RECT 2.586 1.368 2.736 1.518 ;
      RECT 2.484 1.061 2.634 1.211 ;
      RECT 2.431 3.173 2.581 3.323 ;
      RECT 2.335 2.87 2.485 3.02 ;
      RECT 1.984 2.708 2.134 2.858 ;
      RECT 1.85 1.643 2 1.793 ;
      RECT 1.698 2.866 1.848 3.016 ;
      RECT 1.697 1.998 1.847 2.148 ;
      RECT 1.69 1.363 1.84 1.513 ;
      RECT 1.393 2.096 1.543 2.246 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
    LAYER NEMANC ;
      RECT 8 0.1 8.4 0.5 ;
      RECT 8 3.88 8.4 4.28 ;
      RECT 4.22 0.1 4.62 0.5 ;
      RECT 4.22 3.88 4.62 4.28 ;
      RECT 0.44 0.1 0.84 0.5 ;
      RECT 0.44 3.88 0.84 4.28 ;
    LAYER NEMCHAN ;
      RECT 7.075 2.22 7.155 2.37 ;
      RECT 7.075 2.22 7.195 2.355 ;
      RECT 7.075 2.22 7.235 2.34 ;
      RECT 7.075 2.22 7.275 2.325 ;
      RECT 7.315 2.14 7.34 2.305 ;
      RECT 7.035 2.23 7.34 2.3 ;
      RECT 7.155 2.195 7.38 2.29 ;
      RECT 7.035 2.26 7.39 2.285 ;
      RECT 7.115 2.205 7.38 2.29 ;
      RECT 7.195 2.18 7.34 2.305 ;
      RECT 7.275 2.155 7.315 2.315 ;
      RECT 7.235 2.165 7.34 2.305 ;
      RECT 7 2.705 7.04 2.975 ;
      RECT 6.96 2.78 7.08 2.95 ;
      RECT 6.96 2.855 7.12 2.93 ;
      RECT 6.96 2.895 7.13 2.915 ;
      RECT 6.92 2.645 6.96 2.88 ;
      RECT 6.88 2.665 7 2.805 ;
      RECT 6.84 2.685 7 2.735 ;
      RECT 6.92 2.65 7 2.88 ;
      RECT 6.835 1.465 6.875 1.64 ;
      RECT 6.795 1.49 6.875 1.625 ;
      RECT 6.795 1.49 6.915 1.62 ;
      RECT 6.795 1.49 6.955 1.595 ;
      RECT 6.755 1.51 6.995 1.565 ;
      RECT 6.995 1.375 7.035 1.55 ;
      RECT 6.995 1.395 7.075 1.525 ;
      RECT 6.835 1.465 7.11 1.51 ;
      RECT 6.875 1.445 7.075 1.525 ;
      RECT 6.955 1.4 6.995 1.57 ;
      RECT 6.915 1.42 7.075 1.525 ;
      RECT 6.39 1.115 6.41 1.46 ;
      RECT 6.39 1.175 6.45 1.445 ;
      RECT 6.35 1.295 6.49 1.435 ;
      RECT 6.35 1.39 6.51 1.425 ;
      RECT 6.31 1.14 6.41 1.345 ;
      RECT 6.27 1.15 6.41 1.22 ;
      RECT 6.35 1.125 6.41 1.435 ;
      RECT 6.24 2.92 6.26 3.26 ;
      RECT 6.24 2.98 6.3 3.25 ;
      RECT 6.2 3.1 6.34 3.24 ;
      RECT 6.2 3.195 6.36 3.23 ;
      RECT 6.16 2.945 6.26 3.16 ;
      RECT 6.12 2.955 6.26 3.035 ;
      RECT 6.2 2.93 6.26 3.24 ;
      RECT 5.595 2.82 5.635 2.99 ;
      RECT 5.555 2.84 5.635 2.975 ;
      RECT 5.555 2.84 5.675 2.97 ;
      RECT 5.555 2.84 5.755 2.93 ;
      RECT 5.515 2.865 5.755 2.915 ;
      RECT 5.515 2.865 5.795 2.905 ;
      RECT 5.795 2.72 5.805 2.895 ;
      RECT 5.715 2.755 5.845 2.88 ;
      RECT 5.595 2.82 5.875 2.86 ;
      RECT 5.635 2.8 5.845 2.88 ;
      RECT 5.675 2.78 5.715 2.95 ;
      RECT 5.755 2.735 5.805 2.895 ;
      RECT 5.64 1.48 5.68 1.745 ;
      RECT 5.6 1.555 5.72 1.72 ;
      RECT 5.6 1.625 5.76 1.7 ;
      RECT 5.6 1.665 5.77 1.685 ;
      RECT 5.56 1.415 5.6 1.65 ;
      RECT 5.52 1.44 5.64 1.58 ;
      RECT 5.48 1.46 5.64 1.51 ;
      RECT 5.56 1.425 5.64 1.65 ;
      RECT 5.265 2.08 5.305 2.23 ;
      RECT 5.265 2.08 5.345 2.225 ;
      RECT 5.265 2.08 5.385 2.21 ;
      RECT 5.265 2.08 5.425 2.2 ;
      RECT 5.505 2 5.53 2.17 ;
      RECT 5.225 2.09 5.53 2.165 ;
      RECT 5.345 2.06 5.57 2.155 ;
      RECT 5.225 2.135 5.575 2.145 ;
      RECT 5.305 2.065 5.57 2.155 ;
      RECT 5.345 2.055 5.53 2.17 ;
      RECT 5.465 2.015 5.505 2.175 ;
      RECT 5.385 2.04 5.53 2.17 ;
      RECT 5.425 2.025 5.465 2.185 ;
      RECT 3.295 2.22 3.375 2.37 ;
      RECT 3.295 2.22 3.415 2.355 ;
      RECT 3.295 2.22 3.455 2.34 ;
      RECT 3.295 2.22 3.495 2.325 ;
      RECT 3.535 2.14 3.56 2.305 ;
      RECT 3.255 2.23 3.56 2.3 ;
      RECT 3.375 2.195 3.6 2.29 ;
      RECT 3.255 2.26 3.61 2.285 ;
      RECT 3.335 2.205 3.6 2.29 ;
      RECT 3.415 2.18 3.56 2.305 ;
      RECT 3.495 2.155 3.535 2.315 ;
      RECT 3.455 2.165 3.56 2.305 ;
      RECT 3.22 2.705 3.26 2.975 ;
      RECT 3.18 2.78 3.3 2.95 ;
      RECT 3.18 2.855 3.34 2.93 ;
      RECT 3.18 2.895 3.35 2.915 ;
      RECT 3.14 2.645 3.18 2.88 ;
      RECT 3.1 2.665 3.22 2.805 ;
      RECT 3.06 2.685 3.22 2.735 ;
      RECT 3.14 2.65 3.22 2.88 ;
      RECT 3.055 1.465 3.095 1.64 ;
      RECT 3.015 1.49 3.095 1.625 ;
      RECT 3.015 1.49 3.135 1.62 ;
      RECT 3.015 1.49 3.175 1.595 ;
      RECT 2.975 1.51 3.215 1.565 ;
      RECT 3.215 1.375 3.255 1.55 ;
      RECT 3.215 1.395 3.295 1.525 ;
      RECT 3.055 1.465 3.33 1.51 ;
      RECT 3.095 1.445 3.295 1.525 ;
      RECT 3.175 1.4 3.215 1.57 ;
      RECT 3.135 1.42 3.295 1.525 ;
      RECT 2.61 1.115 2.63 1.46 ;
      RECT 2.61 1.175 2.67 1.445 ;
      RECT 2.57 1.295 2.71 1.435 ;
      RECT 2.57 1.39 2.73 1.425 ;
      RECT 2.53 1.14 2.63 1.345 ;
      RECT 2.49 1.15 2.63 1.22 ;
      RECT 2.57 1.125 2.63 1.435 ;
      RECT 2.46 2.92 2.48 3.26 ;
      RECT 2.46 2.98 2.52 3.25 ;
      RECT 2.42 3.1 2.56 3.24 ;
      RECT 2.42 3.195 2.58 3.23 ;
      RECT 2.38 2.945 2.48 3.16 ;
      RECT 2.34 2.955 2.48 3.035 ;
      RECT 2.42 2.93 2.48 3.24 ;
      RECT 1.815 2.82 1.855 2.99 ;
      RECT 1.775 2.84 1.855 2.975 ;
      RECT 1.775 2.84 1.895 2.97 ;
      RECT 1.775 2.84 1.975 2.93 ;
      RECT 1.735 2.865 1.975 2.915 ;
      RECT 1.735 2.865 2.015 2.905 ;
      RECT 2.015 2.72 2.025 2.895 ;
      RECT 1.935 2.755 2.065 2.88 ;
      RECT 1.815 2.82 2.095 2.86 ;
      RECT 1.855 2.8 2.065 2.88 ;
      RECT 1.895 2.78 1.935 2.95 ;
      RECT 1.975 2.735 2.025 2.895 ;
      RECT 1.86 1.48 1.9 1.745 ;
      RECT 1.82 1.555 1.94 1.72 ;
      RECT 1.82 1.625 1.98 1.7 ;
      RECT 1.82 1.665 1.99 1.685 ;
      RECT 1.78 1.415 1.82 1.65 ;
      RECT 1.74 1.44 1.86 1.58 ;
      RECT 1.7 1.46 1.86 1.51 ;
      RECT 1.78 1.425 1.86 1.65 ;
      RECT 1.485 2.08 1.525 2.23 ;
      RECT 1.485 2.08 1.565 2.225 ;
      RECT 1.485 2.08 1.605 2.21 ;
      RECT 1.485 2.08 1.645 2.2 ;
      RECT 1.725 2 1.75 2.17 ;
      RECT 1.445 2.09 1.75 2.165 ;
      RECT 1.565 2.06 1.79 2.155 ;
      RECT 1.445 2.135 1.795 2.145 ;
      RECT 1.525 2.065 1.79 2.155 ;
      RECT 1.565 2.055 1.75 2.17 ;
      RECT 1.685 2.015 1.725 2.175 ;
      RECT 1.605 2.04 1.75 2.17 ;
      RECT 1.645 2.025 1.685 2.185 ;
    LAYER NEMBODY ;
      RECT 7.9 3.78 8.5 4.38 ;
      RECT 4.12 3.78 4.72 4.38 ;
      RECT 4.52 0.8 4.72 4.38 ;
      RECT 0.34 3.78 0.94 4.38 ;
      RECT 0.74 0.8 0.94 4.38 ;
      RECT 4.92 3.78 8.5 3.98 ;
      RECT 1.14 3.78 4.72 3.98 ;
      RECT 4.92 0.8 5.12 3.98 ;
      RECT 1.14 0.8 1.34 3.98 ;
      RECT 4.92 3.38 8.1 3.58 ;
      RECT 7.9 0 8.1 3.58 ;
      RECT 1.14 3.38 4.32 3.58 ;
      RECT 4.12 0 4.32 3.58 ;
      RECT 4.92 0.8 7.7 3.58 ;
      RECT 7.5 0.4 7.7 3.58 ;
      RECT 1.14 0.8 3.92 3.58 ;
      RECT 3.72 0.4 3.92 3.58 ;
      RECT 4.52 0.8 7.7 1 ;
      RECT 0.74 0.8 3.92 1 ;
      RECT 7.9 0 8.5 0.6 ;
      RECT 4.12 0.4 7.7 0.6 ;
      RECT 0.34 0.4 3.92 0.6 ;
      RECT 4.12 0 4.72 0.6 ;
      RECT 0.34 0 0.94 0.6 ;
  END
END nem_ohmux_invd1_2i_8b

END LIBRARY
