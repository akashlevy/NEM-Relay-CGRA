###############################################################################
#TSMC Library/IP Product
#Filename: tcbn40ulpbwp40_c170815.lef
#Technology: CLN40UP
#Product Type: Standard Cell
#Product Name: tcbn40ulpbwp40_c170815
#Version: 130a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################
SITE core
    SIZE 0.140 BY 1.260 ;
    SYMMETRY Y ;
    CLASS CORE ;
END core

SITE gacore
    SIZE 0.700 BY 1.260 ;
    SYMMETRY Y ;
    CLASS CORE ;
END gacore

MACRO AN2D0BWP40
    CLASS CORE ;
    FOREIGN AN2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.050000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.700 0.185 0.735 0.305 ;
        RECT  0.705 0.905 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.490 0.420 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 -0.115 0.840 0.115 ;
        RECT  0.455 -0.115 0.575 0.215 ;
        RECT  0.000 -0.115 0.455 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.150 1.145 0.480 1.375 ;
        RECT  0.070 0.985 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.520 0.655 0.640 ;
        RECT  0.535 0.305 0.605 0.915 ;
        RECT  0.165 0.305 0.535 0.375 ;
        RECT  0.340 0.845 0.535 0.915 ;
        RECT  0.260 0.845 0.340 1.050 ;
        RECT  0.070 0.185 0.165 0.375 ;
    END
END AN2D0BWP40

MACRO AN2D12BWP40
    CLASS CORE ;
    FOREIGN AN2D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.700 3.820 1.025 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.415 0.345 3.745 0.465 ;
        RECT  3.415 0.700 3.740 0.820 ;
        RECT  3.345 0.185 3.415 0.465 ;
        RECT  3.340 0.700 3.415 1.045 ;
        RECT  3.045 0.345 3.345 0.465 ;
        RECT  3.020 0.700 3.340 0.820 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.700 3.020 1.045 ;
        RECT  2.945 0.185 2.975 1.045 ;
        RECT  2.940 0.345 2.945 1.045 ;
        RECT  2.765 0.345 2.940 0.820 ;
        RECT  2.635 0.345 2.765 0.465 ;
        RECT  2.640 0.700 2.765 0.820 ;
        RECT  2.560 0.700 2.640 1.025 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.345 2.565 0.465 ;
        RECT  2.260 0.700 2.560 0.820 ;
        RECT  2.180 0.700 2.260 1.025 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.880 0.345 2.185 0.465 ;
        RECT  1.880 0.700 2.180 0.820 ;
        RECT  1.805 0.185 1.880 0.465 ;
        RECT  1.800 0.700 1.880 1.025 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.495 1.555 0.625 ;
        RECT  1.145 0.495 1.240 0.765 ;
        RECT  0.245 0.695 1.145 0.765 ;
        RECT  0.105 0.525 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.405 0.495 1.000 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.465 ;
        RECT  3.640 -0.115 3.930 0.115 ;
        RECT  3.520 -0.115 3.640 0.265 ;
        RECT  3.240 -0.115 3.520 0.115 ;
        RECT  3.120 -0.115 3.240 0.265 ;
        RECT  2.850 -0.115 3.120 0.115 ;
        RECT  2.730 -0.115 2.850 0.265 ;
        RECT  2.450 -0.115 2.730 0.115 ;
        RECT  2.370 -0.115 2.450 0.275 ;
        RECT  2.070 -0.115 2.370 0.115 ;
        RECT  1.990 -0.115 2.070 0.275 ;
        RECT  1.690 -0.115 1.990 0.115 ;
        RECT  1.610 -0.115 1.690 0.275 ;
        RECT  1.310 -0.115 1.610 0.115 ;
        RECT  1.190 -0.115 1.310 0.125 ;
        RECT  0.125 -0.115 1.190 0.115 ;
        RECT  0.055 -0.115 0.125 0.435 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.670 4.010 1.375 ;
        RECT  3.640 1.145 3.930 1.375 ;
        RECT  3.520 0.890 3.640 1.375 ;
        RECT  3.240 1.145 3.520 1.375 ;
        RECT  3.120 0.890 3.240 1.375 ;
        RECT  2.850 1.145 3.120 1.375 ;
        RECT  2.730 0.890 2.850 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 0.890 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 0.890 2.090 1.375 ;
        RECT  1.690 1.145 1.970 1.375 ;
        RECT  1.610 0.985 1.690 1.375 ;
        RECT  1.270 1.145 1.610 1.375 ;
        RECT  1.190 0.985 1.270 1.375 ;
        RECT  0.890 1.145 1.190 1.375 ;
        RECT  0.810 0.985 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.985 0.510 1.375 ;
        RECT  0.125 1.145 0.430 1.375 ;
        RECT  0.055 0.845 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.740 0.700 3.820 1.025 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.415 0.345 3.745 0.465 ;
        RECT  3.415 0.700 3.740 0.820 ;
        RECT  3.345 0.185 3.415 0.465 ;
        RECT  3.340 0.700 3.415 1.045 ;
        RECT  3.045 0.345 3.345 0.465 ;
        RECT  3.045 0.700 3.340 0.820 ;
        RECT  2.635 0.345 2.695 0.465 ;
        RECT  2.640 0.700 2.695 0.820 ;
        RECT  2.560 0.700 2.640 1.025 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.345 2.565 0.465 ;
        RECT  2.260 0.700 2.560 0.820 ;
        RECT  2.180 0.700 2.260 1.025 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.880 0.345 2.185 0.465 ;
        RECT  1.880 0.700 2.180 0.820 ;
        RECT  1.805 0.185 1.880 0.465 ;
        RECT  1.800 0.700 1.880 1.025 ;
        RECT  1.705 0.545 2.505 0.615 ;
        RECT  1.635 0.345 1.705 0.915 ;
        RECT  0.410 0.345 1.635 0.415 ;
        RECT  1.495 0.845 1.635 0.915 ;
        RECT  0.220 0.205 1.520 0.275 ;
        RECT  1.425 0.845 1.495 1.075 ;
        RECT  1.075 0.845 1.425 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.320 0.845 0.625 0.915 ;
        RECT  0.220 0.845 0.320 1.075 ;
    END
END AN2D12BWP40

MACRO AN2D16BWP40
    CLASS CORE ;
    FOREIGN AN2D16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.275 0.185 5.370 0.465 ;
        RECT  5.280 0.700 5.360 1.025 ;
        RECT  4.980 0.700 5.280 0.820 ;
        RECT  4.985 0.345 5.275 0.465 ;
        RECT  4.900 0.185 4.985 0.465 ;
        RECT  4.900 0.700 4.980 1.025 ;
        RECT  4.600 0.345 4.900 0.465 ;
        RECT  4.600 0.700 4.900 0.820 ;
        RECT  4.525 0.185 4.600 0.465 ;
        RECT  4.520 0.700 4.600 1.025 ;
        RECT  4.215 0.345 4.525 0.465 ;
        RECT  4.215 0.700 4.520 0.820 ;
        RECT  4.145 0.185 4.215 0.465 ;
        RECT  4.140 0.700 4.215 1.045 ;
        RECT  4.095 0.345 4.145 0.465 ;
        RECT  4.095 0.700 4.140 0.820 ;
        RECT  3.885 0.345 4.095 0.820 ;
        RECT  3.820 0.345 3.885 0.465 ;
        RECT  3.820 0.700 3.885 0.820 ;
        RECT  3.745 0.185 3.820 0.465 ;
        RECT  3.740 0.700 3.820 1.025 ;
        RECT  3.435 0.345 3.745 0.465 ;
        RECT  3.440 0.700 3.740 0.820 ;
        RECT  3.360 0.700 3.440 1.025 ;
        RECT  3.365 0.185 3.435 0.465 ;
        RECT  3.055 0.345 3.365 0.465 ;
        RECT  3.060 0.700 3.360 0.820 ;
        RECT  2.980 0.700 3.060 1.025 ;
        RECT  2.985 0.185 3.055 0.465 ;
        RECT  2.680 0.345 2.985 0.465 ;
        RECT  2.680 0.700 2.980 0.820 ;
        RECT  2.605 0.185 2.680 0.465 ;
        RECT  2.600 0.700 2.680 1.025 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.495 2.355 0.625 ;
        RECT  1.435 0.495 1.540 0.765 ;
        RECT  0.245 0.695 1.435 0.765 ;
        RECT  0.105 0.525 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 1.325 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.550 0.465 ;
        RECT  5.190 -0.115 5.470 0.115 ;
        RECT  5.070 -0.115 5.190 0.265 ;
        RECT  4.810 -0.115 5.070 0.115 ;
        RECT  4.690 -0.115 4.810 0.265 ;
        RECT  4.430 -0.115 4.690 0.115 ;
        RECT  4.310 -0.115 4.430 0.265 ;
        RECT  4.040 -0.115 4.310 0.115 ;
        RECT  3.920 -0.115 4.040 0.265 ;
        RECT  3.650 -0.115 3.920 0.115 ;
        RECT  3.530 -0.115 3.650 0.265 ;
        RECT  3.270 -0.115 3.530 0.115 ;
        RECT  3.150 -0.115 3.270 0.265 ;
        RECT  2.890 -0.115 3.150 0.115 ;
        RECT  2.770 -0.115 2.890 0.265 ;
        RECT  2.490 -0.115 2.770 0.115 ;
        RECT  2.410 -0.115 2.490 0.275 ;
        RECT  2.110 -0.115 2.410 0.115 ;
        RECT  1.990 -0.115 2.110 0.125 ;
        RECT  1.690 -0.115 1.990 0.115 ;
        RECT  1.570 -0.115 1.690 0.125 ;
        RECT  0.125 -0.115 1.570 0.115 ;
        RECT  0.055 -0.115 0.125 0.430 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 1.145 5.600 1.375 ;
        RECT  5.470 0.670 5.550 1.375 ;
        RECT  5.190 1.145 5.470 1.375 ;
        RECT  5.070 0.890 5.190 1.375 ;
        RECT  4.810 1.145 5.070 1.375 ;
        RECT  4.690 0.890 4.810 1.375 ;
        RECT  4.430 1.145 4.690 1.375 ;
        RECT  4.310 0.890 4.430 1.375 ;
        RECT  4.040 1.145 4.310 1.375 ;
        RECT  3.920 0.890 4.040 1.375 ;
        RECT  3.650 1.145 3.920 1.375 ;
        RECT  3.530 0.890 3.650 1.375 ;
        RECT  3.270 1.145 3.530 1.375 ;
        RECT  3.150 0.890 3.270 1.375 ;
        RECT  2.890 1.145 3.150 1.375 ;
        RECT  2.770 0.890 2.890 1.375 ;
        RECT  2.490 1.145 2.770 1.375 ;
        RECT  2.410 0.985 2.490 1.375 ;
        RECT  2.090 1.145 2.410 1.375 ;
        RECT  2.010 0.985 2.090 1.375 ;
        RECT  1.670 1.145 2.010 1.375 ;
        RECT  1.580 0.985 1.670 1.375 ;
        RECT  1.270 1.145 1.580 1.375 ;
        RECT  1.190 0.985 1.270 1.375 ;
        RECT  0.890 1.145 1.190 1.375 ;
        RECT  0.810 0.985 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.985 0.510 1.375 ;
        RECT  0.125 1.145 0.430 1.375 ;
        RECT  0.055 0.845 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.275 0.185 5.370 0.465 ;
        RECT  5.280 0.700 5.360 1.025 ;
        RECT  4.980 0.700 5.280 0.820 ;
        RECT  4.985 0.345 5.275 0.465 ;
        RECT  4.900 0.185 4.985 0.465 ;
        RECT  4.900 0.700 4.980 1.025 ;
        RECT  4.600 0.345 4.900 0.465 ;
        RECT  4.600 0.700 4.900 0.820 ;
        RECT  4.525 0.185 4.600 0.465 ;
        RECT  4.520 0.700 4.600 1.025 ;
        RECT  4.215 0.345 4.525 0.465 ;
        RECT  4.215 0.700 4.520 0.820 ;
        RECT  4.165 0.185 4.215 0.465 ;
        RECT  4.165 0.700 4.215 1.045 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.740 0.700 3.815 1.025 ;
        RECT  3.435 0.345 3.745 0.465 ;
        RECT  3.440 0.700 3.740 0.820 ;
        RECT  3.360 0.700 3.440 1.025 ;
        RECT  3.365 0.185 3.435 0.465 ;
        RECT  3.055 0.345 3.365 0.465 ;
        RECT  3.060 0.700 3.360 0.820 ;
        RECT  2.980 0.700 3.060 1.025 ;
        RECT  2.985 0.185 3.055 0.465 ;
        RECT  2.680 0.345 2.985 0.465 ;
        RECT  2.680 0.700 2.980 0.820 ;
        RECT  2.605 0.185 2.680 0.465 ;
        RECT  2.600 0.700 2.680 1.025 ;
        RECT  2.505 0.545 3.735 0.615 ;
        RECT  2.435 0.345 2.505 0.915 ;
        RECT  0.410 0.345 2.435 0.415 ;
        RECT  2.295 0.845 2.435 0.915 ;
        RECT  0.220 0.205 2.320 0.275 ;
        RECT  2.225 0.845 2.295 1.075 ;
        RECT  1.880 0.845 2.225 0.915 ;
        RECT  1.800 0.845 1.880 1.075 ;
        RECT  1.455 0.845 1.800 0.915 ;
        RECT  1.385 0.845 1.455 1.075 ;
        RECT  1.075 0.845 1.385 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.320 0.845 0.625 0.915 ;
        RECT  0.220 0.845 0.320 1.075 ;
    END
END AN2D16BWP40

MACRO AN2D1BWP40
    CLASS CORE ;
    FOREIGN AN2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.700 0.185 0.735 0.465 ;
        RECT  0.705 0.745 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.490 0.420 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 -0.115 0.840 0.115 ;
        RECT  0.455 -0.115 0.575 0.215 ;
        RECT  0.000 -0.115 0.455 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.150 1.145 0.480 1.375 ;
        RECT  0.070 0.965 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.520 0.655 0.640 ;
        RECT  0.535 0.305 0.605 0.915 ;
        RECT  0.165 0.305 0.535 0.375 ;
        RECT  0.340 0.845 0.535 0.915 ;
        RECT  0.260 0.845 0.340 1.050 ;
        RECT  0.070 0.195 0.165 0.375 ;
    END
END AN2D1BWP40

MACRO AN2D2BWP40
    CLASS CORE ;
    FOREIGN AN2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.785 ;
        RECT  0.715 0.355 0.735 0.455 ;
        RECT  0.715 0.715 0.735 0.785 ;
        RECT  0.645 0.185 0.715 0.455 ;
        RECT  0.645 0.715 0.715 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.395 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.280 ;
        RECT  0.550 -0.115 0.830 0.115 ;
        RECT  0.410 -0.115 0.550 0.265 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.865 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.985 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 0.525 0.665 0.635 ;
        RECT  0.470 0.345 0.540 0.915 ;
        RECT  0.145 0.345 0.470 0.415 ;
        RECT  0.340 0.845 0.470 0.915 ;
        RECT  0.220 0.845 0.340 1.055 ;
        RECT  0.035 0.195 0.145 0.415 ;
    END
END AN2D2BWP40

MACRO AN2D3BWP40
    CLASS CORE ;
    FOREIGN AN2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.268000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.185 1.205 0.475 ;
        RECT  1.130 0.700 1.205 1.045 ;
        RECT  1.015 0.355 1.135 0.475 ;
        RECT  1.015 0.700 1.130 0.820 ;
        RECT  0.805 0.355 1.015 0.820 ;
        RECT  0.715 0.355 0.805 0.475 ;
        RECT  0.715 0.700 0.805 0.820 ;
        RECT  0.645 0.185 0.715 0.475 ;
        RECT  0.645 0.700 0.715 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.395 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 -0.115 1.260 0.115 ;
        RECT  0.870 -0.115 0.950 0.280 ;
        RECT  0.550 -0.115 0.870 0.115 ;
        RECT  0.410 -0.115 0.550 0.265 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.145 1.260 1.375 ;
        RECT  0.850 0.890 0.970 1.375 ;
        RECT  0.540 1.145 0.850 1.375 ;
        RECT  0.420 0.985 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.185 1.205 0.475 ;
        RECT  1.130 0.700 1.205 1.045 ;
        RECT  1.085 0.355 1.135 0.475 ;
        RECT  1.085 0.700 1.130 0.820 ;
        RECT  0.715 0.355 0.735 0.475 ;
        RECT  0.715 0.700 0.735 0.820 ;
        RECT  0.645 0.185 0.715 0.475 ;
        RECT  0.645 0.700 0.715 1.045 ;
        RECT  0.540 0.545 0.700 0.615 ;
        RECT  0.470 0.345 0.540 0.915 ;
        RECT  0.145 0.345 0.470 0.415 ;
        RECT  0.340 0.845 0.470 0.915 ;
        RECT  0.220 0.845 0.340 1.055 ;
        RECT  0.035 0.195 0.145 0.415 ;
    END
END AN2D3BWP40

MACRO AN2D4BWP40
    CLASS CORE ;
    FOREIGN AN2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.185 1.515 0.485 ;
        RECT  1.445 0.700 1.515 1.030 ;
        RECT  1.435 0.355 1.445 0.485 ;
        RECT  1.435 0.700 1.445 0.820 ;
        RECT  1.225 0.355 1.435 0.820 ;
        RECT  1.135 0.355 1.225 0.475 ;
        RECT  1.135 0.700 1.225 0.820 ;
        RECT  1.065 0.185 1.135 0.475 ;
        RECT  1.065 0.700 1.135 1.030 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.780 0.640 ;
        RECT  0.625 0.520 0.695 0.790 ;
        RECT  0.245 0.720 0.625 0.790 ;
        RECT  0.170 0.495 0.245 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.480 0.545 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.730 -0.115 1.820 0.115 ;
        RECT  1.650 -0.115 1.730 0.475 ;
        RECT  1.350 -0.115 1.650 0.115 ;
        RECT  1.230 -0.115 1.350 0.280 ;
        RECT  0.940 -0.115 1.230 0.115 ;
        RECT  0.820 -0.115 0.940 0.265 ;
        RECT  0.130 -0.115 0.820 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.145 1.820 1.375 ;
        RECT  1.655 0.670 1.735 1.375 ;
        RECT  1.350 1.145 1.655 1.375 ;
        RECT  1.230 0.890 1.350 1.375 ;
        RECT  0.920 1.145 1.230 1.375 ;
        RECT  0.840 1.000 0.920 1.375 ;
        RECT  0.510 1.145 0.840 1.375 ;
        RECT  0.430 1.000 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.185 1.515 0.485 ;
        RECT  1.505 0.700 1.515 1.030 ;
        RECT  1.135 0.355 1.155 0.475 ;
        RECT  1.135 0.700 1.155 0.820 ;
        RECT  1.065 0.185 1.135 0.475 ;
        RECT  1.065 0.700 1.135 1.030 ;
        RECT  0.925 0.545 1.145 0.615 ;
        RECT  0.855 0.335 0.925 0.930 ;
        RECT  0.410 0.335 0.855 0.405 ;
        RECT  0.720 0.860 0.855 0.930 ;
        RECT  0.220 0.195 0.720 0.265 ;
        RECT  0.600 0.860 0.720 1.065 ;
        RECT  0.340 0.860 0.600 0.930 ;
        RECT  0.220 0.860 0.340 1.065 ;
    END
END AN2D4BWP40

MACRO AN2D6BWP40
    CLASS CORE ;
    FOREIGN AN2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.700 1.855 1.030 ;
        RECT  1.575 0.355 1.785 0.465 ;
        RECT  1.575 0.700 1.785 0.820 ;
        RECT  1.475 0.355 1.575 0.820 ;
        RECT  1.405 0.185 1.475 1.030 ;
        RECT  1.365 0.355 1.405 0.820 ;
        RECT  1.095 0.355 1.365 0.475 ;
        RECT  1.095 0.700 1.365 0.820 ;
        RECT  1.025 0.185 1.095 0.475 ;
        RECT  1.025 0.700 1.095 1.030 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.780 0.640 ;
        RECT  0.625 0.520 0.695 0.790 ;
        RECT  0.245 0.720 0.625 0.790 ;
        RECT  0.170 0.495 0.245 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.480 0.545 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.475 ;
        RECT  1.690 -0.115 1.970 0.115 ;
        RECT  1.570 -0.115 1.690 0.280 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.280 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.800 -0.115 0.920 0.265 ;
        RECT  0.130 -0.115 0.800 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.670 2.050 1.375 ;
        RECT  1.690 1.145 1.970 1.375 ;
        RECT  1.570 0.890 1.690 1.375 ;
        RECT  1.310 1.145 1.570 1.375 ;
        RECT  1.190 0.890 1.310 1.375 ;
        RECT  0.900 1.145 1.190 1.375 ;
        RECT  0.820 1.000 0.900 1.375 ;
        RECT  0.510 1.145 0.820 1.375 ;
        RECT  0.430 1.000 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.700 1.855 1.030 ;
        RECT  1.645 0.355 1.785 0.465 ;
        RECT  1.645 0.700 1.785 0.820 ;
        RECT  1.095 0.355 1.295 0.475 ;
        RECT  1.095 0.700 1.295 0.820 ;
        RECT  1.025 0.185 1.095 0.475 ;
        RECT  1.025 0.700 1.095 1.030 ;
        RECT  0.925 0.545 1.255 0.615 ;
        RECT  0.855 0.335 0.925 0.930 ;
        RECT  0.410 0.335 0.855 0.405 ;
        RECT  0.720 0.860 0.855 0.930 ;
        RECT  0.220 0.195 0.720 0.265 ;
        RECT  0.600 0.860 0.720 1.065 ;
        RECT  0.340 0.860 0.600 0.930 ;
        RECT  0.220 0.860 0.340 1.065 ;
    END
END AN2D6BWP40

MACRO AN2D8BWP40
    CLASS CORE ;
    FOREIGN AN2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.135 0.325 2.220 0.445 ;
        RECT  2.135 0.700 2.220 0.820 ;
        RECT  1.925 0.325 2.135 0.820 ;
        RECT  1.900 0.325 1.925 0.445 ;
        RECT  1.900 0.700 1.925 0.820 ;
        RECT  1.805 0.185 1.900 0.445 ;
        RECT  1.805 0.700 1.900 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.094400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.160 0.770 ;
        RECT  0.535 0.700 1.015 0.770 ;
        RECT  0.445 0.495 0.535 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.094400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.545 0.915 0.625 ;
        RECT  0.730 0.350 0.815 0.625 ;
        RECT  0.275 0.350 0.730 0.420 ;
        RECT  0.195 0.350 0.275 0.620 ;
        RECT  0.100 0.550 0.195 0.620 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.445 ;
        RECT  2.520 -0.115 2.810 0.115 ;
        RECT  2.400 -0.115 2.520 0.255 ;
        RECT  2.120 -0.115 2.400 0.115 ;
        RECT  2.000 -0.115 2.120 0.255 ;
        RECT  1.720 -0.115 2.000 0.115 ;
        RECT  1.600 -0.115 1.720 0.255 ;
        RECT  1.300 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.300 0.265 ;
        RECT  0.540 -0.115 1.220 0.115 ;
        RECT  0.420 -0.115 0.540 0.140 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.680 2.890 1.375 ;
        RECT  2.520 1.145 2.810 1.375 ;
        RECT  2.400 0.890 2.520 1.375 ;
        RECT  2.120 1.145 2.400 1.375 ;
        RECT  2.000 0.890 2.120 1.375 ;
        RECT  1.720 1.145 2.000 1.375 ;
        RECT  1.600 0.890 1.720 1.375 ;
        RECT  1.300 1.145 1.600 1.375 ;
        RECT  1.220 0.980 1.300 1.375 ;
        RECT  0.910 1.145 1.220 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.520 1.145 0.830 1.375 ;
        RECT  0.440 0.980 0.520 1.375 ;
        RECT  0.130 1.145 0.440 1.375 ;
        RECT  0.050 0.735 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.205 0.325 2.220 0.445 ;
        RECT  2.205 0.700 2.220 0.820 ;
        RECT  1.805 0.185 1.855 0.445 ;
        RECT  1.805 0.700 1.855 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        RECT  1.320 0.545 1.775 0.615 ;
        RECT  0.740 0.840 1.000 0.910 ;
        RECT  0.620 0.840 0.740 1.050 ;
        RECT  0.315 0.840 0.620 0.910 ;
        RECT  0.245 0.735 0.315 1.035 ;
        RECT  0.055 0.210 0.125 0.470 ;
        RECT  1.250 0.345 1.320 0.910 ;
        RECT  1.095 0.345 1.250 0.415 ;
        RECT  1.120 0.840 1.250 0.910 ;
        RECT  1.000 0.840 1.120 1.050 ;
        RECT  1.025 0.210 1.095 0.415 ;
        RECT  0.125 0.210 1.025 0.280 ;
    END
END AN2D8BWP40

MACRO AN3D0BWP40
    CLASS CORE ;
    FOREIGN AN3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.195 0.945 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.565 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 -0.115 0.980 0.115 ;
        RECT  0.630 -0.115 0.750 0.235 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.145 0.980 1.375 ;
        RECT  0.630 0.990 0.750 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.305 0.790 0.915 ;
        RECT  0.140 0.305 0.720 0.375 ;
        RECT  0.510 0.845 0.720 0.915 ;
        RECT  0.430 0.845 0.510 1.035 ;
        RECT  0.130 0.845 0.430 0.915 ;
        RECT  0.050 0.200 0.140 0.375 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END AN3D0BWP40

MACRO AN3D1BWP40
    CLASS CORE ;
    FOREIGN AN3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.195 0.945 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.565 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 -0.115 0.980 0.115 ;
        RECT  0.630 -0.115 0.750 0.235 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.145 0.980 1.375 ;
        RECT  0.630 0.990 0.750 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.305 0.790 0.915 ;
        RECT  0.140 0.305 0.720 0.375 ;
        RECT  0.510 0.845 0.720 0.915 ;
        RECT  0.430 0.845 0.510 1.035 ;
        RECT  0.130 0.845 0.430 0.915 ;
        RECT  0.050 0.200 0.140 0.375 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END AN3D1BWP40

MACRO AN3D2BWP40
    CLASS CORE ;
    FOREIGN AN3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.128000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.965 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.190 -0.115 1.260 0.115 ;
        RECT  1.110 -0.115 1.190 0.410 ;
        RECT  0.750 -0.115 1.110 0.115 ;
        RECT  0.630 -0.115 0.750 0.235 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.195 1.145 1.260 1.375 ;
        RECT  1.115 0.715 1.195 1.375 ;
        RECT  0.750 1.145 1.115 1.375 ;
        RECT  0.630 0.990 0.750 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.305 0.805 0.915 ;
        RECT  0.145 0.305 0.735 0.375 ;
        RECT  0.525 0.845 0.735 0.915 ;
        RECT  0.415 0.845 0.525 1.065 ;
        RECT  0.130 0.845 0.415 0.915 ;
        RECT  0.035 0.195 0.145 0.415 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END AN3D2BWP40

MACRO AN3D3BWP40
    CLASS CORE ;
    FOREIGN AN3D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.195 1.365 0.485 ;
        RECT  1.295 0.700 1.365 1.055 ;
        RECT  1.275 0.195 1.295 1.055 ;
        RECT  1.270 0.365 1.275 1.055 ;
        RECT  1.085 0.365 1.270 0.820 ;
        RECT  0.955 0.365 1.085 0.475 ;
        RECT  0.955 0.700 1.085 0.820 ;
        RECT  0.885 0.195 0.955 0.475 ;
        RECT  0.885 0.700 0.955 1.055 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 -0.115 1.400 0.115 ;
        RECT  1.060 -0.115 1.180 0.285 ;
        RECT  0.750 -0.115 1.060 0.115 ;
        RECT  0.630 -0.115 0.750 0.235 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.145 1.400 1.375 ;
        RECT  1.060 0.890 1.180 1.375 ;
        RECT  0.750 1.145 1.060 1.375 ;
        RECT  0.630 0.990 0.750 1.375 ;
        RECT  0.340 1.145 0.630 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.365 0.975 0.475 ;
        RECT  0.955 0.700 0.975 0.820 ;
        RECT  0.885 0.195 0.955 0.475 ;
        RECT  0.885 0.700 0.955 1.055 ;
        RECT  0.805 0.545 0.975 0.615 ;
        RECT  0.735 0.305 0.805 0.915 ;
        RECT  0.145 0.305 0.735 0.375 ;
        RECT  0.525 0.845 0.735 0.915 ;
        RECT  0.415 0.845 0.525 1.065 ;
        RECT  0.130 0.845 0.415 0.915 ;
        RECT  0.035 0.195 0.145 0.410 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END AN3D3BWP40

MACRO AN3D4BWP40
    CLASS CORE ;
    FOREIGN AN3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.185 1.945 0.465 ;
        RECT  1.875 0.700 1.945 1.065 ;
        RECT  1.855 0.355 1.875 0.465 ;
        RECT  1.855 0.700 1.875 0.820 ;
        RECT  1.645 0.355 1.855 0.820 ;
        RECT  1.535 0.355 1.645 0.465 ;
        RECT  1.535 0.700 1.645 0.820 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.700 1.535 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.495 1.225 0.790 ;
        RECT  0.260 0.720 1.105 0.790 ;
        RECT  0.170 0.495 0.260 0.790 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.350 1.000 0.640 ;
        RECT  0.430 0.350 0.875 0.420 ;
        RECT  0.350 0.350 0.430 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 -0.115 2.240 0.115 ;
        RECT  2.090 -0.115 2.170 0.475 ;
        RECT  1.760 -0.115 2.090 0.115 ;
        RECT  1.640 -0.115 1.760 0.275 ;
        RECT  1.320 -0.115 1.640 0.115 ;
        RECT  1.240 -0.115 1.320 0.265 ;
        RECT  0.125 -0.115 1.240 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.145 2.240 1.375 ;
        RECT  2.090 0.670 2.170 1.375 ;
        RECT  1.760 1.145 2.090 1.375 ;
        RECT  1.640 0.890 1.760 1.375 ;
        RECT  1.320 1.145 1.640 1.375 ;
        RECT  1.240 1.000 1.320 1.375 ;
        RECT  0.910 1.145 1.240 1.375 ;
        RECT  0.830 1.000 0.910 1.375 ;
        RECT  0.510 1.145 0.830 1.375 ;
        RECT  0.430 1.000 0.510 1.375 ;
        RECT  0.125 1.145 0.430 1.375 ;
        RECT  0.055 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.185 1.945 0.465 ;
        RECT  1.535 0.700 1.575 0.820 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.700 1.535 1.065 ;
        RECT  1.375 0.535 1.550 0.630 ;
        RECT  1.305 0.345 1.375 0.930 ;
        RECT  1.145 0.345 1.305 0.415 ;
        RECT  1.120 0.860 1.305 0.930 ;
        RECT  1.075 0.210 1.145 0.415 ;
        RECT  1.000 0.860 1.120 1.070 ;
        RECT  0.610 0.210 1.075 0.280 ;
        RECT  0.730 0.860 1.000 0.930 ;
        RECT  0.610 0.860 0.730 1.070 ;
        RECT  0.340 0.860 0.610 0.930 ;
        RECT  0.220 0.860 0.340 1.070 ;
        RECT  1.925 0.700 1.945 1.065 ;
        RECT  1.535 0.355 1.575 0.465 ;
    END
END AN3D4BWP40

MACRO AN3D6BWP40
    CLASS CORE ;
    FOREIGN AN3D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.185 2.275 0.465 ;
        RECT  2.205 0.700 2.275 1.065 ;
        RECT  1.995 0.355 2.205 0.465 ;
        RECT  1.995 0.700 2.205 0.820 ;
        RECT  1.895 0.355 1.995 0.820 ;
        RECT  1.825 0.185 1.895 1.065 ;
        RECT  1.785 0.355 1.825 0.820 ;
        RECT  1.495 0.355 1.785 0.465 ;
        RECT  1.495 0.700 1.785 0.820 ;
        RECT  1.425 0.185 1.495 0.465 ;
        RECT  1.425 0.700 1.495 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.495 1.185 0.790 ;
        RECT  0.260 0.720 1.105 0.790 ;
        RECT  0.170 0.495 0.260 0.790 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.350 1.000 0.640 ;
        RECT  0.430 0.350 0.875 0.420 ;
        RECT  0.350 0.350 0.430 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.110 -0.115 2.390 0.115 ;
        RECT  1.990 -0.115 2.110 0.275 ;
        RECT  1.720 -0.115 1.990 0.115 ;
        RECT  1.600 -0.115 1.720 0.275 ;
        RECT  1.300 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.300 0.265 ;
        RECT  0.125 -0.115 1.220 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.720 2.470 1.375 ;
        RECT  2.110 1.145 2.390 1.375 ;
        RECT  1.990 0.890 2.110 1.375 ;
        RECT  1.720 1.145 1.990 1.375 ;
        RECT  1.600 0.890 1.720 1.375 ;
        RECT  1.290 1.145 1.600 1.375 ;
        RECT  1.210 1.000 1.290 1.375 ;
        RECT  0.910 1.145 1.210 1.375 ;
        RECT  0.830 1.000 0.910 1.375 ;
        RECT  0.510 1.145 0.830 1.375 ;
        RECT  0.430 1.000 0.510 1.375 ;
        RECT  0.125 1.145 0.430 1.375 ;
        RECT  0.055 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.185 2.275 0.465 ;
        RECT  2.205 0.700 2.275 1.065 ;
        RECT  2.065 0.355 2.205 0.465 ;
        RECT  2.065 0.700 2.205 0.820 ;
        RECT  1.495 0.355 1.715 0.465 ;
        RECT  1.495 0.700 1.715 0.820 ;
        RECT  1.425 0.185 1.495 0.465 ;
        RECT  1.265 0.345 1.335 0.930 ;
        RECT  1.145 0.345 1.265 0.415 ;
        RECT  1.120 0.860 1.265 0.930 ;
        RECT  1.075 0.210 1.145 0.415 ;
        RECT  1.000 0.860 1.120 1.070 ;
        RECT  0.610 0.210 1.075 0.280 ;
        RECT  0.730 0.860 1.000 0.930 ;
        RECT  0.610 0.860 0.730 1.070 ;
        RECT  0.340 0.860 0.610 0.930 ;
        RECT  0.220 0.860 0.340 1.070 ;
        RECT  1.425 0.700 1.495 1.065 ;
        RECT  1.335 0.545 1.710 0.615 ;
    END
END AN3D6BWP40

MACRO AN3D8BWP40
    CLASS CORE ;
    FOREIGN AN3D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 0.700 3.260 1.025 ;
        RECT  3.185 0.185 3.255 0.465 ;
        RECT  2.855 0.345 3.185 0.465 ;
        RECT  2.855 0.700 3.180 0.820 ;
        RECT  2.835 0.185 2.855 0.465 ;
        RECT  2.835 0.700 2.855 1.045 ;
        RECT  2.785 0.185 2.835 1.045 ;
        RECT  2.780 0.345 2.785 1.045 ;
        RECT  2.625 0.345 2.780 0.820 ;
        RECT  2.455 0.345 2.625 0.465 ;
        RECT  2.460 0.700 2.625 0.820 ;
        RECT  2.380 0.700 2.460 1.025 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.055 0.345 2.385 0.465 ;
        RECT  2.060 0.700 2.380 0.820 ;
        RECT  1.980 0.700 2.060 1.025 ;
        RECT  1.985 0.185 2.055 0.465 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.760 ;
        RECT  1.295 0.495 1.575 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.495 1.225 0.765 ;
        RECT  0.780 0.495 1.145 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.540 0.625 ;
        RECT  0.175 0.495 0.245 0.760 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.465 ;
        RECT  3.080 -0.115 3.370 0.115 ;
        RECT  2.960 -0.115 3.080 0.265 ;
        RECT  2.680 -0.115 2.960 0.115 ;
        RECT  2.560 -0.115 2.680 0.265 ;
        RECT  2.280 -0.115 2.560 0.115 ;
        RECT  2.160 -0.115 2.280 0.265 ;
        RECT  1.855 -0.115 2.160 0.115 ;
        RECT  1.775 -0.115 1.855 0.400 ;
        RECT  1.460 -0.115 1.775 0.115 ;
        RECT  1.380 -0.115 1.460 0.275 ;
        RECT  0.000 -0.115 1.380 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.670 3.450 1.375 ;
        RECT  3.080 1.145 3.370 1.375 ;
        RECT  2.960 0.890 3.080 1.375 ;
        RECT  2.680 1.145 2.960 1.375 ;
        RECT  2.560 0.890 2.680 1.375 ;
        RECT  2.280 1.145 2.560 1.375 ;
        RECT  2.160 0.890 2.280 1.375 ;
        RECT  1.875 1.145 2.160 1.375 ;
        RECT  1.755 1.010 1.875 1.375 ;
        RECT  1.480 1.145 1.755 1.375 ;
        RECT  1.360 1.010 1.480 1.375 ;
        RECT  1.100 1.145 1.360 1.375 ;
        RECT  0.980 1.010 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 1.010 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.180 0.700 3.260 1.025 ;
        RECT  3.185 0.185 3.255 0.465 ;
        RECT  2.905 0.345 3.185 0.465 ;
        RECT  2.905 0.700 3.180 0.820 ;
        RECT  2.455 0.345 2.555 0.465 ;
        RECT  2.460 0.700 2.555 0.820 ;
        RECT  2.380 0.700 2.460 1.025 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.055 0.345 2.385 0.465 ;
        RECT  2.060 0.700 2.380 0.820 ;
        RECT  1.980 0.700 2.060 1.025 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.880 0.545 2.485 0.615 ;
        RECT  1.810 0.545 1.880 0.910 ;
        RECT  1.665 0.840 1.810 0.910 ;
        RECT  1.550 0.205 1.670 0.415 ;
        RECT  1.555 0.840 1.665 1.075 ;
        RECT  1.285 0.840 1.555 0.910 ;
        RECT  1.265 0.345 1.550 0.415 ;
        RECT  1.175 0.840 1.285 1.075 ;
        RECT  1.195 0.185 1.265 0.415 ;
        RECT  0.790 0.345 1.195 0.415 ;
        RECT  0.905 0.840 1.175 0.910 ;
        RECT  0.225 0.205 1.100 0.275 ;
        RECT  0.795 0.840 0.905 1.075 ;
        RECT  0.700 0.840 0.795 0.910 ;
        RECT  0.620 0.345 0.700 0.910 ;
        RECT  0.145 0.345 0.620 0.415 ;
        RECT  0.525 0.840 0.620 0.910 ;
        RECT  0.415 0.840 0.525 1.075 ;
        RECT  0.145 0.840 0.415 0.910 ;
        RECT  0.035 0.195 0.145 0.415 ;
        RECT  0.035 0.840 0.145 1.075 ;
    END
END AN3D8BWP40

MACRO AN4D0BWP40
    CLASS CORE ;
    FOREIGN AN4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.054000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.195 1.225 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.850 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.635 0.665 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.450 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.115 1.260 0.115 ;
        RECT  0.880 -0.115 1.000 0.210 ;
        RECT  0.000 -0.115 0.880 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.145 1.260 1.375 ;
        RECT  0.880 0.985 1.000 1.375 ;
        RECT  0.550 1.145 0.880 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.985 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 0.280 1.050 0.915 ;
        RECT  0.140 0.280 0.980 0.350 ;
        RECT  0.750 0.845 0.980 0.915 ;
        RECT  0.670 0.845 0.750 1.045 ;
        RECT  0.320 0.845 0.670 0.915 ;
        RECT  0.240 0.845 0.320 1.045 ;
        RECT  0.040 0.200 0.140 0.350 ;
    END
END AN4D0BWP40

MACRO AN4D1BWP40
    CLASS CORE ;
    FOREIGN AN4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.108000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.195 1.225 1.065 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.850 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.635 0.665 0.765 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.115 1.260 0.115 ;
        RECT  0.880 -0.115 1.000 0.210 ;
        RECT  0.000 -0.115 0.880 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.145 1.260 1.375 ;
        RECT  0.880 0.985 1.000 1.375 ;
        RECT  0.550 1.145 0.880 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.985 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 0.280 1.050 0.915 ;
        RECT  0.035 0.280 0.980 0.350 ;
        RECT  0.750 0.845 0.980 0.915 ;
        RECT  0.670 0.845 0.750 1.045 ;
        RECT  0.320 0.845 0.670 0.915 ;
        RECT  0.240 0.845 0.320 1.045 ;
    END
END AN4D1BWP40

MACRO AN4D2BWP40
    CLASS CORE ;
    FOREIGN AN4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.495 1.225 0.765 ;
        RECT  1.090 0.195 1.160 1.065 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.850 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.275 -0.115 1.345 0.415 ;
        RECT  0.970 -0.115 1.275 0.115 ;
        RECT  0.850 -0.115 0.970 0.210 ;
        RECT  0.000 -0.115 0.850 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.270 0.860 1.345 1.375 ;
        RECT  0.980 1.145 1.270 1.375 ;
        RECT  0.860 0.985 0.980 1.375 ;
        RECT  0.550 1.145 0.860 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.125 1.145 0.430 1.375 ;
        RECT  0.050 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.280 1.020 0.915 ;
        RECT  0.145 0.280 0.950 0.350 ;
        RECT  0.765 0.845 0.950 0.915 ;
        RECT  0.655 0.845 0.765 1.065 ;
        RECT  0.335 0.845 0.655 0.915 ;
        RECT  0.225 0.845 0.335 1.065 ;
        RECT  0.035 0.195 0.145 0.410 ;
    END
END AN4D2BWP40

MACRO AN4D3BWP40
    CLASS CORE ;
    FOREIGN AN4D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.195 1.505 0.455 ;
        RECT  1.435 0.710 1.505 1.045 ;
        RECT  1.415 0.195 1.435 1.045 ;
        RECT  1.225 0.355 1.415 0.810 ;
        RECT  1.110 0.355 1.225 0.455 ;
        RECT  1.110 0.710 1.225 0.810 ;
        RECT  1.040 0.195 1.110 0.455 ;
        RECT  1.040 0.710 1.110 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.810 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.320 0.240 ;
        RECT  0.930 -0.115 1.200 0.115 ;
        RECT  0.810 -0.115 0.930 0.210 ;
        RECT  0.000 -0.115 0.810 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.540 1.375 ;
        RECT  1.200 0.890 1.320 1.375 ;
        RECT  0.930 1.145 1.200 1.375 ;
        RECT  0.810 0.985 0.930 1.375 ;
        RECT  0.530 1.145 0.810 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.110 0.355 1.155 0.455 ;
        RECT  1.110 0.710 1.155 0.810 ;
        RECT  1.040 0.195 1.110 0.455 ;
        RECT  1.040 0.710 1.110 1.045 ;
        RECT  0.970 0.545 1.110 0.615 ;
        RECT  0.900 0.280 0.970 0.915 ;
        RECT  0.145 0.280 0.900 0.350 ;
        RECT  0.715 0.845 0.900 0.915 ;
        RECT  0.605 0.845 0.715 1.065 ;
        RECT  0.335 0.845 0.605 0.915 ;
        RECT  0.225 0.845 0.335 1.065 ;
        RECT  0.035 0.195 0.145 0.410 ;
    END
END AN4D3BWP40

MACRO AN4D4BWP40
    CLASS CORE ;
    FOREIGN AN4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.249600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.395 0.465 ;
        RECT  2.325 0.690 2.395 1.025 ;
        RECT  2.275 0.355 2.325 0.465 ;
        RECT  2.275 0.690 2.325 0.790 ;
        RECT  2.065 0.355 2.275 0.790 ;
        RECT  2.015 0.355 2.065 0.465 ;
        RECT  2.005 0.690 2.065 0.790 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.690 2.005 1.025 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.520 1.650 0.915 ;
        RECT  0.245 0.845 1.565 0.915 ;
        RECT  0.165 0.495 0.245 0.915 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.430 0.765 ;
        RECT  0.420 0.345 1.295 0.415 ;
        RECT  0.315 0.345 0.420 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.495 1.225 0.765 ;
        RECT  0.665 0.695 1.120 0.765 ;
        RECT  0.575 0.495 0.665 0.765 ;
        RECT  0.545 0.495 0.575 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.985 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.475 ;
        RECT  2.230 -0.115 2.530 0.115 ;
        RECT  2.110 -0.115 2.230 0.275 ;
        RECT  1.780 -0.115 2.110 0.115 ;
        RECT  1.700 -0.115 1.780 0.300 ;
        RECT  0.125 -0.115 1.700 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.700 2.610 1.375 ;
        RECT  2.230 1.145 2.530 1.375 ;
        RECT  2.110 0.870 2.230 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.125 1.800 1.375 ;
        RECT  1.360 1.145 1.680 1.375 ;
        RECT  1.240 1.125 1.360 1.375 ;
        RECT  0.940 1.145 1.240 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.530 1.145 0.820 1.375 ;
        RECT  0.410 1.125 0.530 1.375 ;
        RECT  0.125 1.145 0.410 1.375 ;
        RECT  0.055 0.980 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.185 2.395 0.465 ;
        RECT  2.345 0.690 2.395 1.025 ;
        RECT  1.945 0.185 1.995 0.465 ;
        RECT  1.935 0.690 1.995 1.025 ;
        RECT  1.855 0.545 1.970 0.615 ;
        RECT  1.785 0.370 1.855 1.055 ;
        RECT  1.600 0.370 1.785 0.440 ;
        RECT  0.220 0.985 1.785 1.055 ;
        RECT  1.530 0.205 1.600 0.440 ;
        RECT  0.825 0.205 1.530 0.275 ;
    END
END AN4D4BWP40

MACRO AN4D6BWP40
    CLASS CORE ;
    FOREIGN AN4D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.366600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.185 2.780 0.470 ;
        RECT  2.700 0.710 2.780 1.025 ;
        RECT  2.415 0.355 2.700 0.470 ;
        RECT  2.415 0.710 2.700 0.810 ;
        RECT  2.405 0.355 2.415 0.810 ;
        RECT  2.400 0.185 2.405 0.810 ;
        RECT  2.325 0.185 2.400 1.025 ;
        RECT  2.205 0.355 2.325 0.810 ;
        RECT  2.015 0.355 2.205 0.465 ;
        RECT  2.005 0.710 2.205 0.810 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.710 2.005 1.025 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.520 1.650 0.915 ;
        RECT  0.245 0.845 1.565 0.915 ;
        RECT  0.165 0.495 0.245 0.915 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.430 0.765 ;
        RECT  0.420 0.345 1.295 0.415 ;
        RECT  0.315 0.345 0.420 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.495 1.225 0.765 ;
        RECT  0.665 0.695 1.120 0.765 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.545 0.495 0.595 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.985 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 -0.115 3.080 0.115 ;
        RECT  2.915 -0.115 2.995 0.475 ;
        RECT  2.610 -0.115 2.915 0.115 ;
        RECT  2.490 -0.115 2.610 0.275 ;
        RECT  2.230 -0.115 2.490 0.115 ;
        RECT  2.110 -0.115 2.230 0.275 ;
        RECT  1.780 -0.115 2.110 0.115 ;
        RECT  1.700 -0.115 1.780 0.300 ;
        RECT  0.125 -0.115 1.700 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 1.145 3.080 1.375 ;
        RECT  2.915 0.695 2.995 1.375 ;
        RECT  2.610 1.145 2.915 1.375 ;
        RECT  2.490 0.890 2.610 1.375 ;
        RECT  2.230 1.145 2.490 1.375 ;
        RECT  2.110 0.890 2.230 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.125 1.800 1.375 ;
        RECT  1.360 1.145 1.680 1.375 ;
        RECT  1.240 1.125 1.360 1.375 ;
        RECT  0.940 1.145 1.240 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.530 1.145 0.820 1.375 ;
        RECT  0.410 1.125 0.530 1.375 ;
        RECT  0.125 1.145 0.410 1.375 ;
        RECT  0.055 0.980 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.700 0.185 2.780 0.470 ;
        RECT  2.700 0.710 2.780 1.025 ;
        RECT  2.485 0.355 2.700 0.470 ;
        RECT  2.485 0.710 2.700 0.810 ;
        RECT  2.015 0.355 2.135 0.465 ;
        RECT  2.005 0.710 2.135 0.810 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.710 2.005 1.025 ;
        RECT  1.855 0.545 2.130 0.615 ;
        RECT  1.785 0.370 1.855 1.055 ;
        RECT  1.600 0.370 1.785 0.440 ;
        RECT  0.220 0.985 1.785 1.055 ;
        RECT  1.530 0.205 1.600 0.440 ;
        RECT  0.825 0.205 1.530 0.275 ;
    END
END AN4D6BWP40

MACRO AN4D8BWP40
    CLASS CORE ;
    FOREIGN AN4D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.496000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.660 0.695 3.750 0.995 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.355 0.345 3.665 0.465 ;
        RECT  3.360 0.695 3.660 0.815 ;
        RECT  3.280 0.695 3.360 0.995 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.255 0.345 3.285 0.465 ;
        RECT  3.255 0.695 3.280 0.815 ;
        RECT  3.045 0.345 3.255 0.815 ;
        RECT  2.975 0.345 3.045 0.465 ;
        RECT  2.975 0.695 3.045 0.815 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.900 0.695 2.975 0.995 ;
        RECT  2.595 0.345 2.905 0.465 ;
        RECT  2.600 0.695 2.900 0.815 ;
        RECT  2.520 0.695 2.600 0.995 ;
        RECT  2.525 0.185 2.595 0.465 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.145 0.495 2.215 0.765 ;
        RECT  1.855 0.495 2.145 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.785 0.765 ;
        RECT  1.365 0.495 1.715 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.135 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.175 0.495 0.455 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.975 -0.115 4.060 0.115 ;
        RECT  3.895 -0.115 3.975 0.465 ;
        RECT  3.570 -0.115 3.895 0.115 ;
        RECT  3.450 -0.115 3.570 0.275 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.275 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.275 ;
        RECT  2.410 -0.115 2.690 0.115 ;
        RECT  2.330 -0.115 2.410 0.455 ;
        RECT  2.030 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.030 0.275 ;
        RECT  0.000 -0.115 1.950 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.975 1.145 4.060 1.375 ;
        RECT  3.895 0.720 3.975 1.375 ;
        RECT  3.570 1.145 3.895 1.375 ;
        RECT  3.450 0.885 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.885 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.885 2.810 1.375 ;
        RECT  2.410 1.145 2.690 1.375 ;
        RECT  2.330 0.985 2.410 1.375 ;
        RECT  2.030 1.145 2.330 1.375 ;
        RECT  1.950 0.985 2.030 1.375 ;
        RECT  1.650 1.145 1.950 1.375 ;
        RECT  1.570 0.985 1.650 1.375 ;
        RECT  1.270 1.145 1.570 1.375 ;
        RECT  1.190 0.985 1.270 1.375 ;
        RECT  0.890 1.145 1.190 1.375 ;
        RECT  0.810 0.985 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.985 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.720 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.660 0.695 3.750 0.995 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.355 0.345 3.665 0.465 ;
        RECT  3.360 0.695 3.660 0.815 ;
        RECT  3.325 0.695 3.360 0.995 ;
        RECT  3.325 0.185 3.355 0.465 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.900 0.695 2.975 0.995 ;
        RECT  2.595 0.345 2.905 0.465 ;
        RECT  2.600 0.695 2.900 0.815 ;
        RECT  2.520 0.695 2.600 0.995 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.400 0.545 2.965 0.615 ;
        RECT  2.320 0.545 2.400 0.915 ;
        RECT  2.240 0.845 2.320 0.915 ;
        RECT  2.120 0.205 2.240 0.415 ;
        RECT  2.120 0.845 2.240 1.055 ;
        RECT  1.855 0.345 2.120 0.415 ;
        RECT  1.860 0.845 2.120 0.915 ;
        RECT  1.740 0.845 1.860 1.055 ;
        RECT  1.745 0.205 1.855 0.415 ;
        RECT  1.360 0.205 1.745 0.275 ;
        RECT  1.480 0.845 1.740 0.915 ;
        RECT  0.790 0.345 1.665 0.415 ;
        RECT  1.360 0.845 1.480 1.055 ;
        RECT  1.100 0.845 1.360 0.915 ;
        RECT  0.225 0.205 1.100 0.275 ;
        RECT  0.980 0.845 1.100 1.055 ;
        RECT  0.720 0.845 0.980 0.915 ;
        RECT  0.665 0.845 0.720 1.055 ;
        RECT  0.600 0.345 0.665 1.055 ;
        RECT  0.595 0.345 0.600 0.915 ;
        RECT  0.145 0.345 0.595 0.415 ;
        RECT  0.340 0.845 0.595 0.915 ;
        RECT  0.220 0.845 0.340 1.055 ;
        RECT  0.035 0.195 0.145 0.415 ;
    END
END AN4D8BWP40

MACRO ANTENNABWP40
    CLASS CORE ;
    FOREIGN ANTENNABWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN I
        ANTENNADIFFAREA 0.120400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.190 0.245 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
END ANTENNABWP40

MACRO AO211D0BWP40
    CLASS CORE ;
    FOREIGN AO211D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.064000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.190 1.225 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.455 0.835 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.940 0.210 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.210 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 1.260 1.375 ;
        RECT  0.820 1.050 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.290 1.020 0.920 ;
        RECT  0.720 0.290 0.950 0.360 ;
        RECT  0.220 0.850 0.950 0.920 ;
        RECT  0.640 0.215 0.720 0.360 ;
        RECT  0.130 0.290 0.640 0.360 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.050 0.195 0.130 0.360 ;
        RECT  0.050 0.915 0.130 1.065 ;
    END
END AO211D0BWP40

MACRO AO211D1BWP40
    CLASS CORE ;
    FOREIGN AO211D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.128000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.190 1.225 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.455 0.875 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.630 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.630 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.940 0.210 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.210 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 1.260 1.375 ;
        RECT  0.820 0.995 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.290 1.020 0.920 ;
        RECT  0.720 0.290 0.950 0.360 ;
        RECT  0.220 0.850 0.950 0.920 ;
        RECT  0.640 0.215 0.720 0.360 ;
        RECT  0.130 0.290 0.640 0.360 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.050 0.195 0.130 0.360 ;
        RECT  0.050 0.915 0.130 1.065 ;
    END
END AO211D1BWP40

MACRO AO211D2BWP40
    CLASS CORE ;
    FOREIGN AO211D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.165 0.495 1.225 0.765 ;
        RECT  1.090 0.190 1.165 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.475 0.835 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.275 -0.115 1.345 0.400 ;
        RECT  0.940 -0.115 1.275 0.115 ;
        RECT  0.820 -0.115 0.940 0.210 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.210 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.275 0.860 1.345 1.375 ;
        RECT  0.940 1.145 1.275 1.375 ;
        RECT  0.820 0.995 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.945 0.290 1.015 0.920 ;
        RECT  0.735 0.290 0.945 0.360 ;
        RECT  0.220 0.850 0.945 0.920 ;
        RECT  0.625 0.195 0.735 0.405 ;
        RECT  0.145 0.290 0.625 0.360 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.035 0.195 0.145 0.405 ;
        RECT  0.050 0.915 0.130 1.065 ;
    END
END AO211D2BWP40

MACRO AO211D4BWP40
    CLASS CORE ;
    FOREIGN AO211D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.237000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.415 1.030 ;
        RECT  2.205 0.355 2.325 0.905 ;
        RECT  2.015 0.355 2.205 0.465 ;
        RECT  2.015 0.745 2.205 0.905 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.745 2.015 1.030 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.555 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.495 0.805 0.765 ;
        RECT  0.245 0.695 0.700 0.765 ;
        RECT  0.170 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.485 0.490 1.680 0.775 ;
        RECT  0.995 0.705 1.485 0.775 ;
        RECT  0.875 0.495 0.995 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.495 1.375 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.475 ;
        RECT  2.230 -0.115 2.530 0.115 ;
        RECT  2.110 -0.115 2.230 0.260 ;
        RECT  1.830 -0.115 2.110 0.115 ;
        RECT  1.750 -0.115 1.830 0.260 ;
        RECT  1.650 -0.115 1.750 0.115 ;
        RECT  1.570 -0.115 1.650 0.260 ;
        RECT  0.890 -0.115 1.570 0.115 ;
        RECT  0.810 -0.115 0.890 0.265 ;
        RECT  0.510 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.720 2.610 1.375 ;
        RECT  2.230 1.145 2.530 1.375 ;
        RECT  2.110 0.985 2.230 1.375 ;
        RECT  1.850 1.145 2.110 1.375 ;
        RECT  1.730 1.125 1.850 1.375 ;
        RECT  0.530 1.145 1.730 1.375 ;
        RECT  0.410 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.015 0.355 2.135 0.465 ;
        RECT  2.015 0.745 2.135 0.905 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.745 2.015 1.030 ;
        RECT  1.860 0.550 2.125 0.625 ;
        RECT  1.790 0.345 1.860 1.055 ;
        RECT  0.720 0.345 1.790 0.415 ;
        RECT  0.985 0.985 1.790 1.055 ;
        RECT  0.905 0.845 1.670 0.915 ;
        RECT  0.980 0.200 1.480 0.275 ;
        RECT  0.795 0.845 0.905 1.075 ;
        RECT  0.600 0.205 0.720 0.415 ;
        RECT  0.340 0.345 0.600 0.415 ;
        RECT  0.220 0.205 0.340 0.415 ;
        RECT  0.035 0.845 0.145 1.075 ;
        RECT  0.145 0.845 0.795 0.915 ;
    END
END AO211D4BWP40

MACRO AO21D0BWP40
    CLASS CORE ;
    FOREIGN AO21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.195 0.945 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.590 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.210 ;
        RECT  0.130 -0.115 0.640 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 1.005 0.760 1.375 ;
        RECT  0.000 1.145 0.640 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.280 0.790 0.915 ;
        RECT  0.525 0.280 0.720 0.350 ;
        RECT  0.220 0.845 0.720 0.915 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.455 0.205 0.525 0.350 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO21D0BWP40

MACRO AO21D1BWP40
    CLASS CORE ;
    FOREIGN AO21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.195 0.945 1.065 ;
        RECT  0.855 0.955 0.860 1.065 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.590 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.210 ;
        RECT  0.130 -0.115 0.640 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 1.005 0.760 1.375 ;
        RECT  0.000 1.145 0.640 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.280 0.790 0.915 ;
        RECT  0.525 0.280 0.720 0.350 ;
        RECT  0.220 0.845 0.720 0.915 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.455 0.205 0.525 0.350 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO21D1BWP40

MACRO AO21D2BWP40
    CLASS CORE ;
    FOREIGN AO21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.950 1.065 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 -0.115 1.260 0.115 ;
        RECT  1.095 -0.115 1.175 0.415 ;
        RECT  0.720 -0.115 1.095 0.115 ;
        RECT  0.600 -0.115 0.720 0.210 ;
        RECT  0.130 -0.115 0.600 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.145 1.260 1.375 ;
        RECT  1.110 0.710 1.180 1.375 ;
        RECT  0.720 1.145 1.110 1.375 ;
        RECT  0.600 1.005 0.720 1.375 ;
        RECT  0.000 1.145 0.600 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.280 0.805 0.915 ;
        RECT  0.405 0.280 0.735 0.350 ;
        RECT  0.200 0.845 0.735 0.915 ;
        RECT  0.130 0.995 0.530 1.065 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO21D2BWP40

MACRO AO21D4BWP40
    CLASS CORE ;
    FOREIGN AO21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.185 1.935 0.465 ;
        RECT  1.865 0.710 1.935 1.030 ;
        RECT  1.855 0.355 1.865 0.465 ;
        RECT  1.855 0.710 1.865 0.830 ;
        RECT  1.645 0.355 1.855 0.830 ;
        RECT  1.535 0.355 1.645 0.465 ;
        RECT  1.535 0.710 1.645 0.830 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.710 1.535 1.030 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.495 1.225 0.780 ;
        RECT  0.245 0.710 1.100 0.780 ;
        RECT  0.145 0.495 0.245 0.780 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.845 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.345 1.020 0.640 ;
        RECT  0.430 0.345 0.915 0.415 ;
        RECT  0.315 0.345 0.430 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.145 -0.115 2.240 0.115 ;
        RECT  2.065 -0.115 2.145 0.475 ;
        RECT  1.760 -0.115 2.065 0.115 ;
        RECT  1.640 -0.115 1.760 0.280 ;
        RECT  1.340 -0.115 1.640 0.115 ;
        RECT  1.220 -0.115 1.340 0.135 ;
        RECT  0.730 -0.115 1.220 0.115 ;
        RECT  0.610 -0.115 0.730 0.135 ;
        RECT  0.125 -0.115 0.610 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 1.145 2.240 1.375 ;
        RECT  2.075 0.680 2.155 1.375 ;
        RECT  1.760 1.145 2.075 1.375 ;
        RECT  1.640 0.910 1.760 1.375 ;
        RECT  1.340 1.145 1.640 1.375 ;
        RECT  1.220 0.990 1.340 1.375 ;
        RECT  0.125 1.145 1.220 1.375 ;
        RECT  0.055 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.185 1.935 0.465 ;
        RECT  1.925 0.710 1.935 1.030 ;
        RECT  1.535 0.355 1.575 0.465 ;
        RECT  1.535 0.710 1.575 0.830 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.710 1.535 1.030 ;
        RECT  1.375 0.550 1.535 0.630 ;
        RECT  1.305 0.205 1.375 0.920 ;
        RECT  0.220 0.205 1.305 0.275 ;
        RECT  0.415 0.850 1.305 0.920 ;
        RECT  0.335 0.990 1.120 1.060 ;
        RECT  0.225 0.850 0.335 1.060 ;
    END
END AO21D4BWP40

MACRO AO221D0BWP40
    CLASS CORE ;
    FOREIGN AO221D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.062000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.195 1.505 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.155 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.795 0.695 0.875 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.195 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.540 0.115 ;
        RECT  1.160 -0.115 1.280 0.230 ;
        RECT  0.690 -0.115 1.160 0.115 ;
        RECT  0.610 -0.115 0.690 0.275 ;
        RECT  0.140 -0.115 0.610 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.160 0.990 1.280 1.375 ;
        RECT  0.000 1.145 1.160 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.345 1.330 0.640 ;
        RECT  1.065 0.345 1.260 0.415 ;
        RECT  0.995 0.195 1.065 0.415 ;
        RECT  0.990 0.845 1.060 1.030 ;
        RECT  0.505 0.345 0.995 0.415 ;
        RECT  0.595 0.845 0.990 0.915 ;
        RECT  0.125 0.995 0.900 1.065 ;
        RECT  0.435 0.195 0.505 0.415 ;
        RECT  0.335 0.345 0.435 0.415 ;
        RECT  0.265 0.345 0.335 0.915 ;
        RECT  0.210 0.845 0.265 0.915 ;
        RECT  0.055 0.925 0.125 1.065 ;
    END
END AO221D0BWP40

MACRO AO221D1BWP40
    CLASS CORE ;
    FOREIGN AO221D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.195 1.505 1.075 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.155 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.805 0.625 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.795 0.695 0.875 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.195 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.540 0.115 ;
        RECT  1.160 -0.115 1.280 0.230 ;
        RECT  0.690 -0.115 1.160 0.115 ;
        RECT  0.610 -0.115 0.690 0.275 ;
        RECT  0.140 -0.115 0.610 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.160 0.910 1.280 1.375 ;
        RECT  0.000 1.145 1.160 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.270 0.345 1.340 0.640 ;
        RECT  1.065 0.345 1.270 0.415 ;
        RECT  0.995 0.195 1.065 0.415 ;
        RECT  0.990 0.845 1.060 1.030 ;
        RECT  0.505 0.345 0.995 0.415 ;
        RECT  0.595 0.845 0.990 0.915 ;
        RECT  0.125 0.995 0.900 1.065 ;
        RECT  0.435 0.195 0.505 0.415 ;
        RECT  0.335 0.345 0.435 0.415 ;
        RECT  0.265 0.345 0.335 0.915 ;
        RECT  0.210 0.845 0.265 0.915 ;
        RECT  0.055 0.755 0.125 1.065 ;
    END
END AO221D1BWP40

MACRO AO221D2BWP40
    CLASS CORE ;
    FOREIGN AO221D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.495 1.785 0.640 ;
        RECT  1.500 0.195 1.595 1.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.775 1.365 0.905 ;
        RECT  1.170 0.495 1.245 0.905 ;
        RECT  1.155 0.495 1.170 0.695 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.805 0.625 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 -0.115 1.820 0.115 ;
        RECT  1.685 -0.115 1.755 0.415 ;
        RECT  1.370 -0.115 1.685 0.115 ;
        RECT  1.250 -0.115 1.370 0.230 ;
        RECT  0.720 -0.115 1.250 0.115 ;
        RECT  0.640 -0.115 0.720 0.275 ;
        RECT  0.125 -0.115 0.640 0.115 ;
        RECT  0.055 -0.115 0.125 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 1.145 1.820 1.375 ;
        RECT  1.685 0.720 1.755 1.375 ;
        RECT  1.370 1.145 1.685 1.375 ;
        RECT  1.250 0.985 1.370 1.375 ;
        RECT  0.000 1.145 1.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.345 0.345 1.425 0.640 ;
        RECT  1.095 0.345 1.345 0.415 ;
        RECT  1.025 0.195 1.095 0.415 ;
        RECT  1.020 0.845 1.090 1.030 ;
        RECT  0.525 0.345 1.025 0.415 ;
        RECT  0.620 0.845 1.020 0.915 ;
        RECT  0.125 0.995 0.930 1.065 ;
        RECT  0.455 0.195 0.525 0.415 ;
        RECT  0.385 0.345 0.455 0.415 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.220 0.845 0.315 0.915 ;
        RECT  0.055 0.915 0.125 1.065 ;
    END
END AO221D2BWP40

MACRO AO221D4BWP40
    CLASS CORE ;
    FOREIGN AO221D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.185 2.835 0.465 ;
        RECT  2.825 0.745 2.835 1.030 ;
        RECT  2.765 0.185 2.825 1.030 ;
        RECT  2.625 0.355 2.765 0.830 ;
        RECT  2.455 0.355 2.625 0.465 ;
        RECT  2.455 0.745 2.625 0.830 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.745 2.455 1.030 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.100 0.630 ;
        RECT  1.855 0.495 1.925 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.495 1.645 0.775 ;
        RECT  1.085 0.705 1.515 0.775 ;
        RECT  0.990 0.495 1.085 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.780 0.640 ;
        RECT  0.625 0.520 0.695 0.775 ;
        RECT  0.245 0.705 0.625 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.485 0.545 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.475 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.550 -0.115 2.670 0.280 ;
        RECT  2.265 -0.115 2.550 0.115 ;
        RECT  2.195 -0.115 2.265 0.275 ;
        RECT  1.820 -0.115 2.195 0.115 ;
        RECT  1.820 0.195 1.910 0.265 ;
        RECT  1.700 -0.115 1.820 0.265 ;
        RECT  0.940 -0.115 1.700 0.115 ;
        RECT  1.610 0.195 1.700 0.265 ;
        RECT  0.820 -0.115 0.940 0.260 ;
        RECT  0.130 -0.115 0.820 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.715 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.550 0.910 2.670 1.375 ;
        RECT  2.270 1.145 2.550 1.375 ;
        RECT  2.190 0.730 2.270 1.375 ;
        RECT  1.890 1.145 2.190 1.375 ;
        RECT  1.810 0.985 1.890 1.375 ;
        RECT  0.000 1.145 1.810 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.455 0.355 2.555 0.465 ;
        RECT  2.455 0.745 2.555 0.830 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.745 2.455 1.030 ;
        RECT  2.305 0.545 2.440 0.615 ;
        RECT  2.235 0.345 2.305 0.615 ;
        RECT  2.075 0.345 2.235 0.415 ;
        RECT  1.985 0.845 2.095 1.060 ;
        RECT  2.005 0.185 2.075 0.415 ;
        RECT  0.920 0.345 2.005 0.415 ;
        RECT  1.040 0.845 1.985 0.915 ;
        RECT  0.130 0.985 1.730 1.055 ;
        RECT  1.020 0.195 1.540 0.265 ;
        RECT  0.850 0.345 0.920 0.915 ;
        RECT  0.415 0.345 0.850 0.415 ;
        RECT  0.220 0.845 0.850 0.915 ;
        RECT  0.335 0.205 0.740 0.275 ;
        RECT  0.225 0.205 0.335 0.415 ;
        RECT  0.050 0.875 0.130 1.055 ;
    END
END AO221D4BWP40

MACRO AO222D0BWP40
    CLASS CORE ;
    FOREIGN AO222D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.064000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.185 1.785 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.635 1.505 0.765 ;
        RECT  1.295 0.495 1.375 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.630 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.620 0.610 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.115 1.820 0.115 ;
        RECT  1.400 -0.115 1.520 0.240 ;
        RECT  0.540 -0.115 1.400 0.115 ;
        RECT  0.420 -0.115 0.540 0.220 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.145 1.820 1.375 ;
        RECT  1.425 1.010 1.545 1.375 ;
        RECT  1.130 1.145 1.425 1.375 ;
        RECT  1.010 1.000 1.130 1.375 ;
        RECT  0.000 1.145 1.010 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.500 0.315 1.590 0.555 ;
        RECT  1.130 0.315 1.500 0.385 ;
        RECT  1.220 0.855 1.300 1.040 ;
        RECT  0.220 0.855 1.220 0.925 ;
        RECT  0.830 0.225 1.130 0.385 ;
        RECT  0.130 0.995 0.930 1.065 ;
        RECT  0.760 0.315 0.830 0.385 ;
        RECT  0.690 0.315 0.760 0.785 ;
        RECT  0.140 0.315 0.690 0.385 ;
        RECT  0.630 0.685 0.690 0.785 ;
        RECT  0.055 0.195 0.140 0.385 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO222D0BWP40

MACRO AO222D1BWP40
    CLASS CORE ;
    FOREIGN AO222D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.128000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.185 1.785 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.710 1.505 0.780 ;
        RECT  1.295 0.495 1.375 0.780 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.620 0.610 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.115 1.820 0.115 ;
        RECT  1.400 -0.115 1.520 0.240 ;
        RECT  0.540 -0.115 1.400 0.115 ;
        RECT  0.420 -0.115 0.540 0.220 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.145 1.820 1.375 ;
        RECT  1.425 0.870 1.545 1.375 ;
        RECT  1.130 1.145 1.425 1.375 ;
        RECT  1.010 1.000 1.130 1.375 ;
        RECT  0.000 1.145 1.010 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.500 0.315 1.590 0.640 ;
        RECT  1.130 0.315 1.500 0.385 ;
        RECT  0.220 0.855 1.320 0.925 ;
        RECT  0.830 0.225 1.130 0.385 ;
        RECT  0.130 0.995 0.930 1.065 ;
        RECT  0.760 0.315 0.830 0.385 ;
        RECT  0.690 0.315 0.760 0.785 ;
        RECT  0.140 0.315 0.690 0.385 ;
        RECT  0.630 0.685 0.690 0.785 ;
        RECT  0.055 0.195 0.140 0.385 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO222D1BWP40

MACRO AO222D2BWP40
    CLASS CORE ;
    FOREIGN AO222D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.735 0.495 1.785 0.765 ;
        RECT  1.645 0.185 1.735 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.710 1.500 0.780 ;
        RECT  1.295 0.495 1.375 0.780 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.620 0.610 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.830 -0.115 1.910 0.395 ;
        RECT  1.515 -0.115 1.830 0.115 ;
        RECT  1.375 -0.115 1.515 0.240 ;
        RECT  0.540 -0.115 1.375 0.115 ;
        RECT  0.420 -0.115 0.540 0.220 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.830 0.860 1.910 1.375 ;
        RECT  1.540 1.145 1.830 1.375 ;
        RECT  1.420 0.870 1.540 1.375 ;
        RECT  1.130 1.145 1.420 1.375 ;
        RECT  1.010 1.000 1.130 1.375 ;
        RECT  0.000 1.145 1.010 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.485 0.315 1.565 0.640 ;
        RECT  1.130 0.315 1.485 0.385 ;
        RECT  1.205 0.855 1.315 1.065 ;
        RECT  0.220 0.855 1.205 0.925 ;
        RECT  0.830 0.225 1.130 0.385 ;
        RECT  0.130 0.995 0.930 1.065 ;
        RECT  0.760 0.315 0.830 0.385 ;
        RECT  0.690 0.315 0.760 0.785 ;
        RECT  0.145 0.315 0.690 0.385 ;
        RECT  0.630 0.685 0.690 0.785 ;
        RECT  0.035 0.195 0.145 0.410 ;
        RECT  0.050 0.925 0.130 1.065 ;
    END
END AO222D2BWP40

MACRO AO222D4BWP40
    CLASS CORE ;
    FOREIGN AO222D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.185 3.255 0.485 ;
        RECT  3.245 0.710 3.255 1.045 ;
        RECT  3.185 0.185 3.245 1.045 ;
        RECT  3.045 0.355 3.185 0.830 ;
        RECT  2.875 0.355 3.045 0.485 ;
        RECT  2.875 0.710 3.045 0.830 ;
        RECT  2.805 0.185 2.875 0.485 ;
        RECT  2.805 0.710 2.875 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.495 2.540 0.640 ;
        RECT  2.385 0.495 2.485 0.775 ;
        RECT  1.920 0.705 2.385 0.775 ;
        RECT  1.795 0.495 1.920 0.775 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.270 0.630 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.670 0.775 ;
        RECT  1.085 0.705 1.575 0.775 ;
        RECT  0.985 0.495 1.085 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.490 1.505 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.765 0.640 ;
        RECT  0.625 0.520 0.695 0.775 ;
        RECT  0.245 0.705 0.625 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.475 ;
        RECT  3.090 -0.115 3.370 0.115 ;
        RECT  2.970 -0.115 3.090 0.280 ;
        RECT  2.680 -0.115 2.970 0.115 ;
        RECT  2.560 -0.115 2.680 0.210 ;
        RECT  1.820 -0.115 2.560 0.115 ;
        RECT  1.820 0.195 1.910 0.265 ;
        RECT  1.700 -0.115 1.820 0.265 ;
        RECT  0.940 -0.115 1.700 0.115 ;
        RECT  1.610 0.195 1.700 0.265 ;
        RECT  0.820 -0.115 0.940 0.210 ;
        RECT  0.130 -0.115 0.820 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.720 3.450 1.375 ;
        RECT  3.090 1.145 3.370 1.375 ;
        RECT  2.970 0.900 3.090 1.375 ;
        RECT  2.660 1.145 2.970 1.375 ;
        RECT  2.580 0.745 2.660 1.375 ;
        RECT  2.270 1.145 2.580 1.375 ;
        RECT  2.190 0.985 2.270 1.375 ;
        RECT  1.890 1.145 2.190 1.375 ;
        RECT  1.810 0.985 1.890 1.375 ;
        RECT  0.000 1.145 1.810 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.875 0.355 2.975 0.485 ;
        RECT  2.875 0.710 2.975 0.830 ;
        RECT  2.805 0.185 2.875 0.485 ;
        RECT  2.805 0.710 2.875 1.045 ;
        RECT  2.645 0.345 2.735 0.640 ;
        RECT  0.915 0.345 2.645 0.415 ;
        RECT  1.980 0.195 2.480 0.265 ;
        RECT  2.360 0.845 2.480 1.055 ;
        RECT  2.100 0.845 2.360 0.915 ;
        RECT  1.980 0.845 2.100 1.055 ;
        RECT  1.040 0.845 1.980 0.915 ;
        RECT  0.130 0.985 1.730 1.055 ;
        RECT  1.030 0.195 1.540 0.265 ;
        RECT  0.845 0.345 0.915 0.915 ;
        RECT  0.410 0.345 0.845 0.415 ;
        RECT  0.220 0.845 0.845 0.915 ;
        RECT  0.210 0.195 0.735 0.265 ;
        RECT  0.050 0.875 0.130 1.055 ;
    END
END AO222D4BWP40

MACRO AO22D0BWP40
    CLASS CORE ;
    FOREIGN AO22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.054000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.185 1.365 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 -0.115 1.400 0.115 ;
        RECT  1.055 -0.115 1.125 0.260 ;
        RECT  0.910 -0.115 1.055 0.115 ;
        RECT  0.835 -0.115 0.910 0.260 ;
        RECT  0.130 -0.115 0.835 0.115 ;
        RECT  0.050 -0.115 0.130 0.260 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 1.145 1.400 1.375 ;
        RECT  1.055 0.990 1.125 1.375 ;
        RECT  0.340 1.145 1.055 1.375 ;
        RECT  0.220 1.045 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.095 0.330 1.165 0.915 ;
        RECT  0.705 0.330 1.095 0.400 ;
        RECT  0.605 0.845 1.095 0.915 ;
        RECT  0.505 0.995 0.930 1.065 ;
        RECT  0.635 0.195 0.705 0.400 ;
        RECT  0.415 0.195 0.635 0.265 ;
        RECT  0.435 0.905 0.505 1.065 ;
        RECT  0.125 0.905 0.435 0.975 ;
        RECT  0.055 0.905 0.125 1.065 ;
    END
END AO22D0BWP40

MACRO AO22D1BWP40
    CLASS CORE ;
    FOREIGN AO22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.108000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.185 1.365 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 -0.115 1.400 0.115 ;
        RECT  1.055 -0.115 1.125 0.260 ;
        RECT  0.910 -0.115 1.055 0.115 ;
        RECT  0.835 -0.115 0.910 0.260 ;
        RECT  0.130 -0.115 0.835 0.115 ;
        RECT  0.050 -0.115 0.130 0.260 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.125 1.145 1.400 1.375 ;
        RECT  1.055 0.990 1.125 1.375 ;
        RECT  0.340 1.145 1.055 1.375 ;
        RECT  0.220 1.045 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.095 0.330 1.165 0.915 ;
        RECT  0.705 0.330 1.095 0.400 ;
        RECT  0.605 0.845 1.095 0.915 ;
        RECT  0.505 0.995 0.930 1.065 ;
        RECT  0.635 0.195 0.705 0.400 ;
        RECT  0.415 0.195 0.635 0.265 ;
        RECT  0.435 0.905 0.505 1.065 ;
        RECT  0.125 0.905 0.435 0.975 ;
        RECT  0.055 0.905 0.125 1.065 ;
    END
END AO22D1BWP40

MACRO AO22D2BWP40
    CLASS CORE ;
    FOREIGN AO22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 0.495 1.365 0.765 ;
        RECT  1.230 0.185 1.300 1.065 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 -0.115 1.540 0.115 ;
        RECT  1.415 -0.115 1.485 0.415 ;
        RECT  1.095 -0.115 1.415 0.115 ;
        RECT  1.025 -0.115 1.095 0.260 ;
        RECT  0.900 -0.115 1.025 0.115 ;
        RECT  0.825 -0.115 0.900 0.260 ;
        RECT  0.130 -0.115 0.825 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 1.145 1.540 1.375 ;
        RECT  1.415 0.860 1.485 1.375 ;
        RECT  1.095 1.145 1.415 1.375 ;
        RECT  1.025 0.990 1.095 1.375 ;
        RECT  0.340 1.145 1.025 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.065 0.330 1.135 0.915 ;
        RECT  0.705 0.330 1.065 0.400 ;
        RECT  0.605 0.845 1.065 0.915 ;
        RECT  0.505 0.995 0.920 1.065 ;
        RECT  0.635 0.195 0.705 0.400 ;
        RECT  0.415 0.195 0.635 0.265 ;
        RECT  0.435 0.845 0.505 1.065 ;
        RECT  0.125 0.845 0.435 0.915 ;
        RECT  0.055 0.845 0.125 1.065 ;
    END
END AO22D2BWP40

MACRO AO22D4BWP40
    CLASS CORE ;
    FOREIGN AO22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.395 0.485 ;
        RECT  2.325 0.710 2.395 1.045 ;
        RECT  2.275 0.355 2.325 0.485 ;
        RECT  2.275 0.710 2.325 0.830 ;
        RECT  2.065 0.355 2.275 0.830 ;
        RECT  2.015 0.355 2.065 0.485 ;
        RECT  2.015 0.710 2.065 0.830 ;
        RECT  1.945 0.185 2.015 0.485 ;
        RECT  1.945 0.710 2.015 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.520 0.790 0.775 ;
        RECT  0.245 0.705 0.670 0.775 ;
        RECT  0.135 0.495 0.245 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.645 0.775 ;
        RECT  0.995 0.705 1.505 0.775 ;
        RECT  0.870 0.495 0.995 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.410 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.475 ;
        RECT  2.230 -0.115 2.510 0.115 ;
        RECT  2.110 -0.115 2.230 0.280 ;
        RECT  1.825 -0.115 2.110 0.115 ;
        RECT  1.755 -0.115 1.825 0.260 ;
        RECT  1.645 -0.115 1.755 0.115 ;
        RECT  1.575 -0.115 1.645 0.260 ;
        RECT  0.885 -0.115 1.575 0.115 ;
        RECT  0.815 -0.115 0.885 0.240 ;
        RECT  0.130 -0.115 0.815 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.720 2.590 1.375 ;
        RECT  2.230 1.145 2.510 1.375 ;
        RECT  2.110 0.900 2.230 1.375 ;
        RECT  1.825 1.145 2.110 1.375 ;
        RECT  1.755 0.990 1.825 1.375 ;
        RECT  0.700 1.145 1.755 1.375 ;
        RECT  0.620 0.985 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 0.985 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.185 2.395 0.485 ;
        RECT  2.345 0.710 2.395 1.045 ;
        RECT  1.945 0.185 1.995 0.485 ;
        RECT  1.945 0.710 1.995 1.045 ;
        RECT  1.780 0.345 1.860 0.915 ;
        RECT  0.400 0.345 1.780 0.415 ;
        RECT  0.980 0.845 1.780 0.915 ;
        RECT  0.885 0.985 1.670 1.055 ;
        RECT  0.980 0.195 1.480 0.265 ;
        RECT  0.815 0.845 0.885 1.055 ;
        RECT  0.530 0.845 0.815 0.915 ;
        RECT  0.220 0.195 0.720 0.265 ;
        RECT  0.410 0.845 0.530 1.055 ;
        RECT  0.145 0.845 0.410 0.915 ;
        RECT  0.035 0.845 0.145 1.055 ;
    END
END AO22D4BWP40

MACRO AO31D0BWP40
    CLASS CORE ;
    FOREIGN AO31D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.054000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.190 1.225 1.045 ;
        RECT  1.120 0.190 1.155 0.470 ;
        RECT  1.120 0.760 1.155 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.485 0.850 0.770 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.415 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.010 -0.115 1.260 0.115 ;
        RECT  0.890 -0.115 1.010 0.210 ;
        RECT  0.140 -0.115 0.890 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 1.145 1.260 1.375 ;
        RECT  0.905 0.995 0.985 1.375 ;
        RECT  0.000 1.145 0.905 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.520 1.060 0.640 ;
        RECT  0.970 0.280 1.040 0.915 ;
        RECT  0.780 0.280 0.970 0.350 ;
        RECT  0.125 0.845 0.970 0.915 ;
        RECT  0.220 0.985 0.795 1.055 ;
        RECT  0.660 0.215 0.780 0.350 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END AO31D0BWP40

MACRO AO31D1BWP40
    CLASS CORE ;
    FOREIGN AO31D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.108000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.190 1.225 1.045 ;
        RECT  1.120 0.190 1.155 0.470 ;
        RECT  1.120 0.760 1.155 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.485 0.850 0.770 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.415 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.010 -0.115 1.260 0.115 ;
        RECT  0.890 -0.115 1.010 0.210 ;
        RECT  0.140 -0.115 0.890 0.115 ;
        RECT  0.040 -0.115 0.140 0.390 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 1.145 1.260 1.375 ;
        RECT  0.905 0.995 0.985 1.375 ;
        RECT  0.000 1.145 0.905 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.520 1.060 0.640 ;
        RECT  0.970 0.335 1.040 0.915 ;
        RECT  0.775 0.335 0.970 0.405 ;
        RECT  0.125 0.845 0.970 0.915 ;
        RECT  0.220 0.985 0.795 1.055 ;
        RECT  0.665 0.195 0.775 0.405 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END AO31D1BWP40

MACRO AO31D2BWP40
    CLASS CORE ;
    FOREIGN AO31D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.495 1.365 0.630 ;
        RECT  1.120 0.190 1.190 1.060 ;
        RECT  1.085 0.190 1.120 0.470 ;
        RECT  1.085 0.775 1.120 1.060 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.485 0.840 0.770 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.415 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 0.495 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.275 -0.115 1.345 0.415 ;
        RECT  0.985 -0.115 1.275 0.115 ;
        RECT  0.865 -0.115 0.985 0.210 ;
        RECT  0.140 -0.115 0.865 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.275 0.720 1.345 1.375 ;
        RECT  0.965 1.145 1.275 1.375 ;
        RECT  0.885 0.995 0.965 1.375 ;
        RECT  0.000 1.145 0.885 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.005 0.520 1.025 0.640 ;
        RECT  0.935 0.335 1.005 0.915 ;
        RECT  0.790 0.335 0.935 0.405 ;
        RECT  0.125 0.845 0.935 0.915 ;
        RECT  0.680 0.195 0.790 0.405 ;
        RECT  0.220 0.985 0.785 1.055 ;
        RECT  0.055 0.845 0.125 1.025 ;
    END
END AO31D2BWP40

MACRO AO31D4BWP40
    CLASS CORE ;
    FOREIGN AO31D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.395 0.465 ;
        RECT  2.325 0.700 2.395 1.035 ;
        RECT  2.275 0.355 2.325 0.465 ;
        RECT  2.275 0.700 2.325 0.820 ;
        RECT  2.065 0.355 2.275 0.820 ;
        RECT  2.015 0.355 2.065 0.465 ;
        RECT  2.015 0.700 2.065 0.820 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.700 2.015 1.035 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.660 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.495 1.225 0.640 ;
        RECT  1.050 0.495 1.120 0.785 ;
        RECT  0.245 0.715 1.050 0.785 ;
        RECT  0.125 0.495 0.245 0.785 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.345 0.975 0.625 ;
        RECT  0.385 0.345 0.865 0.415 ;
        RECT  0.315 0.345 0.385 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.700 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.475 ;
        RECT  2.230 -0.115 2.510 0.115 ;
        RECT  2.110 -0.115 2.230 0.250 ;
        RECT  1.830 -0.115 2.110 0.115 ;
        RECT  1.750 -0.115 1.830 0.260 ;
        RECT  1.650 -0.115 1.750 0.115 ;
        RECT  1.570 -0.115 1.650 0.265 ;
        RECT  1.290 -0.115 1.570 0.115 ;
        RECT  1.200 -0.115 1.290 0.280 ;
        RECT  0.130 -0.115 1.200 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.720 2.590 1.375 ;
        RECT  2.230 1.145 2.510 1.375 ;
        RECT  2.110 0.890 2.230 1.375 ;
        RECT  1.850 1.145 2.110 1.375 ;
        RECT  1.750 0.855 1.850 1.375 ;
        RECT  1.360 0.855 1.750 0.925 ;
        RECT  0.000 1.145 1.750 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.185 2.395 0.465 ;
        RECT  2.345 0.700 2.395 1.035 ;
        RECT  1.945 0.185 1.995 0.465 ;
        RECT  1.945 0.700 1.995 1.035 ;
        RECT  1.855 0.550 1.985 0.630 ;
        RECT  1.785 0.350 1.855 0.780 ;
        RECT  1.120 0.350 1.785 0.420 ;
        RECT  1.270 0.710 1.785 0.780 ;
        RECT  0.125 0.995 1.670 1.065 ;
        RECT  1.200 0.710 1.270 0.925 ;
        RECT  0.220 0.855 1.200 0.925 ;
        RECT  1.050 0.195 1.120 0.420 ;
        RECT  0.600 0.195 1.050 0.265 ;
        RECT  0.055 0.880 0.125 1.065 ;
    END
END AO31D4BWP40

MACRO AO32D0BWP40
    CLASS CORE ;
    FOREIGN AO32D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.068000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.190 1.645 1.045 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.115 1.680 0.115 ;
        RECT  1.295 -0.115 1.395 0.260 ;
        RECT  1.170 -0.115 1.295 0.115 ;
        RECT  1.070 -0.115 1.170 0.260 ;
        RECT  0.130 -0.115 1.070 0.115 ;
        RECT  0.050 -0.115 0.130 0.270 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.145 1.680 1.375 ;
        RECT  1.285 1.005 1.405 1.375 ;
        RECT  0.980 1.145 1.285 1.375 ;
        RECT  0.860 1.125 0.980 1.375 ;
        RECT  0.000 1.145 0.860 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.345 1.420 0.915 ;
        RECT  0.765 0.345 1.350 0.415 ;
        RECT  0.125 0.845 1.350 0.915 ;
        RECT  0.230 0.985 1.180 1.055 ;
        RECT  0.650 0.210 0.765 0.415 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO32D0BWP40

MACRO AO32D1BWP40
    CLASS CORE ;
    FOREIGN AO32D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.190 1.645 1.065 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.115 1.680 0.115 ;
        RECT  1.295 -0.115 1.395 0.260 ;
        RECT  1.165 -0.115 1.295 0.115 ;
        RECT  1.075 -0.115 1.165 0.260 ;
        RECT  0.130 -0.115 1.075 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.145 1.680 1.375 ;
        RECT  1.285 1.005 1.405 1.375 ;
        RECT  0.980 1.145 1.285 1.375 ;
        RECT  0.860 1.125 0.980 1.375 ;
        RECT  0.000 1.145 0.860 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.345 1.420 0.915 ;
        RECT  0.765 0.345 1.350 0.415 ;
        RECT  0.125 0.845 1.350 0.915 ;
        RECT  0.230 0.985 1.180 1.055 ;
        RECT  0.655 0.195 0.765 0.415 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO32D1BWP40

MACRO AO32D2BWP40
    CLASS CORE ;
    FOREIGN AO32D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.495 1.645 0.765 ;
        RECT  1.500 0.190 1.570 1.065 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.760 0.415 ;
        RECT  1.385 -0.115 1.690 0.115 ;
        RECT  1.305 -0.115 1.385 0.260 ;
        RECT  1.160 -0.115 1.305 0.115 ;
        RECT  1.090 -0.115 1.160 0.260 ;
        RECT  0.130 -0.115 1.090 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.145 1.820 1.375 ;
        RECT  1.690 0.860 1.760 1.375 ;
        RECT  1.405 1.145 1.690 1.375 ;
        RECT  1.285 1.005 1.405 1.375 ;
        RECT  0.980 1.145 1.285 1.375 ;
        RECT  0.860 1.125 0.980 1.375 ;
        RECT  0.000 1.145 0.860 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.345 1.420 0.915 ;
        RECT  0.765 0.345 1.350 0.415 ;
        RECT  0.125 0.845 1.350 0.915 ;
        RECT  0.230 0.985 1.180 1.055 ;
        RECT  0.655 0.205 0.765 0.415 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END AO32D2BWP40

MACRO AO32D4BWP40
    CLASS CORE ;
    FOREIGN AO32D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.185 2.835 0.485 ;
        RECT  2.765 0.710 2.835 1.050 ;
        RECT  2.695 0.355 2.765 0.485 ;
        RECT  2.695 0.710 2.765 0.830 ;
        RECT  2.485 0.355 2.695 0.830 ;
        RECT  2.455 0.355 2.485 0.485 ;
        RECT  2.455 0.710 2.485 0.830 ;
        RECT  2.385 0.185 2.455 0.485 ;
        RECT  2.385 0.710 2.455 1.050 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 0.495 2.095 0.770 ;
        RECT  1.420 0.700 1.940 0.770 ;
        RECT  1.295 0.495 1.420 0.770 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.495 1.870 0.630 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.070 0.495 1.145 0.775 ;
        RECT  0.245 0.705 1.070 0.775 ;
        RECT  0.110 0.495 0.245 0.775 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 0.975 0.630 ;
        RECT  0.425 0.345 0.875 0.415 ;
        RECT  0.315 0.345 0.425 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.475 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.550 -0.115 2.670 0.280 ;
        RECT  2.265 -0.115 2.550 0.115 ;
        RECT  2.195 -0.115 2.265 0.260 ;
        RECT  2.085 -0.115 2.195 0.115 ;
        RECT  2.015 -0.115 2.085 0.260 ;
        RECT  1.330 -0.115 2.015 0.115 ;
        RECT  1.250 -0.115 1.330 0.265 ;
        RECT  0.130 -0.115 1.250 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.720 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.550 0.900 2.670 1.375 ;
        RECT  2.270 1.145 2.550 1.375 ;
        RECT  2.190 0.990 2.270 1.375 ;
        RECT  1.910 1.145 2.190 1.375 ;
        RECT  1.790 1.125 1.910 1.375 ;
        RECT  1.510 1.145 1.790 1.375 ;
        RECT  1.390 1.125 1.510 1.375 ;
        RECT  0.000 1.145 1.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.185 2.835 0.485 ;
        RECT  2.765 0.710 2.835 1.050 ;
        RECT  2.385 0.185 2.415 0.485 ;
        RECT  2.385 0.710 2.415 1.050 ;
        RECT  2.225 0.345 2.295 0.915 ;
        RECT  1.170 0.345 2.225 0.415 ;
        RECT  0.220 0.845 2.225 0.915 ;
        RECT  0.125 0.985 2.110 1.055 ;
        RECT  1.415 0.195 1.925 0.265 ;
        RECT  1.090 0.195 1.170 0.415 ;
        RECT  0.600 0.195 1.090 0.265 ;
        RECT  0.055 0.900 0.125 1.055 ;
    END
END AO32D4BWP40

MACRO AO33D0BWP40
    CLASS CORE ;
    FOREIGN AO33D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.070000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.185 1.645 1.075 ;
        RECT  1.535 0.185 1.575 0.255 ;
        RECT  1.530 0.985 1.575 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.365 0.625 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.450 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 -0.115 1.680 0.115 ;
        RECT  1.280 -0.115 1.400 0.210 ;
        RECT  0.130 -0.115 1.280 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.145 1.680 1.375 ;
        RECT  1.280 0.985 1.400 1.375 ;
        RECT  0.940 1.145 1.280 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.435 0.320 1.505 0.915 ;
        RECT  1.165 0.320 1.435 0.390 ;
        RECT  0.130 0.845 1.435 0.915 ;
        RECT  1.095 0.215 1.165 0.390 ;
        RECT  0.220 0.985 1.150 1.055 ;
        RECT  0.610 0.215 1.095 0.285 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO33D0BWP40

MACRO AO33D1BWP40
    CLASS CORE ;
    FOREIGN AO33D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.128000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.195 1.645 1.065 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.455 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 -0.115 1.680 0.115 ;
        RECT  1.280 -0.115 1.400 0.210 ;
        RECT  0.130 -0.115 1.280 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.145 1.680 1.375 ;
        RECT  1.280 0.985 1.400 1.375 ;
        RECT  0.940 1.145 1.280 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.395 0.285 1.465 0.915 ;
        RECT  0.610 0.285 1.395 0.355 ;
        RECT  0.130 0.845 1.395 0.915 ;
        RECT  0.220 0.985 1.150 1.055 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO33D1BWP40

MACRO AO33D2BWP40
    CLASS CORE ;
    FOREIGN AO33D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.495 1.645 0.765 ;
        RECT  1.510 0.195 1.580 1.065 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.285 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.455 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.215 0.525 0.345 ;
        RECT  0.315 0.215 0.385 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.115 1.820 0.115 ;
        RECT  1.695 -0.115 1.765 0.405 ;
        RECT  1.395 -0.115 1.695 0.115 ;
        RECT  1.275 -0.115 1.395 0.210 ;
        RECT  0.130 -0.115 1.275 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.695 0.860 1.770 1.375 ;
        RECT  1.395 1.145 1.695 1.375 ;
        RECT  1.275 0.985 1.395 1.375 ;
        RECT  0.940 1.145 1.275 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.355 0.285 1.425 0.915 ;
        RECT  0.610 0.285 1.355 0.355 ;
        RECT  0.130 0.845 1.355 0.915 ;
        RECT  0.220 0.985 1.150 1.055 ;
        RECT  0.050 0.845 0.130 0.995 ;
    END
END AO33D2BWP40

MACRO AO33D4BWP40
    CLASS CORE ;
    FOREIGN AO33D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.185 0.185 3.255 0.485 ;
        RECT  3.185 0.710 3.255 1.050 ;
        RECT  3.115 0.355 3.185 0.485 ;
        RECT  3.115 0.710 3.185 0.830 ;
        RECT  2.905 0.355 3.115 0.830 ;
        RECT  2.875 0.355 2.905 0.485 ;
        RECT  2.875 0.710 2.905 0.830 ;
        RECT  2.805 0.185 2.875 0.485 ;
        RECT  2.805 0.710 2.875 1.050 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 0.495 2.485 0.780 ;
        RECT  1.505 0.710 2.360 0.780 ;
        RECT  1.375 0.495 1.505 0.780 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.345 2.225 0.640 ;
        RECT  1.675 0.345 2.135 0.415 ;
        RECT  1.575 0.345 1.675 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 2.065 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.225 0.780 ;
        RECT  0.195 0.710 1.130 0.780 ;
        RECT  0.125 0.520 0.195 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.345 1.015 0.640 ;
        RECT  0.405 0.345 0.915 0.415 ;
        RECT  0.305 0.345 0.405 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.565 0.495 0.845 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.475 ;
        RECT  3.090 -0.115 3.370 0.115 ;
        RECT  2.970 -0.115 3.090 0.280 ;
        RECT  2.685 -0.115 2.970 0.115 ;
        RECT  2.615 -0.115 2.685 0.280 ;
        RECT  2.505 -0.115 2.615 0.115 ;
        RECT  2.435 -0.115 2.505 0.260 ;
        RECT  1.345 -0.115 2.435 0.115 ;
        RECT  1.275 -0.115 1.345 0.275 ;
        RECT  0.130 -0.115 1.275 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.720 3.450 1.375 ;
        RECT  3.090 1.145 3.370 1.375 ;
        RECT  2.970 0.900 3.090 1.375 ;
        RECT  2.685 1.145 2.970 1.375 ;
        RECT  2.615 0.990 2.685 1.375 ;
        RECT  2.340 1.145 2.615 1.375 ;
        RECT  2.210 1.130 2.340 1.375 ;
        RECT  1.950 1.145 2.210 1.375 ;
        RECT  1.830 1.130 1.950 1.375 ;
        RECT  1.550 1.145 1.830 1.375 ;
        RECT  1.430 1.130 1.550 1.375 ;
        RECT  0.000 1.145 1.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.185 3.255 0.485 ;
        RECT  3.185 0.710 3.255 1.050 ;
        RECT  2.805 0.185 2.835 0.485 ;
        RECT  2.805 0.710 2.835 1.050 ;
        RECT  2.645 0.350 2.715 0.920 ;
        RECT  2.365 0.350 2.645 0.420 ;
        RECT  0.220 0.850 2.645 0.920 ;
        RECT  0.125 0.990 2.530 1.060 ;
        RECT  2.295 0.205 2.365 0.420 ;
        RECT  1.505 0.205 2.295 0.275 ;
        RECT  1.435 0.205 1.505 0.415 ;
        RECT  1.165 0.345 1.435 0.415 ;
        RECT  1.095 0.205 1.165 0.415 ;
        RECT  0.640 0.205 1.095 0.275 ;
        RECT  0.055 0.910 0.125 1.060 ;
    END
END AO33D4BWP40

MACRO AOI211D0BWP40
    CLASS CORE ;
    FOREIGN AOI211D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.092625 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.195 0.750 0.360 ;
        RECT  0.525 0.290 0.650 0.360 ;
        RECT  0.455 0.290 0.525 0.915 ;
        RECT  0.145 0.290 0.455 0.360 ;
        RECT  0.220 0.845 0.455 0.915 ;
        RECT  0.035 0.200 0.145 0.360 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.775 0.805 0.915 ;
        RECT  0.595 0.485 0.665 0.915 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.440 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.280 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.210 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.990 0.930 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.995 0.560 1.065 ;
        RECT  0.055 0.915 0.125 1.065 ;
    END
END AOI211D0BWP40

MACRO AOI211D1BWP40
    CLASS CORE ;
    FOREIGN AOI211D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.169250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.290 0.760 0.360 ;
        RECT  0.455 0.290 0.525 0.915 ;
        RECT  0.145 0.290 0.455 0.360 ;
        RECT  0.220 0.845 0.455 0.915 ;
        RECT  0.035 0.215 0.145 0.360 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.775 0.805 0.915 ;
        RECT  0.595 0.485 0.665 0.915 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.440 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.420 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.210 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.990 0.930 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.995 0.560 1.065 ;
        RECT  0.055 0.915 0.125 1.065 ;
    END
END AOI211D1BWP40

MACRO AOI211D2BWP40
    CLASS CORE ;
    FOREIGN AOI211D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.292500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.845 1.540 0.925 ;
        RECT  1.235 0.185 1.365 0.415 ;
        RECT  0.930 0.345 1.235 0.415 ;
        RECT  0.930 0.775 1.085 0.925 ;
        RECT  0.845 0.345 0.930 0.925 ;
        RECT  0.710 0.345 0.845 0.415 ;
        RECT  0.765 0.775 0.845 0.925 ;
        RECT  0.595 0.185 0.710 0.415 ;
        RECT  0.340 0.345 0.595 0.415 ;
        RECT  0.220 0.205 0.340 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.765 0.640 ;
        RECT  0.625 0.520 0.695 0.775 ;
        RECT  0.245 0.705 0.625 0.775 ;
        RECT  0.130 0.495 0.245 0.775 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.655 0.775 ;
        RECT  1.225 0.705 1.575 0.775 ;
        RECT  1.155 0.495 1.225 0.775 ;
        RECT  1.000 0.495 1.155 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.505 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.115 1.820 0.115 ;
        RECT  1.685 -0.115 1.765 0.420 ;
        RECT  0.915 -0.115 1.685 0.115 ;
        RECT  0.845 -0.115 0.915 0.275 ;
        RECT  0.505 -0.115 0.845 0.115 ;
        RECT  0.435 -0.115 0.505 0.275 ;
        RECT  0.130 -0.115 0.435 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.145 1.820 1.375 ;
        RECT  0.410 0.990 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.635 0.905 1.705 1.065 ;
        RECT  0.695 0.995 1.635 1.065 ;
        RECT  0.625 0.845 0.695 1.065 ;
        RECT  0.125 0.845 0.625 0.915 ;
        RECT  0.055 0.845 0.125 0.995 ;
    END
END AOI211D2BWP40

MACRO AOI211D3BWP40
    CLASS CORE ;
    FOREIGN AOI211D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.458300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.355 2.270 0.425 ;
        RECT  1.085 0.845 1.125 0.915 ;
        RECT  1.000 0.355 1.085 0.915 ;
        RECT  0.145 0.355 1.000 0.425 ;
        RECT  0.225 0.845 1.000 0.915 ;
        RECT  0.035 0.215 0.145 0.425 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.345 0.640 ;
        RECT  1.855 0.495 1.925 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.785 0.640 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.093600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.495 0.930 0.640 ;
        RECT  0.580 0.495 0.685 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.095200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.450 0.640 ;
        RECT  0.150 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.115 2.520 0.115 ;
        RECT  2.365 -0.115 2.435 0.380 ;
        RECT  2.070 -0.115 2.365 0.115 ;
        RECT  1.940 -0.115 2.070 0.210 ;
        RECT  1.685 -0.115 1.940 0.115 ;
        RECT  1.555 -0.115 1.685 0.210 ;
        RECT  1.300 -0.115 1.555 0.115 ;
        RECT  1.180 -0.115 1.300 0.230 ;
        RECT  0.920 -0.115 1.180 0.115 ;
        RECT  0.800 -0.115 0.920 0.135 ;
        RECT  0.000 -0.115 0.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.445 1.145 2.520 1.375 ;
        RECT  2.365 0.720 2.445 1.375 ;
        RECT  2.065 1.145 2.365 1.375 ;
        RECT  1.945 1.050 2.065 1.375 ;
        RECT  0.000 1.145 1.945 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.370 0.845 2.265 0.915 ;
        RECT  0.125 0.995 1.690 1.065 ;
        RECT  0.220 0.205 1.110 0.275 ;
        RECT  0.055 0.915 0.125 1.065 ;
    END
END AOI211D3BWP40

MACRO AOI211D4BWP40
    CLASS CORE ;
    FOREIGN AOI211D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.627300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 0.190 3.280 0.415 ;
        RECT  2.870 0.345 3.160 0.415 ;
        RECT  2.750 0.190 2.870 0.415 ;
        RECT  2.480 0.345 2.750 0.415 ;
        RECT  2.360 0.190 2.480 0.415 ;
        RECT  2.100 0.345 2.360 0.415 ;
        RECT  1.980 0.190 2.100 0.415 ;
        RECT  0.735 0.345 1.980 0.415 ;
        RECT  1.595 0.700 1.705 0.915 ;
        RECT  0.735 0.845 1.595 0.915 ;
        RECT  0.525 0.345 0.735 0.915 ;
        RECT  0.220 0.345 0.525 0.415 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.495 3.250 0.625 ;
        RECT  2.695 0.495 2.765 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.455 0.625 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  0.885 0.495 1.295 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.765 ;
        RECT  0.035 0.495 0.315 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.460 ;
        RECT  3.060 -0.115 3.370 0.115 ;
        RECT  2.980 -0.115 3.060 0.275 ;
        RECT  2.650 -0.115 2.980 0.115 ;
        RECT  2.570 -0.115 2.650 0.275 ;
        RECT  2.270 -0.115 2.570 0.115 ;
        RECT  2.190 -0.115 2.270 0.275 ;
        RECT  1.890 -0.115 2.190 0.115 ;
        RECT  1.810 -0.115 1.890 0.275 ;
        RECT  1.510 -0.115 1.810 0.115 ;
        RECT  1.390 -0.115 1.510 0.130 ;
        RECT  1.110 -0.115 1.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.130 ;
        RECT  0.000 -0.115 0.990 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.145 3.500 1.375 ;
        RECT  3.180 0.860 3.260 1.375 ;
        RECT  2.850 1.145 3.180 1.375 ;
        RECT  2.770 1.005 2.850 1.375 ;
        RECT  0.000 1.145 2.770 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.160 0.190 3.280 0.415 ;
        RECT  2.870 0.345 3.160 0.415 ;
        RECT  2.750 0.190 2.870 0.415 ;
        RECT  2.480 0.345 2.750 0.415 ;
        RECT  2.360 0.190 2.480 0.415 ;
        RECT  2.100 0.345 2.360 0.415 ;
        RECT  1.980 0.190 2.100 0.415 ;
        RECT  0.805 0.345 1.980 0.415 ;
        RECT  1.595 0.700 1.705 0.915 ;
        RECT  0.805 0.845 1.595 0.915 ;
        RECT  0.220 0.345 0.455 0.415 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        RECT  3.370 0.720 3.450 1.010 ;
        RECT  3.060 0.720 3.370 0.790 ;
        RECT  2.980 0.720 3.060 1.010 ;
        RECT  1.905 0.855 2.980 0.925 ;
        RECT  0.220 0.995 2.480 1.065 ;
        RECT  1.795 0.715 1.905 0.925 ;
        RECT  0.130 0.205 1.710 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI211D4BWP40

MACRO AOI211D6BWP40
    CLASS CORE ;
    FOREIGN AOI211D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.923800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 0.190 4.820 0.415 ;
        RECT  4.410 0.345 4.700 0.415 ;
        RECT  4.290 0.190 4.410 0.415 ;
        RECT  4.010 0.345 4.290 0.415 ;
        RECT  3.890 0.190 4.010 0.415 ;
        RECT  3.630 0.345 3.890 0.415 ;
        RECT  3.510 0.190 3.630 0.415 ;
        RECT  3.250 0.345 3.510 0.415 ;
        RECT  3.130 0.190 3.250 0.415 ;
        RECT  2.870 0.345 3.130 0.415 ;
        RECT  2.750 0.190 2.870 0.415 ;
        RECT  0.735 0.345 2.750 0.415 ;
        RECT  2.365 0.650 2.475 0.915 ;
        RECT  2.075 0.845 2.365 0.915 ;
        RECT  1.965 0.705 2.075 0.915 ;
        RECT  1.675 0.845 1.965 0.915 ;
        RECT  1.565 0.705 1.675 0.915 ;
        RECT  0.735 0.845 1.565 0.915 ;
        RECT  0.525 0.345 0.735 0.915 ;
        RECT  0.220 0.345 0.525 0.415 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.495 4.725 0.765 ;
        RECT  3.840 0.495 4.655 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.495 3.700 0.625 ;
        RECT  2.835 0.495 2.905 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 2.205 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.191200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.765 ;
        RECT  0.035 0.495 0.315 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.460 ;
        RECT  4.600 -0.115 4.910 0.115 ;
        RECT  4.520 -0.115 4.600 0.275 ;
        RECT  4.190 -0.115 4.520 0.115 ;
        RECT  4.110 -0.115 4.190 0.275 ;
        RECT  3.800 -0.115 4.110 0.115 ;
        RECT  3.720 -0.115 3.800 0.275 ;
        RECT  3.420 -0.115 3.720 0.115 ;
        RECT  3.340 -0.115 3.420 0.275 ;
        RECT  3.040 -0.115 3.340 0.115 ;
        RECT  2.960 -0.115 3.040 0.275 ;
        RECT  2.660 -0.115 2.960 0.115 ;
        RECT  2.580 -0.115 2.660 0.275 ;
        RECT  2.280 -0.115 2.580 0.115 ;
        RECT  2.160 -0.115 2.280 0.130 ;
        RECT  1.880 -0.115 2.160 0.115 ;
        RECT  1.760 -0.115 1.880 0.130 ;
        RECT  1.495 -0.115 1.760 0.115 ;
        RECT  1.365 -0.115 1.495 0.130 ;
        RECT  0.000 -0.115 1.365 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.800 1.145 5.040 1.375 ;
        RECT  4.720 1.010 4.800 1.375 ;
        RECT  4.390 1.145 4.720 1.375 ;
        RECT  4.310 1.010 4.390 1.375 ;
        RECT  3.990 1.145 4.310 1.375 ;
        RECT  3.910 0.860 3.990 1.375 ;
        RECT  0.000 1.145 3.910 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.700 0.190 4.820 0.415 ;
        RECT  4.410 0.345 4.700 0.415 ;
        RECT  4.290 0.190 4.410 0.415 ;
        RECT  4.010 0.345 4.290 0.415 ;
        RECT  3.890 0.190 4.010 0.415 ;
        RECT  3.630 0.345 3.890 0.415 ;
        RECT  3.510 0.190 3.630 0.415 ;
        RECT  3.250 0.345 3.510 0.415 ;
        RECT  3.130 0.190 3.250 0.415 ;
        RECT  2.870 0.345 3.130 0.415 ;
        RECT  2.750 0.190 2.870 0.415 ;
        RECT  0.805 0.345 2.750 0.415 ;
        RECT  2.365 0.650 2.475 0.915 ;
        RECT  2.075 0.845 2.365 0.915 ;
        RECT  1.965 0.705 2.075 0.915 ;
        RECT  1.675 0.845 1.965 0.915 ;
        RECT  1.565 0.705 1.675 0.915 ;
        RECT  0.805 0.845 1.565 0.915 ;
        RECT  0.220 0.345 0.455 0.415 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        RECT  4.910 0.675 4.990 1.065 ;
        RECT  4.200 0.855 4.910 0.925 ;
        RECT  4.120 0.720 4.200 1.010 ;
        RECT  3.800 0.720 4.120 0.790 ;
        RECT  3.720 0.720 3.800 1.010 ;
        RECT  3.440 0.720 3.720 0.790 ;
        RECT  0.220 0.995 3.635 1.065 ;
        RECT  3.320 0.720 3.440 0.925 ;
        RECT  2.680 0.855 3.320 0.925 ;
        RECT  2.560 0.650 2.680 0.925 ;
        RECT  0.130 0.205 2.480 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI211D6BWP40

MACRO AOI211D8BWP40
    CLASS CORE ;
    FOREIGN AOI211D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.213300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.240 0.190 6.360 0.415 ;
        RECT  5.950 0.345 6.240 0.415 ;
        RECT  5.830 0.190 5.950 0.415 ;
        RECT  5.550 0.345 5.830 0.415 ;
        RECT  5.430 0.190 5.550 0.415 ;
        RECT  5.150 0.345 5.430 0.415 ;
        RECT  5.035 0.190 5.150 0.415 ;
        RECT  4.770 0.345 5.035 0.415 ;
        RECT  4.650 0.190 4.770 0.415 ;
        RECT  4.390 0.345 4.650 0.415 ;
        RECT  4.270 0.190 4.390 0.415 ;
        RECT  4.010 0.345 4.270 0.415 ;
        RECT  3.890 0.190 4.010 0.415 ;
        RECT  3.630 0.345 3.890 0.415 ;
        RECT  3.510 0.190 3.630 0.415 ;
        RECT  1.015 0.345 3.510 0.415 ;
        RECT  3.125 0.705 3.235 0.915 ;
        RECT  2.835 0.845 3.125 0.915 ;
        RECT  2.725 0.705 2.835 0.915 ;
        RECT  2.435 0.845 2.725 0.915 ;
        RECT  2.325 0.705 2.435 0.915 ;
        RECT  2.055 0.845 2.325 0.915 ;
        RECT  1.945 0.705 2.055 0.915 ;
        RECT  1.675 0.845 1.945 0.915 ;
        RECT  1.565 0.705 1.675 0.915 ;
        RECT  1.015 0.845 1.565 0.915 ;
        RECT  0.805 0.345 1.015 0.915 ;
        RECT  0.220 0.345 0.805 0.415 ;
        RECT  0.125 0.845 0.805 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.495 6.125 0.765 ;
        RECT  4.990 0.495 6.055 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.495 4.805 0.625 ;
        RECT  3.675 0.495 3.745 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.249600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.625 0.765 ;
        RECT  1.690 0.495 2.555 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.253600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.035 0.495 0.455 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 -0.115 6.580 0.115 ;
        RECT  6.450 -0.115 6.530 0.460 ;
        RECT  6.140 -0.115 6.450 0.115 ;
        RECT  6.060 -0.115 6.140 0.275 ;
        RECT  5.730 -0.115 6.060 0.115 ;
        RECT  5.650 -0.115 5.730 0.275 ;
        RECT  5.330 -0.115 5.650 0.115 ;
        RECT  5.250 -0.115 5.330 0.275 ;
        RECT  4.940 -0.115 5.250 0.115 ;
        RECT  4.860 -0.115 4.940 0.275 ;
        RECT  4.560 -0.115 4.860 0.115 ;
        RECT  4.480 -0.115 4.560 0.275 ;
        RECT  4.180 -0.115 4.480 0.115 ;
        RECT  4.100 -0.115 4.180 0.275 ;
        RECT  3.800 -0.115 4.100 0.115 ;
        RECT  3.720 -0.115 3.800 0.275 ;
        RECT  3.420 -0.115 3.720 0.115 ;
        RECT  3.340 -0.115 3.420 0.275 ;
        RECT  3.040 -0.115 3.340 0.115 ;
        RECT  2.920 -0.115 3.040 0.130 ;
        RECT  2.640 -0.115 2.920 0.115 ;
        RECT  2.520 -0.115 2.640 0.130 ;
        RECT  2.255 -0.115 2.520 0.115 ;
        RECT  2.125 -0.115 2.255 0.130 ;
        RECT  1.875 -0.115 2.125 0.115 ;
        RECT  1.745 -0.115 1.875 0.130 ;
        RECT  0.000 -0.115 1.745 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.340 1.145 6.580 1.375 ;
        RECT  6.260 1.000 6.340 1.375 ;
        RECT  5.930 1.145 6.260 1.375 ;
        RECT  5.850 1.000 5.930 1.375 ;
        RECT  5.530 1.145 5.850 1.375 ;
        RECT  5.450 0.860 5.530 1.375 ;
        RECT  5.130 1.145 5.450 1.375 ;
        RECT  5.050 0.860 5.130 1.375 ;
        RECT  0.000 1.145 5.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 0.190 6.360 0.415 ;
        RECT  5.950 0.345 6.240 0.415 ;
        RECT  5.830 0.190 5.950 0.415 ;
        RECT  5.550 0.345 5.830 0.415 ;
        RECT  5.430 0.190 5.550 0.415 ;
        RECT  5.150 0.345 5.430 0.415 ;
        RECT  5.035 0.190 5.150 0.415 ;
        RECT  4.770 0.345 5.035 0.415 ;
        RECT  4.650 0.190 4.770 0.415 ;
        RECT  4.390 0.345 4.650 0.415 ;
        RECT  4.270 0.190 4.390 0.415 ;
        RECT  4.010 0.345 4.270 0.415 ;
        RECT  3.890 0.190 4.010 0.415 ;
        RECT  3.630 0.345 3.890 0.415 ;
        RECT  3.510 0.190 3.630 0.415 ;
        RECT  1.085 0.345 3.510 0.415 ;
        RECT  3.125 0.705 3.235 0.915 ;
        RECT  2.835 0.845 3.125 0.915 ;
        RECT  2.725 0.705 2.835 0.915 ;
        RECT  2.435 0.845 2.725 0.915 ;
        RECT  2.325 0.705 2.435 0.915 ;
        RECT  2.055 0.845 2.325 0.915 ;
        RECT  1.945 0.705 2.055 0.915 ;
        RECT  1.675 0.845 1.945 0.915 ;
        RECT  1.565 0.705 1.675 0.915 ;
        RECT  1.085 0.845 1.565 0.915 ;
        RECT  0.220 0.345 0.735 0.415 ;
        RECT  0.125 0.845 0.735 0.915 ;
        RECT  0.055 0.845 0.125 1.070 ;
        RECT  6.450 0.675 6.530 1.065 ;
        RECT  5.730 0.850 6.450 0.920 ;
        RECT  5.650 0.720 5.730 1.010 ;
        RECT  5.340 0.720 5.650 0.790 ;
        RECT  5.260 0.720 5.340 1.010 ;
        RECT  4.940 0.720 5.260 0.790 ;
        RECT  4.860 0.720 4.940 1.010 ;
        RECT  4.585 0.720 4.860 0.790 ;
        RECT  0.220 0.995 4.780 1.065 ;
        RECT  4.455 0.720 4.585 0.925 ;
        RECT  4.205 0.720 4.455 0.790 ;
        RECT  4.080 0.720 4.205 0.925 ;
        RECT  3.440 0.855 4.080 0.925 ;
        RECT  3.320 0.720 3.440 0.925 ;
        RECT  0.130 0.205 3.240 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI211D8BWP40

MACRO AOI21D0BWP40
    CLASS CORE ;
    FOREIGN AOI21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.079300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.205 0.570 0.330 ;
        RECT  0.455 0.205 0.525 0.905 ;
        RECT  0.250 0.775 0.455 0.905 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.250 0.385 0.650 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.840 0.115 ;
        RECT  0.680 -0.115 0.760 0.250 ;
        RECT  0.130 -0.115 0.680 0.115 ;
        RECT  0.050 -0.115 0.130 0.260 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.840 1.375 ;
        RECT  0.680 1.005 0.760 1.375 ;
        RECT  0.000 1.145 0.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.590 1.055 ;
        RECT  0.055 0.885 0.125 1.055 ;
    END
END AOI21D0BWP40

MACRO AOI21D1BWP40
    CLASS CORE ;
    FOREIGN AOI21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.127000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.215 0.530 0.340 ;
        RECT  0.455 0.215 0.525 0.905 ;
        RECT  0.250 0.775 0.455 0.905 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.250 0.385 0.650 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.840 0.115 ;
        RECT  0.680 -0.115 0.760 0.410 ;
        RECT  0.130 -0.115 0.680 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.840 1.375 ;
        RECT  0.680 0.845 0.760 1.375 ;
        RECT  0.000 1.145 0.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.125 0.985 0.545 1.055 ;
        RECT  0.055 0.885 0.125 1.055 ;
    END
END AOI21D1BWP40

MACRO AOI21D2BWP40
    CLASS CORE ;
    FOREIGN AOI21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.301000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.195 1.365 0.415 ;
        RECT  0.525 0.345 1.240 0.415 ;
        RECT  0.610 0.845 1.100 0.915 ;
        RECT  0.530 0.710 0.610 0.915 ;
        RECT  0.410 0.710 0.530 0.780 ;
        RECT  0.415 0.195 0.525 0.415 ;
        RECT  0.410 0.345 0.415 0.415 ;
        RECT  0.315 0.345 0.410 0.780 ;
        RECT  0.145 0.345 0.315 0.415 ;
        RECT  0.035 0.195 0.145 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.495 1.085 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.365 0.625 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  0.750 0.695 1.155 0.765 ;
        RECT  0.680 0.495 0.750 0.765 ;
        RECT  0.550 0.495 0.680 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.915 -0.115 1.400 0.115 ;
        RECT  0.785 -0.115 0.915 0.240 ;
        RECT  0.340 -0.115 0.785 0.115 ;
        RECT  0.220 -0.115 0.340 0.240 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.310 1.145 1.400 1.375 ;
        RECT  0.240 1.010 0.310 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.270 0.915 1.340 1.055 ;
        RECT  0.460 0.985 1.270 1.055 ;
        RECT  0.380 0.860 0.460 1.055 ;
        RECT  0.125 0.860 0.380 0.930 ;
        RECT  0.055 0.860 0.125 1.015 ;
    END
END AOI21D2BWP40

MACRO AOI21D3BWP40
    CLASS CORE ;
    FOREIGN AOI21D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.345 1.680 0.420 ;
        RECT  1.295 0.345 1.365 0.815 ;
        RECT  0.785 0.345 1.295 0.420 ;
        RECT  1.095 0.735 1.295 0.815 ;
        RECT  0.990 0.735 1.095 0.915 ;
        RECT  0.215 0.845 0.990 0.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.845 0.625 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.135 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.495 1.155 0.650 ;
        RECT  0.735 0.495 0.840 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.115 1.960 0.115 ;
        RECT  1.800 -0.115 1.880 0.410 ;
        RECT  1.485 -0.115 1.800 0.115 ;
        RECT  1.360 -0.115 1.485 0.210 ;
        RECT  0.530 -0.115 1.360 0.115 ;
        RECT  0.410 -0.115 0.530 0.210 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.145 1.960 1.375 ;
        RECT  1.800 0.725 1.880 1.375 ;
        RECT  1.485 1.145 1.800 1.375 ;
        RECT  1.355 1.050 1.485 1.375 ;
        RECT  0.000 1.145 1.355 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.285 0.890 1.675 0.960 ;
        RECT  1.215 0.890 1.285 1.065 ;
        RECT  0.125 0.995 1.215 1.065 ;
        RECT  0.695 0.195 1.130 0.265 ;
        RECT  0.625 0.195 0.695 0.360 ;
        RECT  0.215 0.290 0.625 0.360 ;
        RECT  0.055 0.790 0.125 1.065 ;
    END
END AOI21D3BWP40

MACRO AOI21D4BWP40
    CLASS CORE ;
    FOREIGN AOI21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.516000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 0.200 2.420 0.410 ;
        RECT  2.035 0.340 2.300 0.410 ;
        RECT  1.925 0.195 2.035 0.410 ;
        RECT  1.855 0.340 1.925 0.410 ;
        RECT  1.785 0.340 1.855 0.765 ;
        RECT  1.520 0.695 1.785 0.765 ;
        RECT  1.450 0.695 1.520 0.915 ;
        RECT  0.735 0.845 1.450 0.915 ;
        RECT  0.525 0.350 0.735 0.915 ;
        RECT  0.220 0.350 0.525 0.420 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.315 0.625 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.440 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.435 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.470 ;
        RECT  2.210 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.210 0.270 ;
        RECT  1.840 -0.115 2.130 0.115 ;
        RECT  1.740 -0.115 1.840 0.270 ;
        RECT  1.460 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.460 0.265 ;
        RECT  1.075 -0.115 1.380 0.115 ;
        RECT  1.005 -0.115 1.075 0.265 ;
        RECT  0.000 -0.115 1.005 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.720 2.590 1.375 ;
        RECT  2.210 1.145 2.510 1.375 ;
        RECT  2.130 1.000 2.210 1.375 ;
        RECT  1.830 1.145 2.130 1.375 ;
        RECT  1.760 0.980 1.830 1.375 ;
        RECT  0.000 1.145 1.760 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.300 0.200 2.420 0.410 ;
        RECT  2.035 0.340 2.300 0.410 ;
        RECT  1.925 0.195 2.035 0.410 ;
        RECT  1.855 0.340 1.925 0.410 ;
        RECT  1.785 0.340 1.855 0.765 ;
        RECT  1.520 0.695 1.785 0.765 ;
        RECT  1.450 0.695 1.520 0.915 ;
        RECT  0.805 0.845 1.450 0.915 ;
        RECT  0.220 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        RECT  2.325 0.700 2.395 1.020 ;
        RECT  1.680 0.840 2.325 0.910 ;
        RECT  1.610 0.840 1.680 1.065 ;
        RECT  1.555 0.205 1.665 0.415 ;
        RECT  0.220 0.995 1.610 1.065 ;
        RECT  1.290 0.345 1.555 0.415 ;
        RECT  1.170 0.205 1.290 0.415 ;
        RECT  0.925 0.345 1.170 0.415 ;
        RECT  0.855 0.205 0.925 0.415 ;
        RECT  0.130 0.205 0.855 0.280 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI21D4BWP40

MACRO AOI21D6BWP40
    CLASS CORE ;
    FOREIGN AOI21D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.756000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.200 3.560 0.410 ;
        RECT  3.175 0.340 3.440 0.410 ;
        RECT  3.065 0.200 3.175 0.410 ;
        RECT  2.795 0.340 3.065 0.410 ;
        RECT  2.685 0.200 2.795 0.410 ;
        RECT  2.615 0.340 2.685 0.410 ;
        RECT  2.545 0.340 2.615 0.765 ;
        RECT  2.280 0.695 2.545 0.765 ;
        RECT  2.210 0.695 2.280 0.915 ;
        RECT  2.045 0.845 2.210 0.915 ;
        RECT  1.935 0.705 2.045 0.915 ;
        RECT  1.665 0.845 1.935 0.915 ;
        RECT  1.555 0.705 1.665 0.915 ;
        RECT  0.735 0.845 1.555 0.915 ;
        RECT  0.735 0.350 1.115 0.420 ;
        RECT  0.525 0.350 0.735 0.915 ;
        RECT  0.220 0.350 0.525 0.420 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.495 3.455 0.625 ;
        RECT  2.695 0.495 2.765 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 2.200 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.435 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.470 ;
        RECT  3.350 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.350 0.270 ;
        RECT  2.980 -0.115 3.270 0.115 ;
        RECT  2.880 -0.115 2.980 0.270 ;
        RECT  2.610 -0.115 2.880 0.115 ;
        RECT  2.500 -0.115 2.610 0.270 ;
        RECT  2.220 -0.115 2.500 0.115 ;
        RECT  2.140 -0.115 2.220 0.265 ;
        RECT  1.835 -0.115 2.140 0.115 ;
        RECT  1.765 -0.115 1.835 0.265 ;
        RECT  1.455 -0.115 1.765 0.115 ;
        RECT  1.385 -0.115 1.455 0.265 ;
        RECT  0.000 -0.115 1.385 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.720 3.730 1.375 ;
        RECT  3.350 1.145 3.650 1.375 ;
        RECT  3.270 0.840 3.350 1.375 ;
        RECT  2.970 1.145 3.270 1.375 ;
        RECT  2.900 0.980 2.970 1.375 ;
        RECT  2.585 1.145 2.900 1.375 ;
        RECT  2.515 0.980 2.585 1.375 ;
        RECT  0.000 1.145 2.515 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.440 0.200 3.560 0.410 ;
        RECT  3.175 0.340 3.440 0.410 ;
        RECT  3.065 0.200 3.175 0.410 ;
        RECT  2.795 0.340 3.065 0.410 ;
        RECT  2.685 0.200 2.795 0.410 ;
        RECT  2.615 0.340 2.685 0.410 ;
        RECT  2.545 0.340 2.615 0.765 ;
        RECT  2.280 0.695 2.545 0.765 ;
        RECT  2.210 0.695 2.280 0.915 ;
        RECT  2.045 0.845 2.210 0.915 ;
        RECT  1.935 0.705 2.045 0.915 ;
        RECT  1.665 0.845 1.935 0.915 ;
        RECT  1.555 0.705 1.665 0.915 ;
        RECT  0.805 0.845 1.555 0.915 ;
        RECT  0.805 0.350 1.115 0.420 ;
        RECT  0.220 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        RECT  3.465 0.700 3.535 1.020 ;
        RECT  3.155 0.700 3.465 0.770 ;
        RECT  3.085 0.700 3.155 1.020 ;
        RECT  2.435 0.840 3.085 0.910 ;
        RECT  2.365 0.840 2.435 1.065 ;
        RECT  2.315 0.205 2.425 0.415 ;
        RECT  0.220 0.995 2.365 1.065 ;
        RECT  2.050 0.345 2.315 0.415 ;
        RECT  1.930 0.205 2.050 0.415 ;
        RECT  1.670 0.345 1.930 0.415 ;
        RECT  1.550 0.205 1.670 0.415 ;
        RECT  1.305 0.345 1.550 0.415 ;
        RECT  1.235 0.205 1.305 0.415 ;
        RECT  0.130 0.205 1.235 0.280 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI21D6BWP40

MACRO AOI21D8BWP40
    CLASS CORE ;
    FOREIGN AOI21D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.011750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 0.200 4.820 0.410 ;
        RECT  4.440 0.340 4.700 0.410 ;
        RECT  4.320 0.200 4.440 0.410 ;
        RECT  4.060 0.340 4.320 0.410 ;
        RECT  3.940 0.200 4.060 0.410 ;
        RECT  3.650 0.340 3.940 0.410 ;
        RECT  3.530 0.200 3.650 0.410 ;
        RECT  3.380 0.340 3.530 0.410 ;
        RECT  3.310 0.340 3.380 0.765 ;
        RECT  3.040 0.695 3.310 0.765 ;
        RECT  2.970 0.695 3.040 0.915 ;
        RECT  2.805 0.845 2.970 0.915 ;
        RECT  2.695 0.700 2.805 0.915 ;
        RECT  2.425 0.845 2.695 0.915 ;
        RECT  2.315 0.700 2.425 0.915 ;
        RECT  2.045 0.845 2.315 0.915 ;
        RECT  1.935 0.700 2.045 0.915 ;
        RECT  1.285 0.845 1.935 0.915 ;
        RECT  0.875 0.350 1.505 0.420 ;
        RECT  1.175 0.700 1.285 0.915 ;
        RECT  0.875 0.845 1.175 0.915 ;
        RECT  0.665 0.350 0.875 0.915 ;
        RECT  0.220 0.350 0.665 0.420 ;
        RECT  0.125 0.845 0.665 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.495 4.715 0.625 ;
        RECT  3.675 0.495 3.745 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 2.960 0.625 ;
        RECT  1.715 0.495 1.785 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.435 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.470 ;
        RECT  4.610 -0.115 4.910 0.115 ;
        RECT  4.530 -0.115 4.610 0.270 ;
        RECT  4.230 -0.115 4.530 0.115 ;
        RECT  4.150 -0.115 4.230 0.270 ;
        RECT  3.850 -0.115 4.150 0.115 ;
        RECT  3.770 -0.115 3.850 0.270 ;
        RECT  3.430 -0.115 3.770 0.115 ;
        RECT  3.295 -0.115 3.430 0.270 ;
        RECT  2.980 -0.115 3.295 0.115 ;
        RECT  2.900 -0.115 2.980 0.265 ;
        RECT  2.595 -0.115 2.900 0.115 ;
        RECT  2.525 -0.115 2.595 0.265 ;
        RECT  2.215 -0.115 2.525 0.115 ;
        RECT  2.145 -0.115 2.215 0.265 ;
        RECT  1.835 -0.115 2.145 0.115 ;
        RECT  1.765 -0.115 1.835 0.265 ;
        RECT  0.000 -0.115 1.765 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.720 4.990 1.375 ;
        RECT  4.610 1.145 4.910 1.375 ;
        RECT  4.530 0.840 4.610 1.375 ;
        RECT  4.225 1.145 4.530 1.375 ;
        RECT  4.155 0.840 4.225 1.375 ;
        RECT  3.845 1.145 4.155 1.375 ;
        RECT  3.775 0.985 3.845 1.375 ;
        RECT  3.405 1.145 3.775 1.375 ;
        RECT  3.325 0.985 3.405 1.375 ;
        RECT  0.000 1.145 3.325 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.700 0.200 4.820 0.410 ;
        RECT  4.440 0.340 4.700 0.410 ;
        RECT  4.320 0.200 4.440 0.410 ;
        RECT  4.060 0.340 4.320 0.410 ;
        RECT  3.940 0.200 4.060 0.410 ;
        RECT  3.650 0.340 3.940 0.410 ;
        RECT  3.530 0.200 3.650 0.410 ;
        RECT  3.380 0.340 3.530 0.410 ;
        RECT  3.310 0.340 3.380 0.765 ;
        RECT  3.040 0.695 3.310 0.765 ;
        RECT  2.970 0.695 3.040 0.915 ;
        RECT  2.805 0.845 2.970 0.915 ;
        RECT  2.695 0.700 2.805 0.915 ;
        RECT  2.425 0.845 2.695 0.915 ;
        RECT  2.315 0.700 2.425 0.915 ;
        RECT  2.045 0.845 2.315 0.915 ;
        RECT  1.935 0.700 2.045 0.915 ;
        RECT  1.285 0.845 1.935 0.915 ;
        RECT  0.945 0.350 1.505 0.420 ;
        RECT  1.175 0.700 1.285 0.915 ;
        RECT  0.945 0.845 1.175 0.915 ;
        RECT  0.220 0.350 0.595 0.420 ;
        RECT  0.125 0.845 0.595 0.915 ;
        RECT  0.055 0.845 0.125 0.955 ;
        RECT  4.725 0.700 4.795 1.020 ;
        RECT  4.415 0.700 4.725 0.770 ;
        RECT  4.345 0.700 4.415 1.020 ;
        RECT  4.035 0.700 4.345 0.770 ;
        RECT  3.965 0.700 4.035 1.020 ;
        RECT  3.200 0.845 3.965 0.915 ;
        RECT  3.130 0.845 3.200 1.065 ;
        RECT  3.075 0.205 3.185 0.415 ;
        RECT  0.220 0.995 3.130 1.065 ;
        RECT  2.810 0.345 3.075 0.415 ;
        RECT  2.690 0.205 2.810 0.415 ;
        RECT  2.430 0.345 2.690 0.415 ;
        RECT  2.310 0.205 2.430 0.415 ;
        RECT  2.050 0.345 2.310 0.415 ;
        RECT  1.930 0.205 2.050 0.415 ;
        RECT  1.685 0.345 1.930 0.415 ;
        RECT  1.615 0.205 1.685 0.415 ;
        RECT  0.130 0.205 1.615 0.280 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI21D8BWP40

MACRO AOI221D0BWP40
    CLASS CORE ;
    FOREIGN AOI221D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.094000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.185 1.085 0.380 ;
        RECT  0.385 0.310 0.990 0.380 ;
        RECT  0.315 0.310 0.385 0.915 ;
        RECT  0.155 0.310 0.315 0.380 ;
        RECT  0.220 0.845 0.315 0.915 ;
        RECT  0.035 0.215 0.155 0.380 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.365 0.630 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.465 0.805 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.630 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.630 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.115 1.400 0.115 ;
        RECT  1.225 -0.115 1.305 0.280 ;
        RECT  0.705 -0.115 1.225 0.115 ;
        RECT  0.595 -0.115 0.705 0.240 ;
        RECT  0.525 -0.115 0.595 0.115 ;
        RECT  0.415 -0.115 0.525 0.240 ;
        RECT  0.000 -0.115 0.415 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.145 1.400 1.375 ;
        RECT  1.225 0.980 1.305 1.375 ;
        RECT  0.000 1.145 1.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.855 1.070 1.025 ;
        RECT  0.590 0.855 0.990 0.925 ;
        RECT  0.125 0.995 0.900 1.065 ;
        RECT  0.055 0.895 0.125 1.065 ;
    END
END AOI221D0BWP40

MACRO AOI221D1BWP40
    CLASS CORE ;
    FOREIGN AOI221D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.167250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.975 0.195 1.085 0.415 ;
        RECT  0.385 0.345 0.975 0.415 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.145 0.345 0.315 0.415 ;
        RECT  0.220 0.845 0.315 0.915 ;
        RECT  0.035 0.195 0.145 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.295 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.695 0.855 0.765 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.875 0.495 1.015 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.115 1.400 0.115 ;
        RECT  1.225 -0.115 1.305 0.400 ;
        RECT  0.685 -0.115 1.225 0.115 ;
        RECT  0.615 -0.115 0.685 0.260 ;
        RECT  0.505 -0.115 0.615 0.115 ;
        RECT  0.435 -0.115 0.505 0.260 ;
        RECT  0.000 -0.115 0.435 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.145 1.400 1.375 ;
        RECT  1.225 0.880 1.305 1.375 ;
        RECT  0.000 1.145 1.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.590 0.845 1.090 0.915 ;
        RECT  0.125 0.985 0.900 1.055 ;
        RECT  0.055 0.895 0.125 1.055 ;
    END
END AOI221D1BWP40

MACRO AOI221D2BWP40
    CLASS CORE ;
    FOREIGN AOI221D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.377500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.195 2.120 0.415 ;
        RECT  0.925 0.345 1.995 0.415 ;
        RECT  0.130 0.845 0.930 0.915 ;
        RECT  0.815 0.190 0.925 0.415 ;
        RECT  0.145 0.345 0.815 0.415 ;
        RECT  0.105 0.190 0.145 0.415 ;
        RECT  0.105 0.845 0.130 1.045 ;
        RECT  0.035 0.190 0.105 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.345 0.645 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.835 0.775 ;
        RECT  1.240 0.705 1.715 0.775 ;
        RECT  1.165 0.495 1.240 0.775 ;
        RECT  1.100 0.495 1.165 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.645 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.695 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.765 0.495 0.845 0.775 ;
        RECT  0.255 0.705 0.765 0.775 ;
        RECT  0.175 0.495 0.255 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 -0.115 2.380 0.115 ;
        RECT  2.235 -0.115 2.315 0.400 ;
        RECT  1.845 -0.115 2.235 0.115 ;
        RECT  1.775 -0.115 1.845 0.265 ;
        RECT  1.110 -0.115 1.775 0.115 ;
        RECT  0.995 -0.115 1.110 0.275 ;
        RECT  0.550 -0.115 0.995 0.115 ;
        RECT  0.430 -0.115 0.550 0.220 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.105 1.145 2.380 1.375 ;
        RECT  2.025 1.000 2.105 1.375 ;
        RECT  0.000 1.145 2.025 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.220 0.845 2.330 1.065 ;
        RECT  1.865 0.845 2.220 0.915 ;
        RECT  1.755 0.845 1.865 1.065 ;
        RECT  1.085 0.845 1.755 0.915 ;
        RECT  1.180 0.195 1.680 0.265 ;
        RECT  0.220 0.985 1.675 1.055 ;
        RECT  1.015 0.775 1.085 0.915 ;
    END
END AOI221D2BWP40

MACRO AOI221D4BWP40
    CLASS CORE ;
    FOREIGN AOI221D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.640700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 3.970 0.425 ;
        RECT  1.575 0.845 1.670 0.915 ;
        RECT  1.365 0.355 1.575 0.915 ;
        RECT  0.145 0.355 1.365 0.425 ;
        RECT  0.130 0.845 1.365 0.915 ;
        RECT  0.035 0.215 0.145 0.425 ;
        RECT  0.035 0.845 0.130 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 4.165 0.645 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.220 0.495 3.340 0.775 ;
        RECT  2.135 0.705 3.220 0.775 ;
        RECT  2.060 0.535 2.135 0.775 ;
        RECT  1.995 0.535 2.060 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.465 0.495 3.060 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.365 0.495 0.960 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.775 ;
        RECT  0.255 0.705 1.155 0.775 ;
        RECT  0.175 0.495 0.255 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 -0.115 4.200 0.115 ;
        RECT  4.060 -0.115 4.140 0.400 ;
        RECT  3.760 -0.115 4.060 0.115 ;
        RECT  3.680 -0.115 3.760 0.280 ;
        RECT  3.355 -0.115 3.680 0.115 ;
        RECT  3.275 -0.115 3.355 0.280 ;
        RECT  2.235 -0.115 3.275 0.115 ;
        RECT  2.105 -0.115 2.235 0.140 ;
        RECT  1.845 -0.115 2.105 0.115 ;
        RECT  1.730 -0.115 1.845 0.275 ;
        RECT  0.910 -0.115 1.730 0.115 ;
        RECT  0.790 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.145 4.200 1.375 ;
        RECT  3.870 1.000 3.950 1.375 ;
        RECT  3.570 1.145 3.870 1.375 ;
        RECT  3.490 1.000 3.570 1.375 ;
        RECT  0.000 1.145 3.490 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.355 3.970 0.425 ;
        RECT  1.645 0.845 1.670 0.915 ;
        RECT  0.145 0.355 1.295 0.425 ;
        RECT  0.130 0.845 1.295 0.915 ;
        RECT  0.035 0.215 0.145 0.425 ;
        RECT  0.035 0.845 0.130 1.045 ;
        RECT  4.045 0.845 4.155 1.065 ;
        RECT  3.775 0.845 4.045 0.915 ;
        RECT  3.665 0.845 3.775 1.065 ;
        RECT  1.825 0.845 3.665 0.915 ;
        RECT  1.925 0.215 3.195 0.285 ;
        RECT  0.220 0.985 3.185 1.055 ;
        RECT  1.755 0.775 1.825 0.915 ;
        RECT  0.225 0.215 1.505 0.285 ;
    END
END AOI221D4BWP40

MACRO AOI222D0BWP40
    CLASS CORE ;
    FOREIGN AOI222D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.089625 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.195 1.110 0.390 ;
        RECT  0.525 0.320 1.030 0.390 ;
        RECT  0.455 0.210 0.525 0.915 ;
        RECT  0.220 0.845 0.455 0.915 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.505 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.695 0.730 0.765 ;
        RECT  0.595 0.470 0.665 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.315 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.300 ;
        RECT  0.950 -0.115 1.400 0.115 ;
        RECT  0.830 -0.115 0.950 0.250 ;
        RECT  0.140 -0.115 0.830 0.115 ;
        RECT  0.040 -0.115 0.140 0.300 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.965 1.500 1.375 ;
        RECT  1.120 1.145 1.400 1.375 ;
        RECT  1.020 0.985 1.120 1.375 ;
        RECT  0.000 1.145 1.020 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.845 1.320 1.055 ;
        RECT  0.620 0.845 1.200 0.915 ;
        RECT  0.130 0.995 0.945 1.065 ;
        RECT  0.050 0.910 0.130 1.065 ;
    END
END AOI222D0BWP40

MACRO AOI222D1BWP40
    CLASS CORE ;
    FOREIGN AOI222D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.167250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.185 1.130 0.390 ;
        RECT  0.525 0.320 1.010 0.390 ;
        RECT  0.455 0.195 0.525 0.915 ;
        RECT  0.220 0.845 0.455 0.915 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.505 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.695 0.710 0.765 ;
        RECT  0.595 0.470 0.665 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.315 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.420 ;
        RECT  0.940 -0.115 1.400 0.115 ;
        RECT  0.840 -0.115 0.940 0.250 ;
        RECT  0.140 -0.115 0.840 0.115 ;
        RECT  0.040 -0.115 0.140 0.425 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.870 1.500 1.375 ;
        RECT  1.120 1.145 1.400 1.375 ;
        RECT  1.020 0.985 1.120 1.375 ;
        RECT  0.000 1.145 1.020 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.845 1.320 1.055 ;
        RECT  0.620 0.845 1.200 0.915 ;
        RECT  0.130 0.995 0.945 1.065 ;
        RECT  0.050 0.865 0.130 1.065 ;
    END
END AOI222D1BWP40

MACRO AOI222D2BWP40
    CLASS CORE ;
    FOREIGN AOI222D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.356500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.345 2.230 0.415 ;
        RECT  0.905 0.345 0.945 0.775 ;
        RECT  0.890 0.205 0.905 0.775 ;
        RECT  0.875 0.205 0.890 0.915 ;
        RECT  0.735 0.205 0.875 0.415 ;
        RECT  0.810 0.705 0.875 0.915 ;
        RECT  0.145 0.845 0.810 0.915 ;
        RECT  0.145 0.345 0.735 0.415 ;
        RECT  0.035 0.205 0.145 0.415 ;
        RECT  0.035 0.845 0.145 1.055 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.455 0.495 2.625 0.625 ;
        RECT  2.385 0.495 2.455 0.775 ;
        RECT  1.925 0.705 2.385 0.775 ;
        RECT  1.845 0.495 1.925 0.775 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.235 0.630 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.705 0.775 ;
        RECT  1.155 0.705 1.575 0.775 ;
        RECT  1.085 0.495 1.155 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.495 1.505 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.740 0.495 0.805 0.615 ;
        RECT  0.670 0.495 0.740 0.775 ;
        RECT  0.245 0.705 0.670 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.420 ;
        RECT  1.825 -0.115 2.510 0.115 ;
        RECT  1.755 -0.115 1.825 0.275 ;
        RECT  1.090 -0.115 1.755 0.115 ;
        RECT  0.975 -0.115 1.090 0.275 ;
        RECT  0.530 -0.115 0.975 0.115 ;
        RECT  0.410 -0.115 0.530 0.220 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 1.145 2.660 1.375 ;
        RECT  2.320 0.985 2.400 1.375 ;
        RECT  2.020 1.145 2.320 1.375 ;
        RECT  1.940 0.985 2.020 1.375 ;
        RECT  0.000 1.145 1.940 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.495 0.845 2.605 1.055 ;
        RECT  2.230 0.845 2.495 0.915 ;
        RECT  1.920 0.195 2.420 0.265 ;
        RECT  2.110 0.845 2.230 1.055 ;
        RECT  1.840 0.845 2.110 0.915 ;
        RECT  1.740 0.845 1.840 1.070 ;
        RECT  0.970 0.845 1.740 0.915 ;
        RECT  1.160 0.195 1.660 0.265 ;
        RECT  0.225 0.995 1.660 1.065 ;
    END
END AOI222D2BWP40

MACRO AOI222D4BWP40
    CLASS CORE ;
    FOREIGN AOI222D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.642350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 4.610 0.415 ;
        RECT  1.575 0.785 1.650 0.915 ;
        RECT  1.365 0.345 1.575 0.915 ;
        RECT  0.145 0.345 1.365 0.415 ;
        RECT  0.145 0.845 1.365 0.915 ;
        RECT  0.035 0.205 0.145 0.415 ;
        RECT  0.035 0.845 0.145 1.055 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.765 0.495 4.890 0.775 ;
        RECT  3.620 0.705 4.765 0.775 ;
        RECT  3.530 0.495 3.620 0.775 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.495 4.625 0.630 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.250 0.775 ;
        RECT  2.090 0.705 3.115 0.775 ;
        RECT  1.975 0.495 2.090 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.495 3.045 0.630 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.895 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.545 1.235 0.615 ;
        RECT  1.015 0.545 1.130 0.775 ;
        RECT  0.245 0.705 1.015 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 -0.115 5.040 0.115 ;
        RECT  4.890 -0.115 4.970 0.420 ;
        RECT  3.750 -0.115 4.890 0.115 ;
        RECT  3.625 -0.115 3.750 0.135 ;
        RECT  3.345 -0.115 3.625 0.115 ;
        RECT  3.275 -0.115 3.345 0.275 ;
        RECT  2.235 -0.115 3.275 0.115 ;
        RECT  2.105 -0.115 2.235 0.135 ;
        RECT  1.845 -0.115 2.105 0.115 ;
        RECT  1.730 -0.115 1.845 0.275 ;
        RECT  0.915 -0.115 1.730 0.115 ;
        RECT  0.785 -0.115 0.915 0.135 ;
        RECT  0.530 -0.115 0.785 0.115 ;
        RECT  0.410 -0.115 0.530 0.135 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.780 1.145 5.040 1.375 ;
        RECT  4.700 0.985 4.780 1.375 ;
        RECT  4.400 1.145 4.700 1.375 ;
        RECT  4.320 0.985 4.400 1.375 ;
        RECT  3.960 1.145 4.320 1.375 ;
        RECT  3.870 0.985 3.960 1.375 ;
        RECT  3.560 1.145 3.870 1.375 ;
        RECT  3.445 0.985 3.560 1.375 ;
        RECT  0.000 1.145 3.445 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.345 4.610 0.415 ;
        RECT  1.645 0.785 1.650 0.915 ;
        RECT  0.145 0.345 1.295 0.415 ;
        RECT  0.145 0.845 1.295 0.915 ;
        RECT  0.035 0.205 0.145 0.415 ;
        RECT  0.035 0.845 0.145 1.055 ;
        RECT  4.875 0.845 4.985 1.055 ;
        RECT  4.610 0.845 4.875 0.915 ;
        RECT  3.440 0.205 4.800 0.275 ;
        RECT  4.490 0.845 4.610 1.055 ;
        RECT  4.175 0.845 4.490 0.915 ;
        RECT  4.070 0.845 4.175 1.070 ;
        RECT  3.740 0.845 4.070 0.915 ;
        RECT  3.635 0.845 3.740 1.070 ;
        RECT  3.360 0.845 3.635 0.915 ;
        RECT  3.260 0.845 3.360 1.070 ;
        RECT  1.730 0.845 3.260 0.915 ;
        RECT  1.925 0.205 3.180 0.275 ;
        RECT  0.225 0.995 3.180 1.065 ;
        RECT  0.225 0.205 1.495 0.275 ;
    END
END AOI222D4BWP40

MACRO AOI22D0BWP40
    CLASS CORE ;
    FOREIGN AOI22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.073000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.720 0.805 0.915 ;
        RECT  0.525 0.720 0.645 0.790 ;
        RECT  0.455 0.195 0.525 0.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.330 0.385 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.640 ;
        RECT  0.780 0.520 0.875 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.695 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.265 ;
        RECT  0.130 -0.115 0.850 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.980 1.375 ;
        RECT  0.240 1.045 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 0.995 0.945 1.065 ;
        RECT  0.460 0.905 0.540 1.065 ;
        RECT  0.130 0.905 0.460 0.975 ;
        RECT  0.050 0.905 0.130 1.045 ;
    END
END AOI22D0BWP40

MACRO AOI22D1BWP40
    CLASS CORE ;
    FOREIGN AOI22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.134000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.720 0.760 0.790 ;
        RECT  0.455 0.195 0.525 0.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.330 0.385 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.640 ;
        RECT  0.780 0.520 0.875 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.695 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.265 ;
        RECT  0.130 -0.115 0.850 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.145 0.980 1.375 ;
        RECT  0.240 1.015 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.835 0.865 0.945 1.075 ;
        RECT  0.555 0.865 0.835 0.935 ;
        RECT  0.445 0.865 0.555 1.075 ;
        RECT  0.145 0.865 0.445 0.935 ;
        RECT  0.035 0.865 0.145 1.075 ;
    END
END AOI22D1BWP40

MACRO AOI22D2BWP40
    CLASS CORE ;
    FOREIGN AOI22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.289200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.205 1.785 0.915 ;
        RECT  0.130 0.205 1.715 0.275 ;
        RECT  1.015 0.845 1.715 0.915 ;
        RECT  0.035 0.205 0.130 0.345 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.495 0.805 0.775 ;
        RECT  0.245 0.705 0.700 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.505 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.775 ;
        RECT  1.085 0.705 1.575 0.775 ;
        RECT  0.950 0.495 1.085 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.820 0.115 ;
        RECT  1.200 -0.115 1.320 0.135 ;
        RECT  0.540 -0.115 1.200 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 1.820 1.375 ;
        RECT  0.620 0.985 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.935 0.985 1.760 1.055 ;
        RECT  1.000 0.345 1.530 0.415 ;
        RECT  0.825 0.845 0.935 1.055 ;
        RECT  0.535 0.845 0.825 0.915 ;
        RECT  0.220 0.345 0.750 0.415 ;
        RECT  0.425 0.845 0.535 1.065 ;
        RECT  0.145 0.845 0.425 0.915 ;
        RECT  0.035 0.845 0.145 1.065 ;
    END
END AOI22D2BWP40

MACRO AOI22D3BWP40
    CLASS CORE ;
    FOREIGN AOI22D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.383000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.720 2.345 0.790 ;
        RECT  1.225 0.345 1.720 0.415 ;
        RECT  1.155 0.345 1.225 0.790 ;
        RECT  0.795 0.345 1.155 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.525 0.645 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.715 0.495 0.875 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 0.495 2.485 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.785 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.400 ;
        RECT  2.085 -0.115 2.390 0.115 ;
        RECT  2.015 -0.115 2.085 0.260 ;
        RECT  0.530 -0.115 2.015 0.115 ;
        RECT  0.410 -0.115 0.530 0.220 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.145 2.520 1.375 ;
        RECT  0.980 1.015 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 1.015 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 1.015 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.375 0.865 2.485 1.075 ;
        RECT  2.105 0.865 2.375 0.935 ;
        RECT  2.185 0.195 2.295 0.410 ;
        RECT  1.915 0.340 2.185 0.410 ;
        RECT  1.995 0.865 2.105 1.075 ;
        RECT  1.705 0.865 1.995 0.935 ;
        RECT  1.805 0.195 1.915 0.410 ;
        RECT  1.405 0.195 1.805 0.265 ;
        RECT  1.595 0.865 1.705 1.075 ;
        RECT  1.315 0.865 1.595 0.935 ;
        RECT  1.205 0.865 1.315 1.075 ;
        RECT  0.905 0.865 1.205 0.935 ;
        RECT  0.715 0.195 1.115 0.265 ;
        RECT  0.795 0.865 0.905 1.075 ;
        RECT  0.525 0.865 0.795 0.935 ;
        RECT  0.605 0.195 0.715 0.415 ;
        RECT  0.335 0.345 0.605 0.415 ;
        RECT  0.415 0.865 0.525 1.075 ;
        RECT  0.145 0.865 0.415 0.935 ;
        RECT  0.225 0.195 0.335 0.415 ;
        RECT  0.035 0.865 0.145 1.075 ;
    END
END AOI22D3BWP40

MACRO AOI22D4BWP40
    CLASS CORE ;
    FOREIGN AOI22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.515300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 0.355 3.270 0.425 ;
        RECT  2.570 0.355 2.640 0.775 ;
        RECT  1.265 0.705 2.570 0.775 ;
        RECT  1.195 0.705 1.265 0.905 ;
        RECT  0.735 0.775 1.195 0.905 ;
        RECT  0.525 0.350 0.735 0.905 ;
        RECT  0.220 0.350 0.525 0.420 ;
        RECT  0.125 0.775 0.525 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.435 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.805 0.495 3.315 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.435 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.445 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 -0.115 3.500 0.115 ;
        RECT  2.330 -0.115 2.450 0.145 ;
        RECT  2.030 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.030 0.275 ;
        RECT  1.460 -0.115 1.950 0.115 ;
        RECT  1.380 -0.115 1.460 0.265 ;
        RECT  1.080 -0.115 1.380 0.115 ;
        RECT  1.000 -0.115 1.080 0.265 ;
        RECT  0.000 -0.115 1.000 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.720 3.450 1.375 ;
        RECT  3.040 1.145 3.370 1.375 ;
        RECT  2.960 0.860 3.040 1.375 ;
        RECT  2.640 1.145 2.960 1.375 ;
        RECT  2.560 0.990 2.640 1.375 ;
        RECT  2.220 1.145 2.560 1.375 ;
        RECT  2.140 0.990 2.220 1.375 ;
        RECT  1.840 1.145 2.140 1.375 ;
        RECT  1.740 0.990 1.840 1.375 ;
        RECT  0.000 1.145 1.740 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.640 0.355 3.270 0.425 ;
        RECT  2.570 0.355 2.640 0.775 ;
        RECT  1.265 0.705 2.570 0.775 ;
        RECT  1.195 0.705 1.265 0.905 ;
        RECT  0.805 0.775 1.195 0.905 ;
        RECT  0.220 0.350 0.455 0.420 ;
        RECT  0.125 0.775 0.455 0.905 ;
        RECT  0.055 0.775 0.125 1.065 ;
        RECT  3.370 0.215 3.450 0.375 ;
        RECT  2.250 0.215 3.370 0.285 ;
        RECT  3.175 0.710 3.245 1.000 ;
        RECT  2.835 0.710 3.175 0.790 ;
        RECT  2.765 0.710 2.835 1.025 ;
        RECT  2.450 0.850 2.765 0.920 ;
        RECT  2.330 0.850 2.450 1.060 ;
        RECT  2.040 0.850 2.330 0.920 ;
        RECT  2.130 0.215 2.250 0.415 ;
        RECT  1.850 0.345 2.130 0.415 ;
        RECT  1.920 0.850 2.040 1.060 ;
        RECT  1.455 0.850 1.920 0.920 ;
        RECT  1.735 0.205 1.850 0.415 ;
        RECT  1.550 0.205 1.665 0.415 ;
        RECT  1.290 0.345 1.550 0.415 ;
        RECT  1.385 0.850 1.455 1.045 ;
        RECT  0.220 0.975 1.385 1.045 ;
        RECT  1.170 0.205 1.290 0.415 ;
        RECT  0.920 0.345 1.170 0.415 ;
        RECT  0.850 0.210 0.920 0.415 ;
        RECT  0.130 0.210 0.850 0.280 ;
        RECT  0.050 0.210 0.130 0.370 ;
    END
END AOI22D4BWP40

MACRO AOI22D6BWP40
    CLASS CORE ;
    FOREIGN AOI22D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.761550 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.790 0.355 4.810 0.425 ;
        RECT  3.720 0.355 3.790 0.775 ;
        RECT  2.030 0.705 3.720 0.775 ;
        RECT  1.960 0.705 2.030 0.915 ;
        RECT  0.735 0.845 1.960 0.915 ;
        RECT  0.735 0.350 1.095 0.420 ;
        RECT  0.525 0.350 0.735 0.915 ;
        RECT  0.220 0.350 0.525 0.420 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 1.010 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.605 0.625 ;
        RECT  2.690 0.495 3.535 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.189600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.025 0.495 4.855 0.625 ;
        RECT  3.955 0.495 4.025 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 2.200 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.610 -0.115 5.040 0.115 ;
        RECT  3.480 -0.115 3.610 0.145 ;
        RECT  3.215 -0.115 3.480 0.115 ;
        RECT  3.095 -0.115 3.215 0.145 ;
        RECT  2.795 -0.115 3.095 0.115 ;
        RECT  2.715 -0.115 2.795 0.275 ;
        RECT  2.225 -0.115 2.715 0.115 ;
        RECT  2.145 -0.115 2.225 0.265 ;
        RECT  1.855 -0.115 2.145 0.115 ;
        RECT  1.775 -0.115 1.855 0.265 ;
        RECT  1.485 -0.115 1.775 0.115 ;
        RECT  1.390 -0.115 1.485 0.265 ;
        RECT  0.000 -0.115 1.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.720 4.990 1.375 ;
        RECT  4.580 1.145 4.910 1.375 ;
        RECT  4.500 0.860 4.580 1.375 ;
        RECT  4.190 1.145 4.500 1.375 ;
        RECT  4.110 0.990 4.190 1.375 ;
        RECT  3.775 1.145 4.110 1.375 ;
        RECT  3.695 0.990 3.775 1.375 ;
        RECT  3.395 1.145 3.695 1.375 ;
        RECT  3.315 0.990 3.395 1.375 ;
        RECT  2.985 1.145 3.315 1.375 ;
        RECT  2.905 0.990 2.985 1.375 ;
        RECT  2.605 1.145 2.905 1.375 ;
        RECT  2.505 0.990 2.605 1.375 ;
        RECT  0.000 1.145 2.505 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.790 0.355 4.810 0.425 ;
        RECT  3.720 0.355 3.790 0.775 ;
        RECT  2.030 0.705 3.720 0.775 ;
        RECT  1.960 0.705 2.030 0.915 ;
        RECT  0.805 0.845 1.960 0.915 ;
        RECT  0.805 0.350 1.095 0.420 ;
        RECT  0.220 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 1.010 ;
        RECT  4.895 0.215 5.005 0.425 ;
        RECT  3.415 0.215 4.895 0.285 ;
        RECT  4.715 0.710 4.785 1.000 ;
        RECT  4.375 0.710 4.715 0.790 ;
        RECT  4.305 0.710 4.375 1.025 ;
        RECT  4.025 0.850 4.305 0.920 ;
        RECT  3.900 0.850 4.025 1.060 ;
        RECT  3.605 0.850 3.900 0.920 ;
        RECT  3.485 0.850 3.605 1.060 ;
        RECT  3.215 0.850 3.485 0.920 ;
        RECT  3.295 0.215 3.415 0.415 ;
        RECT  3.015 0.345 3.295 0.415 ;
        RECT  3.095 0.850 3.215 1.060 ;
        RECT  2.805 0.850 3.095 0.920 ;
        RECT  2.895 0.215 3.015 0.415 ;
        RECT  2.615 0.345 2.895 0.415 ;
        RECT  2.685 0.850 2.805 1.060 ;
        RECT  2.220 0.850 2.685 0.920 ;
        RECT  2.500 0.205 2.615 0.415 ;
        RECT  2.315 0.205 2.430 0.415 ;
        RECT  2.055 0.345 2.315 0.415 ;
        RECT  2.150 0.850 2.220 1.065 ;
        RECT  0.220 0.995 2.150 1.065 ;
        RECT  1.935 0.205 2.055 0.415 ;
        RECT  1.675 0.345 1.935 0.415 ;
        RECT  1.555 0.205 1.675 0.415 ;
        RECT  1.290 0.345 1.555 0.415 ;
        RECT  1.175 0.210 1.290 0.415 ;
        RECT  0.130 0.210 1.175 0.280 ;
        RECT  0.050 0.210 0.130 0.370 ;
    END
END AOI22D6BWP40

MACRO AOI22D8BWP40
    CLASS CORE ;
    FOREIGN AOI22D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.002300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.925 0.355 6.350 0.425 ;
        RECT  4.855 0.355 4.925 0.775 ;
        RECT  2.805 0.705 4.855 0.775 ;
        RECT  2.695 0.705 2.805 0.915 ;
        RECT  2.425 0.845 2.695 0.915 ;
        RECT  2.315 0.705 2.425 0.915 ;
        RECT  2.045 0.845 2.315 0.915 ;
        RECT  1.935 0.705 2.045 0.915 ;
        RECT  1.285 0.845 1.935 0.915 ;
        RECT  0.875 0.350 1.490 0.420 ;
        RECT  1.175 0.705 1.285 0.915 ;
        RECT  0.875 0.845 1.175 0.915 ;
        RECT  0.665 0.350 0.875 0.915 ;
        RECT  0.220 0.350 0.665 0.420 ;
        RECT  0.125 0.845 0.665 0.915 ;
        RECT  0.055 0.845 0.125 1.015 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.249600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.355 4.725 0.625 ;
        RECT  3.445 0.495 4.655 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.255200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.145 0.495 6.395 0.625 ;
        RECT  5.075 0.495 5.145 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 2.955 0.625 ;
        RECT  1.715 0.495 1.785 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.740 -0.115 6.580 0.115 ;
        RECT  4.620 -0.115 4.740 0.145 ;
        RECT  4.365 -0.115 4.620 0.115 ;
        RECT  4.235 -0.115 4.365 0.145 ;
        RECT  3.970 -0.115 4.235 0.115 ;
        RECT  3.850 -0.115 3.970 0.145 ;
        RECT  3.550 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.550 0.275 ;
        RECT  2.980 -0.115 3.470 0.115 ;
        RECT  2.900 -0.115 2.980 0.265 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.520 -0.115 2.600 0.265 ;
        RECT  2.220 -0.115 2.520 0.115 ;
        RECT  2.145 -0.115 2.220 0.265 ;
        RECT  1.840 -0.115 2.145 0.115 ;
        RECT  1.760 -0.115 1.840 0.265 ;
        RECT  0.000 -0.115 1.760 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.580 1.375 ;
        RECT  6.450 0.720 6.530 1.375 ;
        RECT  6.120 1.145 6.450 1.375 ;
        RECT  6.040 0.860 6.120 1.375 ;
        RECT  5.730 1.145 6.040 1.375 ;
        RECT  5.650 0.860 5.730 1.375 ;
        RECT  5.350 1.145 5.650 1.375 ;
        RECT  5.270 0.990 5.350 1.375 ;
        RECT  4.910 1.145 5.270 1.375 ;
        RECT  4.830 0.990 4.910 1.375 ;
        RECT  4.530 1.145 4.830 1.375 ;
        RECT  4.450 0.990 4.530 1.375 ;
        RECT  4.150 1.145 4.450 1.375 ;
        RECT  4.070 0.990 4.150 1.375 ;
        RECT  3.740 1.145 4.070 1.375 ;
        RECT  3.660 0.990 3.740 1.375 ;
        RECT  3.360 1.145 3.660 1.375 ;
        RECT  3.260 0.990 3.360 1.375 ;
        RECT  0.000 1.145 3.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.925 0.355 6.350 0.425 ;
        RECT  4.855 0.355 4.925 0.775 ;
        RECT  2.805 0.705 4.855 0.775 ;
        RECT  2.695 0.705 2.805 0.915 ;
        RECT  2.425 0.845 2.695 0.915 ;
        RECT  2.315 0.705 2.425 0.915 ;
        RECT  2.045 0.845 2.315 0.915 ;
        RECT  1.935 0.705 2.045 0.915 ;
        RECT  1.285 0.845 1.935 0.915 ;
        RECT  0.945 0.350 1.490 0.420 ;
        RECT  1.175 0.705 1.285 0.915 ;
        RECT  0.945 0.845 1.175 0.915 ;
        RECT  0.220 0.350 0.595 0.420 ;
        RECT  0.125 0.845 0.595 0.915 ;
        RECT  0.055 0.845 0.125 1.015 ;
        RECT  6.435 0.215 6.545 0.425 ;
        RECT  4.550 0.215 6.435 0.285 ;
        RECT  6.255 0.710 6.325 1.000 ;
        RECT  5.915 0.710 6.255 0.790 ;
        RECT  5.845 0.710 5.915 1.025 ;
        RECT  5.540 0.710 5.845 0.780 ;
        RECT  5.460 0.710 5.540 1.025 ;
        RECT  5.180 0.850 5.460 0.920 ;
        RECT  5.060 0.850 5.180 1.060 ;
        RECT  4.740 0.850 5.060 0.920 ;
        RECT  4.620 0.850 4.740 1.060 ;
        RECT  4.360 0.850 4.620 0.920 ;
        RECT  4.430 0.215 4.550 0.415 ;
        RECT  4.170 0.345 4.430 0.415 ;
        RECT  4.240 0.850 4.360 1.060 ;
        RECT  3.970 0.850 4.240 0.920 ;
        RECT  4.050 0.215 4.170 0.415 ;
        RECT  3.770 0.345 4.050 0.415 ;
        RECT  3.850 0.850 3.970 1.060 ;
        RECT  3.560 0.850 3.850 0.920 ;
        RECT  3.650 0.215 3.770 0.415 ;
        RECT  3.370 0.345 3.650 0.415 ;
        RECT  3.440 0.850 3.560 1.060 ;
        RECT  2.975 0.850 3.440 0.920 ;
        RECT  3.255 0.205 3.370 0.415 ;
        RECT  3.070 0.205 3.185 0.415 ;
        RECT  2.810 0.345 3.070 0.415 ;
        RECT  2.905 0.850 2.975 1.065 ;
        RECT  0.220 0.995 2.905 1.065 ;
        RECT  2.690 0.205 2.810 0.415 ;
        RECT  2.430 0.345 2.690 0.415 ;
        RECT  2.310 0.205 2.430 0.415 ;
        RECT  2.050 0.345 2.310 0.415 ;
        RECT  1.930 0.205 2.050 0.415 ;
        RECT  1.685 0.345 1.930 0.415 ;
        RECT  1.615 0.210 1.685 0.415 ;
        RECT  0.130 0.210 1.615 0.280 ;
        RECT  0.050 0.210 0.130 0.370 ;
    END
END AOI22D8BWP40

MACRO AOI31D0BWP40
    CLASS CORE ;
    FOREIGN AOI31D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.099750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.200 0.740 0.270 ;
        RECT  0.455 0.200 0.525 0.915 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.805 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.930 0.295 ;
        RECT  0.150 -0.115 0.830 0.115 ;
        RECT  0.050 -0.115 0.150 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 1.145 0.980 1.375 ;
        RECT  0.835 0.965 0.935 1.375 ;
        RECT  0.000 1.145 0.835 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.915 0.740 1.055 ;
        RECT  0.230 0.985 0.620 1.055 ;
    END
END AOI31D0BWP40

MACRO AOI31D1BWP40
    CLASS CORE ;
    FOREIGN AOI31D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.181500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.215 0.740 0.305 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.455 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.930 0.400 ;
        RECT  0.150 -0.115 0.830 0.115 ;
        RECT  0.050 -0.115 0.150 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 1.145 0.980 1.375 ;
        RECT  0.835 0.860 0.935 1.375 ;
        RECT  0.000 1.145 0.835 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.845 0.740 1.055 ;
        RECT  0.230 0.985 0.620 1.055 ;
    END
END AOI31D1BWP40

MACRO AOI31D2BWP40
    CLASS CORE ;
    FOREIGN AOI31D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.305700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.195 1.525 0.405 ;
        RECT  1.365 0.335 1.415 0.405 ;
        RECT  1.285 0.335 1.365 0.920 ;
        RECT  1.140 0.335 1.285 0.405 ;
        RECT  0.220 0.850 1.285 0.920 ;
        RECT  1.070 0.205 1.140 0.405 ;
        RECT  0.595 0.205 1.070 0.275 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.785 0.625 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.195 0.780 ;
        RECT  0.255 0.710 1.115 0.780 ;
        RECT  0.170 0.495 0.255 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 1.000 0.630 ;
        RECT  0.435 0.345 0.875 0.415 ;
        RECT  0.345 0.345 0.435 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 -0.115 1.820 0.115 ;
        RECT  1.670 -0.115 1.750 0.400 ;
        RECT  1.290 -0.115 1.670 0.115 ;
        RECT  1.220 -0.115 1.290 0.255 ;
        RECT  0.130 -0.115 1.220 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.145 1.820 1.375 ;
        RECT  1.425 1.130 1.545 1.375 ;
        RECT  0.000 1.145 1.425 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.675 0.760 1.745 1.060 ;
        RECT  0.130 0.990 1.675 1.060 ;
        RECT  0.050 0.880 0.130 1.060 ;
    END
END AOI31D2BWP40

MACRO AOI31D4BWP40
    CLASS CORE ;
    FOREIGN AOI31D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.641200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.205 3.270 0.415 ;
        RECT  2.850 0.345 3.150 0.415 ;
        RECT  2.730 0.205 2.850 0.415 ;
        RECT  2.605 0.345 2.730 0.415 ;
        RECT  2.535 0.345 2.605 0.915 ;
        RECT  1.665 0.845 2.535 0.915 ;
        RECT  1.555 0.700 1.665 0.915 ;
        RECT  1.285 0.845 1.555 0.915 ;
        RECT  1.175 0.700 1.285 0.915 ;
        RECT  0.735 0.845 1.175 0.915 ;
        RECT  0.525 0.350 0.735 0.915 ;
        RECT  0.220 0.350 0.525 0.420 ;
        RECT  0.125 0.845 0.525 0.915 ;
        RECT  0.055 0.845 0.125 1.065 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.495 3.315 0.625 ;
        RECT  2.695 0.495 2.765 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.455 0.625 ;
        RECT  1.855 0.495 1.925 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.435 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.455 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.430 ;
        RECT  3.040 -0.115 3.370 0.115 ;
        RECT  2.960 -0.115 3.040 0.275 ;
        RECT  2.630 -0.115 2.960 0.115 ;
        RECT  2.550 -0.115 2.630 0.275 ;
        RECT  2.220 -0.115 2.550 0.115 ;
        RECT  2.140 -0.115 2.220 0.275 ;
        RECT  1.825 -0.115 2.140 0.115 ;
        RECT  1.755 -0.115 1.825 0.270 ;
        RECT  0.000 -0.115 1.755 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.145 3.500 1.375 ;
        RECT  3.150 0.890 3.270 1.375 ;
        RECT  2.850 1.145 3.150 1.375 ;
        RECT  2.730 1.125 2.850 1.375 ;
        RECT  0.000 1.145 2.730 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.205 3.270 0.415 ;
        RECT  2.850 0.345 3.150 0.415 ;
        RECT  2.730 0.205 2.850 0.415 ;
        RECT  2.605 0.345 2.730 0.415 ;
        RECT  2.535 0.345 2.605 0.915 ;
        RECT  1.665 0.845 2.535 0.915 ;
        RECT  1.555 0.700 1.665 0.915 ;
        RECT  1.285 0.845 1.555 0.915 ;
        RECT  1.175 0.700 1.285 0.915 ;
        RECT  0.805 0.845 1.175 0.915 ;
        RECT  0.220 0.350 0.455 0.420 ;
        RECT  0.125 0.845 0.455 0.915 ;
        RECT  0.055 0.845 0.125 1.065 ;
        RECT  3.370 0.750 3.450 1.030 ;
        RECT  3.040 0.750 3.370 0.820 ;
        RECT  2.965 0.750 3.040 1.055 ;
        RECT  0.220 0.985 2.965 1.055 ;
        RECT  2.325 0.205 2.445 0.415 ;
        RECT  2.040 0.345 2.325 0.415 ;
        RECT  1.920 0.205 2.040 0.415 ;
        RECT  0.980 0.345 1.920 0.415 ;
        RECT  0.130 0.205 1.670 0.275 ;
        RECT  0.050 0.205 0.130 0.370 ;
    END
END AOI31D4BWP40

MACRO AOI32D0BWP40
    CLASS CORE ;
    FOREIGN AOI32D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.099825 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.205 0.805 0.295 ;
        RECT  0.130 0.855 0.545 0.925 ;
        RECT  0.315 0.205 0.385 0.365 ;
        RECT  0.105 0.295 0.315 0.365 ;
        RECT  0.105 0.855 0.130 1.045 ;
        RECT  0.035 0.295 0.105 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.455 0.245 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.455 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.270 ;
        RECT  0.170 -0.115 1.130 0.115 ;
        RECT  0.050 -0.115 0.170 0.215 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 1.145 1.260 1.375 ;
        RECT  0.885 1.010 0.955 1.375 ;
        RECT  0.000 1.145 0.885 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.860 1.205 1.030 ;
        RECT  0.750 0.860 1.135 0.930 ;
        RECT  0.680 0.860 0.750 1.065 ;
        RECT  0.220 0.995 0.680 1.065 ;
    END
END AOI32D0BWP40

MACRO AOI32D1BWP40
    CLASS CORE ;
    FOREIGN AOI32D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.189250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.295 0.805 0.365 ;
        RECT  0.130 0.845 0.545 0.915 ;
        RECT  0.105 0.845 0.130 1.045 ;
        RECT  0.035 0.295 0.105 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.455 0.665 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 -0.115 1.260 0.115 ;
        RECT  1.130 -0.115 1.210 0.410 ;
        RECT  0.170 -0.115 1.130 0.115 ;
        RECT  0.050 -0.115 0.170 0.215 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 1.145 1.260 1.375 ;
        RECT  0.885 0.985 0.955 1.375 ;
        RECT  0.000 1.145 0.885 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.115 0.845 1.225 1.055 ;
        RECT  0.750 0.845 1.115 0.915 ;
        RECT  0.635 0.845 0.750 1.055 ;
        RECT  0.220 0.985 0.635 1.055 ;
    END
END AOI32D1BWP40

MACRO AOI32D2BWP40
    CLASS CORE ;
    FOREIGN AOI32D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.301100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.205 1.770 0.275 ;
        RECT  1.330 0.205 1.575 0.345 ;
        RECT  1.330 0.850 1.365 0.920 ;
        RECT  1.260 0.205 1.330 0.920 ;
        RECT  0.595 0.205 1.260 0.275 ;
        RECT  0.220 0.850 1.260 0.920 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.495 2.065 0.775 ;
        RECT  1.575 0.705 1.945 0.775 ;
        RECT  1.505 0.495 1.575 0.775 ;
        RECT  1.400 0.495 1.505 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.355 1.785 0.630 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 0.495 1.190 0.780 ;
        RECT  0.255 0.710 1.110 0.780 ;
        RECT  0.170 0.495 0.255 0.780 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.345 1.015 0.640 ;
        RECT  0.435 0.345 0.875 0.415 ;
        RECT  0.325 0.345 0.435 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 -0.115 2.240 0.115 ;
        RECT  2.110 -0.115 2.190 0.420 ;
        RECT  1.360 -0.115 2.110 0.115 ;
        RECT  1.240 -0.115 1.360 0.135 ;
        RECT  0.130 -0.115 1.240 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.970 1.145 2.240 1.375 ;
        RECT  1.850 1.015 1.970 1.375 ;
        RECT  1.570 1.145 1.850 1.375 ;
        RECT  1.450 1.130 1.570 1.375 ;
        RECT  0.000 1.145 1.450 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.110 0.875 2.190 1.055 ;
        RECT  1.515 0.875 2.110 0.945 ;
        RECT  1.445 0.875 1.515 1.060 ;
        RECT  0.130 0.990 1.445 1.060 ;
        RECT  0.050 0.875 0.130 1.060 ;
    END
END AOI32D2BWP40

MACRO AOI32D4BWP40
    CLASS CORE ;
    FOREIGN AOI32D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.643000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.195 3.370 0.265 ;
        RECT  2.555 0.195 2.560 0.415 ;
        RECT  2.490 0.195 2.555 0.815 ;
        RECT  2.345 0.345 2.490 0.815 ;
        RECT  1.735 0.345 2.345 0.415 ;
        RECT  2.275 0.745 2.345 0.815 ;
        RECT  2.205 0.745 2.275 0.915 ;
        RECT  0.220 0.845 2.205 0.915 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 4.165 0.630 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.495 3.325 0.630 ;
        RECT  2.695 0.495 2.765 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.805 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.765 ;
        RECT  0.940 0.495 1.435 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.210 0.625 ;
        RECT  1.855 0.495 1.925 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.210 -0.115 4.290 0.420 ;
        RECT  3.935 -0.115 4.210 0.115 ;
        RECT  3.810 -0.115 3.935 0.255 ;
        RECT  3.530 -0.115 3.810 0.115 ;
        RECT  3.450 -0.115 3.530 0.265 ;
        RECT  0.725 -0.115 3.450 0.115 ;
        RECT  0.595 -0.115 0.725 0.230 ;
        RECT  0.345 -0.115 0.595 0.115 ;
        RECT  0.215 -0.115 0.345 0.230 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.145 4.340 1.375 ;
        RECT  3.995 1.030 4.125 1.375 ;
        RECT  3.740 1.145 3.995 1.375 ;
        RECT  3.615 1.025 3.740 1.375 ;
        RECT  3.180 1.145 3.615 1.375 ;
        RECT  3.060 1.025 3.180 1.375 ;
        RECT  2.800 1.145 3.060 1.375 ;
        RECT  2.680 1.025 2.800 1.375 ;
        RECT  0.000 1.145 2.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.625 0.195 3.370 0.265 ;
        RECT  1.735 0.345 2.275 0.415 ;
        RECT  2.205 0.745 2.275 0.915 ;
        RECT  0.220 0.845 2.205 0.915 ;
        RECT  4.195 0.745 4.305 0.955 ;
        RECT  3.925 0.885 4.195 0.955 ;
        RECT  2.665 0.345 4.125 0.415 ;
        RECT  3.815 0.745 3.925 0.955 ;
        RECT  3.365 0.885 3.815 0.955 ;
        RECT  3.255 0.745 3.365 0.955 ;
        RECT  2.985 0.885 3.255 0.955 ;
        RECT  2.875 0.745 2.985 0.955 ;
        RECT  2.600 0.885 2.875 0.955 ;
        RECT  2.510 0.885 2.600 1.065 ;
        RECT  0.130 0.995 2.510 1.065 ;
        RECT  0.975 0.195 2.420 0.265 ;
        RECT  0.035 0.345 1.665 0.415 ;
        RECT  0.050 0.940 0.130 1.065 ;
    END
END AOI32D4BWP40

MACRO AOI33D0BWP40
    CLASS CORE ;
    FOREIGN AOI33D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.110975 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.235 0.760 0.325 ;
        RECT  0.455 0.235 0.525 0.815 ;
        RECT  0.125 0.745 0.455 0.815 ;
        RECT  0.035 0.745 0.125 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.365 0.625 ;
        RECT  1.155 0.495 1.225 0.770 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.390 1.085 0.770 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.770 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.440 0.665 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.315 ;
        RECT  0.140 -0.115 1.260 0.115 ;
        RECT  0.040 -0.115 0.140 0.325 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.985 1.360 1.375 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.840 0.990 0.960 1.375 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.850 1.170 1.060 ;
        RECT  0.735 0.850 1.050 0.920 ;
        RECT  0.665 0.850 0.735 1.065 ;
        RECT  0.220 0.995 0.665 1.065 ;
    END
END AOI33D0BWP40

MACRO AOI33D1BWP40
    CLASS CORE ;
    FOREIGN AOI33D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.183250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.235 0.760 0.325 ;
        RECT  0.455 0.235 0.525 0.815 ;
        RECT  0.125 0.745 0.455 0.815 ;
        RECT  0.035 0.745 0.125 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.390 1.085 0.770 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.770 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.440 0.665 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.415 ;
        RECT  0.140 -0.115 1.260 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.705 1.360 1.375 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.840 0.990 0.960 1.375 ;
        RECT  0.000 1.145 0.840 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.850 1.170 1.060 ;
        RECT  0.755 0.850 1.050 0.920 ;
        RECT  0.645 0.850 0.755 1.065 ;
        RECT  0.220 0.995 0.645 1.065 ;
    END
END AOI33D1BWP40

MACRO AOI33D2BWP40
    CLASS CORE ;
    FOREIGN AOI33D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.304450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.340 2.485 0.795 ;
        RECT  2.270 0.340 2.415 0.410 ;
        RECT  2.300 0.725 2.415 0.795 ;
        RECT  2.230 0.725 2.300 0.925 ;
        RECT  2.200 0.200 2.270 0.410 ;
        RECT  1.365 0.855 2.230 0.925 ;
        RECT  0.595 0.200 2.200 0.270 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.525 1.225 0.640 ;
        RECT  1.085 0.340 1.155 0.640 ;
        RECT  0.245 0.340 1.085 0.410 ;
        RECT  0.175 0.340 0.245 0.765 ;
        RECT  0.130 0.520 0.175 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.495 1.015 0.775 ;
        RECT  0.405 0.705 0.915 0.775 ;
        RECT  0.315 0.495 0.405 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.495 0.845 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.059600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.480 2.345 0.645 ;
        RECT  2.130 0.480 2.245 0.550 ;
        RECT  1.995 0.340 2.130 0.550 ;
        RECT  1.365 0.340 1.995 0.410 ;
        RECT  1.295 0.340 1.365 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.059600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.620 2.150 0.775 ;
        RECT  1.585 0.705 1.995 0.775 ;
        RECT  1.435 0.495 1.585 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.059600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.495 1.925 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.460 -0.115 2.520 0.115 ;
        RECT  2.360 -0.115 2.460 0.270 ;
        RECT  1.300 -0.115 2.360 0.115 ;
        RECT  1.180 -0.115 1.300 0.130 ;
        RECT  0.130 -0.115 1.180 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.145 2.520 1.375 ;
        RECT  0.980 0.985 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 0.985 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.380 0.915 2.450 1.065 ;
        RECT  1.265 0.995 2.380 1.065 ;
        RECT  0.125 0.845 1.195 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
        RECT  1.195 0.755 1.265 1.065 ;
    END
END AOI33D2BWP40

MACRO AOI33D4BWP40
    CLASS CORE ;
    FOREIGN AOI33D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.643000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.345 3.365 0.415 ;
        RECT  2.345 0.345 2.555 0.815 ;
        RECT  1.735 0.345 2.345 0.415 ;
        RECT  2.275 0.745 2.345 0.815 ;
        RECT  2.205 0.745 2.275 0.915 ;
        RECT  0.220 0.845 2.205 0.915 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.495 5.005 0.630 ;
        RECT  4.375 0.495 4.445 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 4.165 0.630 ;
        RECT  3.535 0.495 3.605 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.185 0.765 ;
        RECT  2.675 0.495 3.115 0.630 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.805 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.765 ;
        RECT  0.940 0.495 1.435 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.210 0.625 ;
        RECT  1.855 0.495 1.925 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.875 -0.115 5.180 0.115 ;
        RECT  4.765 -0.115 4.875 0.240 ;
        RECT  4.495 -0.115 4.765 0.115 ;
        RECT  4.385 -0.115 4.495 0.240 ;
        RECT  0.725 -0.115 4.385 0.115 ;
        RECT  0.595 -0.115 0.725 0.265 ;
        RECT  0.345 -0.115 0.595 0.115 ;
        RECT  0.215 -0.115 0.345 0.265 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.885 1.145 5.180 1.375 ;
        RECT  4.755 1.030 4.885 1.375 ;
        RECT  4.505 1.145 4.755 1.375 ;
        RECT  4.375 1.030 4.505 1.375 ;
        RECT  4.125 1.145 4.375 1.375 ;
        RECT  3.995 1.030 4.125 1.375 ;
        RECT  3.740 1.145 3.995 1.375 ;
        RECT  3.615 1.025 3.740 1.375 ;
        RECT  3.180 1.145 3.615 1.375 ;
        RECT  3.060 1.025 3.180 1.375 ;
        RECT  2.800 1.145 3.060 1.375 ;
        RECT  2.680 1.025 2.800 1.375 ;
        RECT  0.000 1.145 2.680 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.625 0.345 3.365 0.415 ;
        RECT  1.735 0.345 2.275 0.415 ;
        RECT  2.205 0.745 2.275 0.915 ;
        RECT  0.220 0.845 2.205 0.915 ;
        RECT  5.010 0.205 5.120 0.415 ;
        RECT  5.005 0.745 5.115 0.955 ;
        RECT  4.685 0.345 5.010 0.415 ;
        RECT  4.685 0.885 5.005 0.955 ;
        RECT  4.575 0.205 4.685 0.415 ;
        RECT  4.575 0.745 4.685 0.955 ;
        RECT  4.305 0.345 4.575 0.415 ;
        RECT  4.305 0.885 4.575 0.955 ;
        RECT  4.195 0.205 4.305 0.415 ;
        RECT  4.195 0.745 4.305 0.955 ;
        RECT  3.435 0.345 4.195 0.415 ;
        RECT  3.925 0.885 4.195 0.955 ;
        RECT  2.665 0.195 4.115 0.265 ;
        RECT  3.815 0.745 3.925 0.955 ;
        RECT  3.365 0.885 3.815 0.955 ;
        RECT  3.255 0.745 3.365 0.955 ;
        RECT  2.985 0.885 3.255 0.955 ;
        RECT  2.875 0.745 2.985 0.955 ;
        RECT  2.590 0.885 2.875 0.955 ;
        RECT  2.510 0.885 2.590 1.065 ;
        RECT  0.130 0.995 2.510 1.065 ;
        RECT  0.975 0.195 2.420 0.265 ;
        RECT  0.035 0.345 1.665 0.415 ;
        RECT  0.050 0.940 0.130 1.065 ;
    END
END AOI33D4BWP40

MACRO BUFFD0BWP40
    CLASS CORE ;
    FOREIGN BUFFD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 1.045 ;
        RECT  0.435 0.185 0.455 0.305 ;
        RECT  0.435 0.905 0.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.520 0.385 0.640 ;
        RECT  0.295 0.335 0.365 0.925 ;
        RECT  0.130 0.335 0.295 0.405 ;
        RECT  0.130 0.855 0.295 0.925 ;
        RECT  0.050 0.195 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END BUFFD0BWP40

MACRO BUFFD10BWP40
    CLASS CORE ;
    FOREIGN BUFFD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.600000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  1.995 0.305 2.195 0.465 ;
        RECT  1.885 0.305 1.995 0.950 ;
        RECT  1.815 0.185 1.885 0.950 ;
        RECT  1.785 0.305 1.815 0.950 ;
        RECT  1.505 0.305 1.785 0.465 ;
        RECT  1.030 0.720 1.785 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 2.940 0.115 ;
        RECT  2.760 -0.115 2.840 0.465 ;
        RECT  2.480 -0.115 2.760 0.115 ;
        RECT  2.360 -0.115 2.480 0.235 ;
        RECT  2.100 -0.115 2.360 0.115 ;
        RECT  1.980 -0.115 2.100 0.235 ;
        RECT  1.720 -0.115 1.980 0.115 ;
        RECT  1.600 -0.115 1.720 0.235 ;
        RECT  1.340 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.340 0.235 ;
        RECT  0.940 -0.115 1.220 0.115 ;
        RECT  0.860 -0.115 0.940 0.465 ;
        RECT  0.565 -0.115 0.860 0.115 ;
        RECT  0.475 -0.115 0.565 0.260 ;
        RECT  0.190 -0.115 0.475 0.115 ;
        RECT  0.090 -0.115 0.190 0.410 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.145 2.940 1.375 ;
        RECT  2.760 0.700 2.840 1.375 ;
        RECT  2.480 1.145 2.760 1.375 ;
        RECT  2.360 1.020 2.480 1.375 ;
        RECT  2.100 1.145 2.360 1.375 ;
        RECT  1.980 1.020 2.100 1.375 ;
        RECT  1.720 1.145 1.980 1.375 ;
        RECT  1.600 1.020 1.720 1.375 ;
        RECT  1.340 1.145 1.600 1.375 ;
        RECT  1.220 1.020 1.340 1.375 ;
        RECT  0.940 1.145 1.220 1.375 ;
        RECT  0.860 0.720 0.940 1.375 ;
        RECT  0.560 1.145 0.860 1.375 ;
        RECT  0.480 0.885 0.560 1.375 ;
        RECT  0.190 1.145 0.480 1.375 ;
        RECT  0.090 0.845 0.190 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.065 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  2.065 0.305 2.195 0.465 ;
        RECT  1.505 0.305 1.715 0.465 ;
        RECT  1.030 0.720 1.715 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  0.770 0.545 1.705 0.615 ;
        RECT  0.660 0.195 0.770 1.050 ;
        RECT  0.390 0.335 0.660 0.415 ;
        RECT  0.365 0.725 0.660 0.805 ;
        RECT  0.270 0.205 0.390 0.415 ;
        RECT  0.295 0.725 0.365 1.050 ;
    END
END BUFFD10BWP40

MACRO BUFFD12BWP40
    CLASS CORE ;
    FOREIGN BUFFD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.275 0.305 2.525 0.465 ;
        RECT  2.215 0.305 2.275 0.950 ;
        RECT  2.135 0.185 2.215 0.950 ;
        RECT  1.925 0.305 2.135 0.950 ;
        RECT  1.835 0.305 1.925 0.465 ;
        RECT  0.980 0.720 1.925 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.465 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.235 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.235 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.890 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.890 0.465 ;
        RECT  0.515 -0.115 0.810 0.115 ;
        RECT  0.425 -0.115 0.515 0.260 ;
        RECT  0.140 -0.115 0.425 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.700 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 1.020 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 1.020 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 1.020 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.020 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 1.020 1.290 1.375 ;
        RECT  0.890 1.145 1.170 1.375 ;
        RECT  0.810 0.720 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.995 0.510 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.345 0.305 2.525 0.465 ;
        RECT  1.835 0.305 1.855 0.465 ;
        RECT  0.980 0.720 1.855 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  0.720 0.545 1.765 0.615 ;
        RECT  0.610 0.195 0.720 1.050 ;
        RECT  0.340 0.335 0.610 0.415 ;
        RECT  0.315 0.775 0.610 0.855 ;
        RECT  0.220 0.205 0.340 0.415 ;
        RECT  0.245 0.775 0.315 1.050 ;
    END
END BUFFD12BWP40

MACRO BUFFD14BWP40
    CLASS CORE ;
    FOREIGN BUFFD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.872000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.835 0.305 3.125 0.465 ;
        RECT  2.815 0.305 2.835 0.945 ;
        RECT  2.745 0.185 2.815 0.945 ;
        RECT  2.485 0.305 2.745 0.945 ;
        RECT  2.435 0.305 2.485 0.465 ;
        RECT  1.200 0.715 2.485 0.945 ;
        RECT  2.365 0.185 2.435 0.465 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.160000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.665 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 -0.115 3.920 0.115 ;
        RECT  3.730 -0.115 3.835 0.465 ;
        RECT  3.410 -0.115 3.730 0.115 ;
        RECT  3.290 -0.115 3.410 0.235 ;
        RECT  3.030 -0.115 3.290 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.650 -0.115 2.910 0.115 ;
        RECT  2.530 -0.115 2.650 0.235 ;
        RECT  2.270 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.270 0.235 ;
        RECT  1.890 -0.115 2.150 0.115 ;
        RECT  1.770 -0.115 1.890 0.235 ;
        RECT  1.510 -0.115 1.770 0.115 ;
        RECT  1.390 -0.115 1.510 0.235 ;
        RECT  1.100 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.100 0.465 ;
        RECT  0.720 -0.115 1.020 0.115 ;
        RECT  0.600 -0.115 0.720 0.265 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 1.145 3.920 1.375 ;
        RECT  3.730 0.690 3.835 1.375 ;
        RECT  3.410 1.145 3.730 1.375 ;
        RECT  3.290 1.015 3.410 1.375 ;
        RECT  3.030 1.145 3.290 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.650 1.145 2.910 1.375 ;
        RECT  2.530 1.015 2.650 1.375 ;
        RECT  2.270 1.145 2.530 1.375 ;
        RECT  2.150 1.015 2.270 1.375 ;
        RECT  1.890 1.145 2.150 1.375 ;
        RECT  1.770 1.015 1.890 1.375 ;
        RECT  1.510 1.145 1.770 1.375 ;
        RECT  1.390 1.015 1.510 1.375 ;
        RECT  1.120 1.145 1.390 1.375 ;
        RECT  1.000 0.710 1.120 1.375 ;
        RECT  0.700 1.145 1.000 1.375 ;
        RECT  0.620 0.860 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 1.000 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.905 0.305 3.125 0.465 ;
        RECT  2.365 0.185 2.415 0.465 ;
        RECT  1.200 0.715 2.415 0.945 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        RECT  0.920 0.545 2.405 0.615 ;
        RECT  0.790 0.195 0.920 1.065 ;
        RECT  0.510 0.335 0.790 0.415 ;
        RECT  0.505 0.705 0.790 0.785 ;
        RECT  0.430 0.185 0.510 0.415 ;
        RECT  0.435 0.705 0.505 1.035 ;
        RECT  0.125 0.850 0.435 0.920 ;
        RECT  0.130 0.335 0.430 0.415 ;
        RECT  0.055 0.255 0.130 0.415 ;
        RECT  0.055 0.850 0.125 1.035 ;
    END
END BUFFD14BWP40

MACRO BUFFD16BWP40
    CLASS CORE ;
    FOREIGN BUFFD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.115 0.305 3.405 0.465 ;
        RECT  3.095 0.305 3.115 0.945 ;
        RECT  3.025 0.185 3.095 0.945 ;
        RECT  2.765 0.305 3.025 0.945 ;
        RECT  2.715 0.305 2.765 0.465 ;
        RECT  1.480 0.715 2.765 0.945 ;
        RECT  2.645 0.185 2.715 0.465 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.945 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.465 ;
        RECT  4.070 -0.115 4.350 0.115 ;
        RECT  3.950 -0.115 4.070 0.235 ;
        RECT  3.690 -0.115 3.950 0.115 ;
        RECT  3.570 -0.115 3.690 0.235 ;
        RECT  3.310 -0.115 3.570 0.115 ;
        RECT  3.190 -0.115 3.310 0.235 ;
        RECT  2.930 -0.115 3.190 0.115 ;
        RECT  2.810 -0.115 2.930 0.235 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.235 ;
        RECT  2.170 -0.115 2.430 0.115 ;
        RECT  2.050 -0.115 2.170 0.235 ;
        RECT  1.790 -0.115 2.050 0.115 ;
        RECT  1.670 -0.115 1.790 0.235 ;
        RECT  1.380 -0.115 1.670 0.115 ;
        RECT  1.300 -0.115 1.380 0.465 ;
        RECT  1.000 -0.115 1.300 0.115 ;
        RECT  0.880 -0.115 1.000 0.265 ;
        RECT  0.620 -0.115 0.880 0.115 ;
        RECT  0.500 -0.115 0.620 0.265 ;
        RECT  0.180 -0.115 0.500 0.115 ;
        RECT  0.060 -0.115 0.180 0.415 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.690 4.430 1.375 ;
        RECT  4.070 1.145 4.350 1.375 ;
        RECT  3.950 1.015 4.070 1.375 ;
        RECT  3.690 1.145 3.950 1.375 ;
        RECT  3.570 1.015 3.690 1.375 ;
        RECT  3.310 1.145 3.570 1.375 ;
        RECT  3.190 1.015 3.310 1.375 ;
        RECT  2.930 1.145 3.190 1.375 ;
        RECT  2.810 1.015 2.930 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 1.015 2.550 1.375 ;
        RECT  2.170 1.145 2.430 1.375 ;
        RECT  2.050 1.015 2.170 1.375 ;
        RECT  1.790 1.145 2.050 1.375 ;
        RECT  1.670 1.015 1.790 1.375 ;
        RECT  1.400 1.145 1.670 1.375 ;
        RECT  1.280 0.710 1.400 1.375 ;
        RECT  0.980 1.145 1.280 1.375 ;
        RECT  0.900 0.860 0.980 1.375 ;
        RECT  0.600 1.145 0.900 1.375 ;
        RECT  0.520 0.860 0.600 1.375 ;
        RECT  0.170 1.145 0.520 1.375 ;
        RECT  0.090 0.845 0.170 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.185 0.305 3.405 0.465 ;
        RECT  2.645 0.185 2.695 0.465 ;
        RECT  1.480 0.715 2.695 0.945 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        RECT  1.200 0.545 2.685 0.615 ;
        RECT  1.070 0.195 1.200 1.065 ;
        RECT  0.790 0.335 1.070 0.415 ;
        RECT  0.785 0.705 1.070 0.785 ;
        RECT  0.710 0.185 0.790 0.415 ;
        RECT  0.715 0.705 0.785 1.035 ;
        RECT  0.405 0.705 0.715 0.785 ;
        RECT  0.410 0.335 0.710 0.415 ;
        RECT  0.310 0.185 0.410 0.415 ;
        RECT  0.335 0.705 0.405 1.035 ;
    END
END BUFFD16BWP40

MACRO BUFFD18BWP40
    CLASS CORE ;
    FOREIGN BUFFD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.080000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.105 0.305 3.305 0.465 ;
        RECT  2.995 0.305 3.105 0.945 ;
        RECT  2.925 0.185 2.995 0.945 ;
        RECT  2.765 0.305 2.925 0.945 ;
        RECT  2.615 0.305 2.765 0.465 ;
        RECT  1.380 0.715 2.765 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  1.405 0.185 1.475 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.855 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.350 -0.115 4.630 0.115 ;
        RECT  4.230 -0.115 4.350 0.235 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.235 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.235 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.235 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.235 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.235 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.235 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.235 ;
        RECT  1.280 -0.115 1.570 0.115 ;
        RECT  1.200 -0.115 1.280 0.465 ;
        RECT  0.910 -0.115 1.200 0.115 ;
        RECT  0.790 -0.115 0.910 0.265 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.265 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.690 4.710 1.375 ;
        RECT  4.350 1.145 4.630 1.375 ;
        RECT  4.230 1.015 4.350 1.375 ;
        RECT  3.970 1.145 4.230 1.375 ;
        RECT  3.850 1.015 3.970 1.375 ;
        RECT  3.590 1.145 3.850 1.375 ;
        RECT  3.470 1.015 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.090 1.015 3.210 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.015 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.330 1.015 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 1.015 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.570 1.015 1.690 1.375 ;
        RECT  1.300 1.145 1.570 1.375 ;
        RECT  1.180 0.710 1.300 1.375 ;
        RECT  0.890 1.145 1.180 1.375 ;
        RECT  0.810 0.860 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.860 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.185 0.305 3.305 0.465 ;
        RECT  2.615 0.305 2.695 0.465 ;
        RECT  1.380 0.715 2.695 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.110 0.545 2.585 0.615 ;
        RECT  0.980 0.195 1.110 1.065 ;
        RECT  0.700 0.335 0.980 0.415 ;
        RECT  0.695 0.705 0.980 0.785 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.625 0.705 0.695 1.035 ;
        RECT  0.315 0.705 0.625 0.785 ;
        RECT  0.320 0.335 0.620 0.415 ;
        RECT  0.220 0.185 0.320 0.415 ;
        RECT  0.245 0.705 0.315 1.035 ;
    END
END BUFFD18BWP40

MACRO BUFFD1BWP40
    CLASS CORE ;
    FOREIGN BUFFD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 1.045 ;
        RECT  0.435 0.185 0.455 0.465 ;
        RECT  0.435 0.735 0.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.520 0.385 0.640 ;
        RECT  0.295 0.335 0.365 0.925 ;
        RECT  0.130 0.335 0.295 0.405 ;
        RECT  0.130 0.855 0.295 0.925 ;
        RECT  0.050 0.195 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END BUFFD1BWP40

MACRO BUFFD20BWP40
    CLASS CORE ;
    FOREIGN BUFFD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.200000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.555 0.305 3.865 0.465 ;
        RECT  3.535 0.185 3.555 0.465 ;
        RECT  3.485 0.185 3.535 0.960 ;
        RECT  3.185 0.305 3.485 0.960 ;
        RECT  3.175 0.305 3.185 0.465 ;
        RECT  1.560 0.730 3.185 0.960 ;
        RECT  3.105 0.185 3.175 0.465 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.224000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.065 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.910 -0.115 5.190 0.115 ;
        RECT  4.790 -0.115 4.910 0.235 ;
        RECT  4.530 -0.115 4.790 0.115 ;
        RECT  4.410 -0.115 4.530 0.235 ;
        RECT  4.150 -0.115 4.410 0.115 ;
        RECT  4.030 -0.115 4.150 0.235 ;
        RECT  3.770 -0.115 4.030 0.115 ;
        RECT  3.650 -0.115 3.770 0.235 ;
        RECT  3.390 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.010 -0.115 3.270 0.115 ;
        RECT  2.890 -0.115 3.010 0.235 ;
        RECT  2.630 -0.115 2.890 0.115 ;
        RECT  2.510 -0.115 2.630 0.235 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.235 ;
        RECT  1.870 -0.115 2.130 0.115 ;
        RECT  1.750 -0.115 1.870 0.235 ;
        RECT  1.465 -0.115 1.750 0.115 ;
        RECT  1.395 -0.115 1.465 0.465 ;
        RECT  1.085 -0.115 1.395 0.115 ;
        RECT  1.015 -0.115 1.085 0.255 ;
        RECT  0.695 -0.115 1.015 0.115 ;
        RECT  0.625 -0.115 0.695 0.255 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.245 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.700 5.270 1.375 ;
        RECT  4.910 1.145 5.190 1.375 ;
        RECT  4.790 1.030 4.910 1.375 ;
        RECT  4.530 1.145 4.790 1.375 ;
        RECT  4.410 1.030 4.530 1.375 ;
        RECT  4.150 1.145 4.410 1.375 ;
        RECT  4.030 1.030 4.150 1.375 ;
        RECT  3.770 1.145 4.030 1.375 ;
        RECT  3.650 1.030 3.770 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.030 3.390 1.375 ;
        RECT  3.010 1.145 3.270 1.375 ;
        RECT  2.890 1.030 3.010 1.375 ;
        RECT  2.630 1.145 2.890 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.250 1.145 2.510 1.375 ;
        RECT  2.130 1.030 2.250 1.375 ;
        RECT  1.870 1.145 2.130 1.375 ;
        RECT  1.750 1.030 1.870 1.375 ;
        RECT  1.465 1.145 1.750 1.375 ;
        RECT  1.395 0.720 1.465 1.375 ;
        RECT  1.085 1.145 1.395 1.375 ;
        RECT  1.015 0.860 1.085 1.375 ;
        RECT  0.710 1.145 1.015 1.375 ;
        RECT  0.610 0.860 0.710 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.605 0.305 3.865 0.465 ;
        RECT  3.105 0.185 3.115 0.465 ;
        RECT  1.560 0.730 3.115 0.960 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        RECT  1.315 0.545 3.105 0.615 ;
        RECT  1.155 0.185 1.315 1.065 ;
        RECT  0.895 0.335 1.155 0.415 ;
        RECT  0.920 0.700 1.155 0.780 ;
        RECT  0.800 0.700 0.920 1.065 ;
        RECT  0.825 0.185 0.895 0.415 ;
        RECT  0.505 0.335 0.825 0.415 ;
        RECT  0.530 0.700 0.800 0.780 ;
        RECT  0.410 0.700 0.530 1.065 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.130 0.335 0.435 0.415 ;
        RECT  0.125 0.845 0.410 0.925 ;
        RECT  0.055 0.275 0.130 0.415 ;
        RECT  0.055 0.845 0.125 0.985 ;
    END
END BUFFD20BWP40

MACRO BUFFD24BWP40
    CLASS CORE ;
    FOREIGN BUFFD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.440000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.155 0.305 4.465 0.465 ;
        RECT  4.095 0.185 4.155 0.465 ;
        RECT  4.085 0.185 4.095 0.945 ;
        RECT  3.775 0.305 4.085 0.945 ;
        RECT  3.745 0.185 3.775 0.945 ;
        RECT  3.705 0.185 3.745 0.465 ;
        RECT  1.780 0.715 3.745 0.945 ;
        RECT  3.395 0.305 3.705 0.465 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.155 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.475 ;
        RECT  5.890 -0.115 6.170 0.115 ;
        RECT  5.770 -0.115 5.890 0.235 ;
        RECT  5.510 -0.115 5.770 0.115 ;
        RECT  5.390 -0.115 5.510 0.235 ;
        RECT  5.130 -0.115 5.390 0.115 ;
        RECT  5.010 -0.115 5.130 0.235 ;
        RECT  4.750 -0.115 5.010 0.115 ;
        RECT  4.630 -0.115 4.750 0.235 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.235 ;
        RECT  3.990 -0.115 4.250 0.115 ;
        RECT  3.870 -0.115 3.990 0.235 ;
        RECT  3.610 -0.115 3.870 0.115 ;
        RECT  3.490 -0.115 3.610 0.235 ;
        RECT  3.230 -0.115 3.490 0.115 ;
        RECT  3.110 -0.115 3.230 0.235 ;
        RECT  2.850 -0.115 3.110 0.115 ;
        RECT  2.730 -0.115 2.850 0.235 ;
        RECT  2.470 -0.115 2.730 0.115 ;
        RECT  2.350 -0.115 2.470 0.235 ;
        RECT  2.090 -0.115 2.350 0.115 ;
        RECT  1.970 -0.115 2.090 0.235 ;
        RECT  1.685 -0.115 1.970 0.115 ;
        RECT  1.615 -0.115 1.685 0.465 ;
        RECT  1.295 -0.115 1.615 0.115 ;
        RECT  1.225 -0.115 1.295 0.245 ;
        RECT  0.895 -0.115 1.225 0.115 ;
        RECT  0.825 -0.115 0.895 0.245 ;
        RECT  0.505 -0.115 0.825 0.115 ;
        RECT  0.435 -0.115 0.505 0.245 ;
        RECT  0.125 -0.115 0.435 0.115 ;
        RECT  0.055 -0.115 0.125 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.720 6.250 1.375 ;
        RECT  5.890 1.145 6.170 1.375 ;
        RECT  5.770 1.015 5.890 1.375 ;
        RECT  5.510 1.145 5.770 1.375 ;
        RECT  5.390 1.015 5.510 1.375 ;
        RECT  5.130 1.145 5.390 1.375 ;
        RECT  5.010 1.015 5.130 1.375 ;
        RECT  4.750 1.145 5.010 1.375 ;
        RECT  4.630 1.015 4.750 1.375 ;
        RECT  4.370 1.145 4.630 1.375 ;
        RECT  4.250 1.015 4.370 1.375 ;
        RECT  3.990 1.145 4.250 1.375 ;
        RECT  3.870 1.015 3.990 1.375 ;
        RECT  3.610 1.145 3.870 1.375 ;
        RECT  3.490 1.015 3.610 1.375 ;
        RECT  3.230 1.145 3.490 1.375 ;
        RECT  3.110 1.015 3.230 1.375 ;
        RECT  2.850 1.145 3.110 1.375 ;
        RECT  2.730 1.015 2.850 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 1.015 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 1.015 2.090 1.375 ;
        RECT  1.685 1.145 1.970 1.375 ;
        RECT  1.615 0.740 1.685 1.375 ;
        RECT  1.295 1.145 1.615 1.375 ;
        RECT  1.225 0.880 1.295 1.375 ;
        RECT  0.900 1.145 1.225 1.375 ;
        RECT  0.820 0.880 0.900 1.375 ;
        RECT  0.510 1.145 0.820 1.375 ;
        RECT  0.430 0.880 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.165 0.305 4.465 0.465 ;
        RECT  3.395 0.305 3.675 0.465 ;
        RECT  1.780 0.715 3.675 0.945 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        RECT  1.535 0.545 3.645 0.615 ;
        RECT  1.365 0.195 1.535 1.070 ;
        RECT  1.100 0.325 1.365 0.415 ;
        RECT  1.120 0.705 1.365 0.795 ;
        RECT  1.000 0.705 1.120 1.070 ;
        RECT  1.020 0.185 1.100 0.415 ;
        RECT  0.700 0.325 1.020 0.415 ;
        RECT  0.720 0.705 1.000 0.795 ;
        RECT  0.600 0.705 0.720 1.070 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.320 0.325 0.620 0.415 ;
        RECT  0.340 0.705 0.600 0.795 ;
        RECT  0.220 0.705 0.340 1.065 ;
        RECT  0.220 0.185 0.320 0.415 ;
    END
END BUFFD24BWP40

MACRO BUFFD2BWP40
    CLASS CORE ;
    FOREIGN BUFFD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.152000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.385 0.805 0.875 ;
        RECT  0.555 0.385 0.735 0.455 ;
        RECT  0.555 0.775 0.735 0.875 ;
        RECT  0.465 0.185 0.555 0.455 ;
        RECT  0.465 0.775 0.555 1.065 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.245 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 -0.115 0.840 0.115 ;
        RECT  0.660 -0.115 0.780 0.265 ;
        RECT  0.340 -0.115 0.660 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.145 0.840 1.375 ;
        RECT  0.660 0.995 0.780 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.395 0.545 0.535 0.615 ;
        RECT  0.325 0.335 0.395 0.925 ;
        RECT  0.130 0.335 0.325 0.405 ;
        RECT  0.130 0.855 0.325 0.925 ;
        RECT  0.050 0.195 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END BUFFD2BWP40

MACRO BUFFD3BWP40
    CLASS CORE ;
    FOREIGN BUFFD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.185 0.945 0.490 ;
        RECT  0.875 0.700 0.945 1.045 ;
        RECT  0.855 0.185 0.875 1.045 ;
        RECT  0.665 0.355 0.855 0.820 ;
        RECT  0.545 0.355 0.665 0.475 ;
        RECT  0.545 0.700 0.665 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.280 ;
        RECT  0.360 -0.115 0.640 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 0.890 0.760 1.375 ;
        RECT  0.360 1.145 0.640 1.375 ;
        RECT  0.240 0.995 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.545 0.355 0.595 0.475 ;
        RECT  0.545 0.700 0.595 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        RECT  0.395 0.545 0.575 0.615 ;
        RECT  0.325 0.345 0.395 0.925 ;
        RECT  0.130 0.345 0.325 0.415 ;
        RECT  0.130 0.855 0.325 0.925 ;
        RECT  0.050 0.245 0.130 0.415 ;
        RECT  0.050 0.855 0.130 1.025 ;
    END
END BUFFD3BWP40

MACRO BUFFD4BWP40
    CLASS CORE ;
    FOREIGN BUFFD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  1.055 0.700 1.125 1.045 ;
        RECT  1.015 0.355 1.055 0.465 ;
        RECT  1.015 0.700 1.055 0.820 ;
        RECT  0.805 0.355 1.015 0.820 ;
        RECT  0.725 0.355 0.805 0.465 ;
        RECT  0.725 0.700 0.805 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.390 0.765 ;
        RECT  0.175 0.495 0.315 0.635 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.475 ;
        RECT  0.950 -0.115 1.270 0.115 ;
        RECT  0.830 -0.115 0.950 0.280 ;
        RECT  0.530 -0.115 0.830 0.115 ;
        RECT  0.450 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.450 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.270 0.700 1.350 1.375 ;
        RECT  0.950 1.145 1.270 1.375 ;
        RECT  0.830 0.890 0.950 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.440 0.975 0.540 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.185 1.125 0.465 ;
        RECT  1.085 0.700 1.125 1.045 ;
        RECT  0.725 0.355 0.735 0.465 ;
        RECT  0.725 0.700 0.735 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  0.585 0.545 0.720 0.615 ;
        RECT  0.510 0.345 0.585 0.905 ;
        RECT  0.325 0.345 0.510 0.415 ;
        RECT  0.325 0.835 0.510 0.905 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.835 0.325 0.995 ;
    END
END BUFFD4BWP40

MACRO BUFFD5BWP40
    CLASS CORE ;
    FOREIGN BUFFD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.340000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.155 0.355 1.415 0.465 ;
        RECT  1.155 0.700 1.415 0.820 ;
        RECT  1.105 0.355 1.155 0.820 ;
        RECT  1.085 0.355 1.105 1.045 ;
        RECT  1.015 0.185 1.085 1.045 ;
        RECT  0.945 0.355 1.015 0.820 ;
        RECT  0.695 0.355 0.945 0.465 ;
        RECT  0.695 0.700 0.945 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.385 0.635 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.320 0.280 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.510 -0.115 0.800 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.540 1.375 ;
        RECT  1.200 0.890 1.320 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.890 0.920 1.375 ;
        RECT  0.530 1.145 0.800 1.375 ;
        RECT  0.410 0.905 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.870 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.225 0.355 1.415 0.465 ;
        RECT  1.225 0.700 1.415 0.820 ;
        RECT  0.695 0.355 0.875 0.465 ;
        RECT  0.695 0.700 0.875 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        RECT  0.535 0.545 0.825 0.615 ;
        RECT  0.465 0.345 0.535 0.815 ;
        RECT  0.315 0.345 0.465 0.415 ;
        RECT  0.315 0.745 0.465 0.815 ;
        RECT  0.245 0.245 0.315 0.415 ;
        RECT  0.245 0.745 0.315 1.045 ;
    END
END BUFFD5BWP40

MACRO BUFFD6BWP40
    CLASS CORE ;
    FOREIGN BUFFD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.384000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.155 0.355 1.455 0.465 ;
        RECT  1.155 0.700 1.455 0.820 ;
        RECT  1.145 0.355 1.155 0.820 ;
        RECT  1.125 0.355 1.145 1.045 ;
        RECT  1.055 0.185 1.125 1.045 ;
        RECT  0.945 0.355 1.055 0.820 ;
        RECT  0.725 0.355 0.945 0.465 ;
        RECT  0.725 0.700 0.945 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.765 ;
        RECT  0.165 0.495 0.315 0.635 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.465 ;
        RECT  1.360 -0.115 1.690 0.115 ;
        RECT  1.240 -0.115 1.360 0.280 ;
        RECT  0.960 -0.115 1.240 0.115 ;
        RECT  0.840 -0.115 0.960 0.280 ;
        RECT  0.540 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.540 0.270 ;
        RECT  0.140 -0.115 0.460 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.720 1.770 1.375 ;
        RECT  1.360 1.145 1.690 1.375 ;
        RECT  1.240 0.890 1.360 1.375 ;
        RECT  0.960 1.145 1.240 1.375 ;
        RECT  0.840 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.000 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.730 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.225 0.355 1.455 0.465 ;
        RECT  1.225 0.700 1.455 0.820 ;
        RECT  0.725 0.355 0.875 0.465 ;
        RECT  0.725 0.700 0.875 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  0.565 0.545 0.865 0.615 ;
        RECT  0.485 0.345 0.565 0.915 ;
        RECT  0.325 0.345 0.485 0.415 ;
        RECT  0.325 0.845 0.485 0.915 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.845 0.325 0.995 ;
    END
END BUFFD6BWP40

MACRO BUFFD8BWP40
    CLASS CORE ;
    FOREIGN BUFFD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.512000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.765 0.305 2.055 0.465 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.655 0.185 1.715 0.950 ;
        RECT  1.365 0.305 1.655 0.950 ;
        RECT  1.325 0.305 1.365 0.465 ;
        RECT  0.825 0.720 1.365 0.950 ;
        RECT  1.235 0.185 1.325 0.465 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.300 0.625 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.960 -0.115 2.250 0.115 ;
        RECT  1.840 -0.115 1.960 0.235 ;
        RECT  1.560 -0.115 1.840 0.115 ;
        RECT  1.440 -0.115 1.560 0.235 ;
        RECT  1.160 -0.115 1.440 0.115 ;
        RECT  1.040 -0.115 1.160 0.235 ;
        RECT  0.730 -0.115 1.040 0.115 ;
        RECT  0.650 -0.115 0.730 0.465 ;
        RECT  0.360 -0.115 0.650 0.115 ;
        RECT  0.240 -0.115 0.360 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.145 2.380 1.375 ;
        RECT  2.250 0.700 2.330 1.375 ;
        RECT  1.960 1.145 2.250 1.375 ;
        RECT  1.840 1.020 1.960 1.375 ;
        RECT  1.560 1.145 1.840 1.375 ;
        RECT  1.440 1.020 1.560 1.375 ;
        RECT  1.160 1.145 1.440 1.375 ;
        RECT  1.040 1.020 1.160 1.375 ;
        RECT  0.730 1.145 1.040 1.375 ;
        RECT  0.650 0.700 0.730 1.375 ;
        RECT  0.360 1.145 0.650 1.375 ;
        RECT  0.240 0.910 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.785 0.305 2.055 0.465 ;
        RECT  1.235 0.185 1.295 0.465 ;
        RECT  0.825 0.720 1.295 0.950 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        RECT  0.535 0.545 1.215 0.615 ;
        RECT  0.445 0.185 0.535 1.055 ;
        RECT  0.125 0.335 0.445 0.415 ;
        RECT  0.125 0.750 0.445 0.830 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.750 0.125 1.055 ;
    END
END BUFFD8BWP40

MACRO CKAN2D1BWP40
    CLASS CORE ;
    FOREIGN CKAN2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.700 0.185 0.735 0.315 ;
        RECT  0.705 0.745 0.735 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.490 0.420 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 -0.115 0.840 0.115 ;
        RECT  0.455 -0.115 0.575 0.215 ;
        RECT  0.000 -0.115 0.455 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.840 1.375 ;
        RECT  0.480 0.990 0.600 1.375 ;
        RECT  0.150 1.145 0.480 1.375 ;
        RECT  0.070 0.985 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.605 0.520 0.655 0.640 ;
        RECT  0.535 0.305 0.605 0.915 ;
        RECT  0.165 0.305 0.535 0.375 ;
        RECT  0.340 0.845 0.535 0.915 ;
        RECT  0.260 0.845 0.340 1.050 ;
        RECT  0.070 0.210 0.165 0.375 ;
    END
END CKAN2D1BWP40

MACRO CKAN2D2BWP40
    CLASS CORE ;
    FOREIGN CKAN2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.905 ;
        RECT  0.715 0.355 0.735 0.475 ;
        RECT  0.715 0.765 0.735 0.905 ;
        RECT  0.645 0.185 0.715 0.475 ;
        RECT  0.645 0.765 0.715 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.024400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.395 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.024400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.280 ;
        RECT  0.550 -0.115 0.830 0.115 ;
        RECT  0.410 -0.115 0.550 0.210 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.420 0.985 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.895 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 0.545 0.640 0.615 ;
        RECT  0.470 0.290 0.540 0.915 ;
        RECT  0.035 0.290 0.470 0.360 ;
        RECT  0.340 0.845 0.470 0.915 ;
        RECT  0.220 0.845 0.340 1.055 ;
    END
END CKAN2D2BWP40

MACRO CKAN2D4BWP40
    CLASS CORE ;
    FOREIGN CKAN2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.185 1.515 0.485 ;
        RECT  1.445 0.700 1.515 1.030 ;
        RECT  1.435 0.355 1.445 0.485 ;
        RECT  1.435 0.700 1.445 0.820 ;
        RECT  1.225 0.355 1.435 0.820 ;
        RECT  1.135 0.355 1.225 0.475 ;
        RECT  1.135 0.700 1.225 0.820 ;
        RECT  1.065 0.185 1.135 0.475 ;
        RECT  1.065 0.700 1.135 1.030 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.048800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.780 0.640 ;
        RECT  0.625 0.520 0.695 0.790 ;
        RECT  0.245 0.720 0.625 0.790 ;
        RECT  0.170 0.495 0.245 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.048800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.480 0.545 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.730 -0.115 1.820 0.115 ;
        RECT  1.650 -0.115 1.730 0.475 ;
        RECT  1.350 -0.115 1.650 0.115 ;
        RECT  1.230 -0.115 1.350 0.280 ;
        RECT  0.940 -0.115 1.230 0.115 ;
        RECT  0.820 -0.115 0.940 0.215 ;
        RECT  0.130 -0.115 0.820 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 1.145 1.820 1.375 ;
        RECT  1.655 0.720 1.735 1.375 ;
        RECT  1.350 1.145 1.655 1.375 ;
        RECT  1.230 0.890 1.350 1.375 ;
        RECT  0.920 1.145 1.230 1.375 ;
        RECT  0.840 1.000 0.920 1.375 ;
        RECT  0.510 1.145 0.840 1.375 ;
        RECT  0.430 1.000 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.185 1.515 0.485 ;
        RECT  1.505 0.700 1.515 1.030 ;
        RECT  1.135 0.355 1.155 0.475 ;
        RECT  1.135 0.700 1.155 0.820 ;
        RECT  1.065 0.185 1.135 0.475 ;
        RECT  1.065 0.700 1.135 1.030 ;
        RECT  0.925 0.545 1.145 0.615 ;
        RECT  0.855 0.335 0.925 0.930 ;
        RECT  0.410 0.335 0.855 0.405 ;
        RECT  0.720 0.860 0.855 0.930 ;
        RECT  0.220 0.195 0.720 0.265 ;
        RECT  0.600 0.860 0.720 1.065 ;
        RECT  0.340 0.860 0.600 0.930 ;
        RECT  0.220 0.860 0.340 1.065 ;
    END
END CKAN2D4BWP40

MACRO CKAN2D8BWP40
    CLASS CORE ;
    FOREIGN CKAN2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.135 0.325 2.220 0.445 ;
        RECT  2.135 0.700 2.220 0.820 ;
        RECT  1.925 0.325 2.135 0.820 ;
        RECT  1.900 0.325 1.925 0.445 ;
        RECT  1.900 0.700 1.925 0.820 ;
        RECT  1.805 0.185 1.900 0.445 ;
        RECT  1.805 0.700 1.900 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.072800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.160 0.770 ;
        RECT  0.535 0.700 1.015 0.770 ;
        RECT  0.445 0.495 0.535 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.072800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.545 0.915 0.625 ;
        RECT  0.730 0.350 0.815 0.625 ;
        RECT  0.275 0.350 0.730 0.420 ;
        RECT  0.195 0.350 0.275 0.640 ;
        RECT  0.125 0.495 0.195 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.445 ;
        RECT  2.520 -0.115 2.810 0.115 ;
        RECT  2.400 -0.115 2.520 0.255 ;
        RECT  2.120 -0.115 2.400 0.115 ;
        RECT  2.000 -0.115 2.120 0.255 ;
        RECT  1.720 -0.115 2.000 0.115 ;
        RECT  1.600 -0.115 1.720 0.255 ;
        RECT  1.300 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.300 0.265 ;
        RECT  0.540 -0.115 1.220 0.115 ;
        RECT  0.420 -0.115 0.540 0.140 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.720 2.890 1.375 ;
        RECT  2.520 1.145 2.810 1.375 ;
        RECT  2.400 0.890 2.520 1.375 ;
        RECT  2.120 1.145 2.400 1.375 ;
        RECT  2.000 0.890 2.120 1.375 ;
        RECT  1.720 1.145 2.000 1.375 ;
        RECT  1.600 0.890 1.720 1.375 ;
        RECT  1.300 1.145 1.600 1.375 ;
        RECT  1.220 0.980 1.300 1.375 ;
        RECT  0.910 1.145 1.220 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.520 1.145 0.830 1.375 ;
        RECT  0.440 0.980 0.520 1.375 ;
        RECT  0.130 1.145 0.440 1.375 ;
        RECT  0.050 0.895 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.205 0.325 2.220 0.445 ;
        RECT  2.205 0.700 2.220 0.820 ;
        RECT  1.805 0.185 1.855 0.445 ;
        RECT  1.805 0.700 1.855 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        RECT  1.320 0.545 1.775 0.615 ;
        RECT  0.740 0.840 1.000 0.910 ;
        RECT  0.620 0.840 0.740 1.050 ;
        RECT  0.315 0.840 0.620 0.910 ;
        RECT  0.245 0.840 0.315 1.035 ;
        RECT  0.055 0.210 0.125 0.380 ;
        RECT  1.250 0.345 1.320 0.910 ;
        RECT  1.095 0.345 1.250 0.415 ;
        RECT  1.120 0.840 1.250 0.910 ;
        RECT  1.000 0.840 1.120 1.050 ;
        RECT  1.025 0.210 1.095 0.415 ;
        RECT  0.125 0.210 1.025 0.280 ;
    END
END CKAN2D8BWP40

MACRO CKBD10BWP40
    CLASS CORE ;
    FOREIGN CKBD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.600000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  1.995 0.305 2.195 0.465 ;
        RECT  1.885 0.305 1.995 0.950 ;
        RECT  1.815 0.185 1.885 0.950 ;
        RECT  1.785 0.305 1.815 0.950 ;
        RECT  1.505 0.305 1.785 0.465 ;
        RECT  1.030 0.720 1.785 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 2.940 0.115 ;
        RECT  2.760 -0.115 2.840 0.465 ;
        RECT  2.480 -0.115 2.760 0.115 ;
        RECT  2.360 -0.115 2.480 0.235 ;
        RECT  2.100 -0.115 2.360 0.115 ;
        RECT  1.980 -0.115 2.100 0.235 ;
        RECT  1.720 -0.115 1.980 0.115 ;
        RECT  1.600 -0.115 1.720 0.235 ;
        RECT  1.340 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.340 0.235 ;
        RECT  0.940 -0.115 1.220 0.115 ;
        RECT  0.860 -0.115 0.940 0.465 ;
        RECT  0.565 -0.115 0.860 0.115 ;
        RECT  0.475 -0.115 0.565 0.260 ;
        RECT  0.190 -0.115 0.475 0.115 ;
        RECT  0.090 -0.115 0.190 0.410 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.145 2.940 1.375 ;
        RECT  2.760 0.700 2.840 1.375 ;
        RECT  2.480 1.145 2.760 1.375 ;
        RECT  2.360 1.020 2.480 1.375 ;
        RECT  2.100 1.145 2.360 1.375 ;
        RECT  1.980 1.020 2.100 1.375 ;
        RECT  1.720 1.145 1.980 1.375 ;
        RECT  1.600 1.020 1.720 1.375 ;
        RECT  1.340 1.145 1.600 1.375 ;
        RECT  1.220 1.020 1.340 1.375 ;
        RECT  0.940 1.145 1.220 1.375 ;
        RECT  0.860 0.720 0.940 1.375 ;
        RECT  0.560 1.145 0.860 1.375 ;
        RECT  0.480 0.995 0.560 1.375 ;
        RECT  0.190 1.145 0.480 1.375 ;
        RECT  0.090 0.845 0.190 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.065 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  2.065 0.305 2.195 0.465 ;
        RECT  1.505 0.305 1.715 0.465 ;
        RECT  1.030 0.720 1.715 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  0.770 0.545 1.705 0.615 ;
        RECT  0.660 0.195 0.770 1.050 ;
        RECT  0.390 0.335 0.660 0.415 ;
        RECT  0.365 0.770 0.660 0.850 ;
        RECT  0.270 0.205 0.390 0.415 ;
        RECT  0.295 0.770 0.365 1.050 ;
    END
END CKBD10BWP40

MACRO CKBD12BWP40
    CLASS CORE ;
    FOREIGN CKBD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.275 0.305 2.525 0.465 ;
        RECT  2.215 0.305 2.275 0.950 ;
        RECT  2.135 0.185 2.215 0.950 ;
        RECT  1.925 0.305 2.135 0.950 ;
        RECT  1.835 0.305 1.925 0.465 ;
        RECT  0.980 0.720 1.925 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.123200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.465 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.235 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.235 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.890 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.890 0.465 ;
        RECT  0.515 -0.115 0.810 0.115 ;
        RECT  0.425 -0.115 0.515 0.260 ;
        RECT  0.140 -0.115 0.425 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.700 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 1.020 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 1.020 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 1.020 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.020 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 1.020 1.290 1.375 ;
        RECT  0.890 1.145 1.170 1.375 ;
        RECT  0.810 0.720 0.890 1.375 ;
        RECT  0.530 1.145 0.810 1.375 ;
        RECT  0.410 0.910 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.345 0.305 2.525 0.465 ;
        RECT  1.835 0.305 1.855 0.465 ;
        RECT  0.980 0.720 1.855 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  0.720 0.545 1.765 0.615 ;
        RECT  0.610 0.195 0.720 1.050 ;
        RECT  0.340 0.335 0.610 0.415 ;
        RECT  0.315 0.750 0.610 0.830 ;
        RECT  0.220 0.205 0.340 0.415 ;
        RECT  0.245 0.750 0.315 1.050 ;
    END
END CKBD12BWP40

MACRO CKBD14BWP40
    CLASS CORE ;
    FOREIGN CKBD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.872000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.835 0.305 3.125 0.465 ;
        RECT  2.815 0.305 2.835 0.945 ;
        RECT  2.745 0.185 2.815 0.945 ;
        RECT  2.485 0.305 2.745 0.945 ;
        RECT  2.435 0.305 2.485 0.465 ;
        RECT  1.200 0.715 2.485 0.945 ;
        RECT  2.365 0.185 2.435 0.465 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.156000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.665 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 -0.115 3.920 0.115 ;
        RECT  3.730 -0.115 3.835 0.465 ;
        RECT  3.410 -0.115 3.730 0.115 ;
        RECT  3.290 -0.115 3.410 0.235 ;
        RECT  3.030 -0.115 3.290 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.650 -0.115 2.910 0.115 ;
        RECT  2.530 -0.115 2.650 0.235 ;
        RECT  2.270 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.270 0.235 ;
        RECT  1.890 -0.115 2.150 0.115 ;
        RECT  1.770 -0.115 1.890 0.235 ;
        RECT  1.510 -0.115 1.770 0.115 ;
        RECT  1.390 -0.115 1.510 0.235 ;
        RECT  1.100 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.100 0.465 ;
        RECT  0.720 -0.115 1.020 0.115 ;
        RECT  0.600 -0.115 0.720 0.265 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.835 1.145 3.920 1.375 ;
        RECT  3.730 0.690 3.835 1.375 ;
        RECT  3.410 1.145 3.730 1.375 ;
        RECT  3.290 1.015 3.410 1.375 ;
        RECT  3.030 1.145 3.290 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.650 1.145 2.910 1.375 ;
        RECT  2.530 1.015 2.650 1.375 ;
        RECT  2.270 1.145 2.530 1.375 ;
        RECT  2.150 1.015 2.270 1.375 ;
        RECT  1.890 1.145 2.150 1.375 ;
        RECT  1.770 1.015 1.890 1.375 ;
        RECT  1.510 1.145 1.770 1.375 ;
        RECT  1.390 1.015 1.510 1.375 ;
        RECT  1.120 1.145 1.390 1.375 ;
        RECT  1.000 0.710 1.120 1.375 ;
        RECT  0.700 1.145 1.000 1.375 ;
        RECT  0.620 1.000 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 1.000 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.905 0.305 3.125 0.465 ;
        RECT  2.365 0.185 2.415 0.465 ;
        RECT  1.200 0.715 2.415 0.945 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        RECT  0.920 0.545 2.405 0.615 ;
        RECT  0.790 0.195 0.920 1.065 ;
        RECT  0.510 0.335 0.790 0.415 ;
        RECT  0.525 0.845 0.790 0.915 ;
        RECT  0.415 0.845 0.525 1.075 ;
        RECT  0.430 0.185 0.510 0.415 ;
        RECT  0.130 0.335 0.430 0.415 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.255 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.075 ;
    END
END CKBD14BWP40

MACRO CKBD16BWP40
    CLASS CORE ;
    FOREIGN CKBD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.115 0.305 3.405 0.465 ;
        RECT  3.095 0.305 3.115 0.945 ;
        RECT  3.025 0.185 3.095 0.945 ;
        RECT  2.765 0.305 3.025 0.945 ;
        RECT  2.715 0.305 2.765 0.465 ;
        RECT  1.480 0.715 2.765 0.945 ;
        RECT  2.645 0.185 2.715 0.465 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.184800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.945 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.115 4.480 0.115 ;
        RECT  4.350 -0.115 4.430 0.465 ;
        RECT  4.070 -0.115 4.350 0.115 ;
        RECT  3.950 -0.115 4.070 0.235 ;
        RECT  3.690 -0.115 3.950 0.115 ;
        RECT  3.570 -0.115 3.690 0.235 ;
        RECT  3.310 -0.115 3.570 0.115 ;
        RECT  3.190 -0.115 3.310 0.235 ;
        RECT  2.930 -0.115 3.190 0.115 ;
        RECT  2.810 -0.115 2.930 0.235 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.235 ;
        RECT  2.170 -0.115 2.430 0.115 ;
        RECT  2.050 -0.115 2.170 0.235 ;
        RECT  1.790 -0.115 2.050 0.115 ;
        RECT  1.670 -0.115 1.790 0.235 ;
        RECT  1.380 -0.115 1.670 0.115 ;
        RECT  1.300 -0.115 1.380 0.465 ;
        RECT  1.000 -0.115 1.300 0.115 ;
        RECT  0.880 -0.115 1.000 0.265 ;
        RECT  0.620 -0.115 0.880 0.115 ;
        RECT  0.500 -0.115 0.620 0.265 ;
        RECT  0.180 -0.115 0.500 0.115 ;
        RECT  0.060 -0.115 0.180 0.415 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.145 4.480 1.375 ;
        RECT  4.350 0.690 4.430 1.375 ;
        RECT  4.070 1.145 4.350 1.375 ;
        RECT  3.950 1.015 4.070 1.375 ;
        RECT  3.690 1.145 3.950 1.375 ;
        RECT  3.570 1.015 3.690 1.375 ;
        RECT  3.310 1.145 3.570 1.375 ;
        RECT  3.190 1.015 3.310 1.375 ;
        RECT  2.930 1.145 3.190 1.375 ;
        RECT  2.810 1.015 2.930 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 1.015 2.550 1.375 ;
        RECT  2.170 1.145 2.430 1.375 ;
        RECT  2.050 1.015 2.170 1.375 ;
        RECT  1.790 1.145 2.050 1.375 ;
        RECT  1.670 1.015 1.790 1.375 ;
        RECT  1.400 1.145 1.670 1.375 ;
        RECT  1.280 0.710 1.400 1.375 ;
        RECT  0.980 1.145 1.280 1.375 ;
        RECT  0.900 0.860 0.980 1.375 ;
        RECT  0.600 1.145 0.900 1.375 ;
        RECT  0.520 0.860 0.600 1.375 ;
        RECT  0.170 1.145 0.520 1.375 ;
        RECT  0.090 0.845 0.170 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.185 0.305 3.405 0.465 ;
        RECT  2.645 0.185 2.695 0.465 ;
        RECT  1.480 0.715 2.695 0.945 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        RECT  1.200 0.545 2.685 0.615 ;
        RECT  1.070 0.195 1.200 1.065 ;
        RECT  0.790 0.335 1.070 0.415 ;
        RECT  0.785 0.705 1.070 0.785 ;
        RECT  0.710 0.185 0.790 0.415 ;
        RECT  0.715 0.705 0.785 1.035 ;
        RECT  0.405 0.705 0.715 0.785 ;
        RECT  0.410 0.335 0.710 0.415 ;
        RECT  0.310 0.185 0.410 0.415 ;
        RECT  0.335 0.705 0.405 1.035 ;
    END
END CKBD16BWP40

MACRO CKBD18BWP40
    CLASS CORE ;
    FOREIGN CKBD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.080000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.105 0.305 3.305 0.465 ;
        RECT  2.995 0.305 3.105 0.945 ;
        RECT  2.925 0.185 2.995 0.945 ;
        RECT  2.765 0.305 2.925 0.945 ;
        RECT  2.615 0.305 2.765 0.465 ;
        RECT  1.380 0.715 2.765 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  1.405 0.185 1.475 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.184800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.855 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.350 -0.115 4.630 0.115 ;
        RECT  4.230 -0.115 4.350 0.235 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.235 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.235 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.235 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.235 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.235 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.235 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.235 ;
        RECT  1.280 -0.115 1.570 0.115 ;
        RECT  1.200 -0.115 1.280 0.465 ;
        RECT  0.910 -0.115 1.200 0.115 ;
        RECT  0.790 -0.115 0.910 0.265 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.265 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.630 0.690 4.710 1.375 ;
        RECT  4.350 1.145 4.630 1.375 ;
        RECT  4.230 1.015 4.350 1.375 ;
        RECT  3.970 1.145 4.230 1.375 ;
        RECT  3.850 1.015 3.970 1.375 ;
        RECT  3.590 1.145 3.850 1.375 ;
        RECT  3.470 1.015 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.090 1.015 3.210 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.015 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.330 1.015 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 1.015 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.570 1.015 1.690 1.375 ;
        RECT  1.300 1.145 1.570 1.375 ;
        RECT  1.180 0.710 1.300 1.375 ;
        RECT  0.890 1.145 1.180 1.375 ;
        RECT  0.810 0.860 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.860 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.185 0.305 3.305 0.465 ;
        RECT  2.615 0.305 2.695 0.465 ;
        RECT  1.380 0.715 2.695 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.110 0.545 2.585 0.615 ;
        RECT  0.980 0.195 1.110 1.065 ;
        RECT  0.700 0.335 0.980 0.415 ;
        RECT  0.695 0.705 0.980 0.785 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.625 0.705 0.695 1.035 ;
        RECT  0.315 0.705 0.625 0.785 ;
        RECT  0.320 0.335 0.620 0.415 ;
        RECT  0.220 0.185 0.320 0.415 ;
        RECT  0.245 0.705 0.315 1.035 ;
    END
END CKBD18BWP40

MACRO CKBD1BWP40
    CLASS CORE ;
    FOREIGN CKBD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.185 0.525 1.045 ;
        RECT  0.435 0.185 0.455 0.465 ;
        RECT  0.435 0.735 0.455 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.190 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.365 0.520 0.385 0.640 ;
        RECT  0.295 0.335 0.365 0.925 ;
        RECT  0.130 0.335 0.295 0.405 ;
        RECT  0.130 0.855 0.295 0.925 ;
        RECT  0.050 0.195 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END CKBD1BWP40

MACRO CKBD20BWP40
    CLASS CORE ;
    FOREIGN CKBD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.200000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.555 0.305 3.865 0.465 ;
        RECT  3.535 0.185 3.555 0.465 ;
        RECT  3.485 0.185 3.535 0.960 ;
        RECT  3.185 0.305 3.485 0.960 ;
        RECT  3.175 0.305 3.185 0.465 ;
        RECT  1.560 0.730 3.185 0.960 ;
        RECT  3.105 0.185 3.175 0.465 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.224000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.065 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 -0.115 5.320 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.910 -0.115 5.190 0.115 ;
        RECT  4.790 -0.115 4.910 0.235 ;
        RECT  4.530 -0.115 4.790 0.115 ;
        RECT  4.410 -0.115 4.530 0.235 ;
        RECT  4.150 -0.115 4.410 0.115 ;
        RECT  4.030 -0.115 4.150 0.235 ;
        RECT  3.770 -0.115 4.030 0.115 ;
        RECT  3.650 -0.115 3.770 0.235 ;
        RECT  3.390 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.010 -0.115 3.270 0.115 ;
        RECT  2.890 -0.115 3.010 0.235 ;
        RECT  2.630 -0.115 2.890 0.115 ;
        RECT  2.510 -0.115 2.630 0.235 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.235 ;
        RECT  1.870 -0.115 2.130 0.115 ;
        RECT  1.750 -0.115 1.870 0.235 ;
        RECT  1.465 -0.115 1.750 0.115 ;
        RECT  1.395 -0.115 1.465 0.465 ;
        RECT  1.085 -0.115 1.395 0.115 ;
        RECT  1.015 -0.115 1.085 0.255 ;
        RECT  0.695 -0.115 1.015 0.115 ;
        RECT  0.625 -0.115 0.695 0.255 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.245 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.270 1.145 5.320 1.375 ;
        RECT  5.190 0.700 5.270 1.375 ;
        RECT  4.910 1.145 5.190 1.375 ;
        RECT  4.790 1.030 4.910 1.375 ;
        RECT  4.530 1.145 4.790 1.375 ;
        RECT  4.410 1.030 4.530 1.375 ;
        RECT  4.150 1.145 4.410 1.375 ;
        RECT  4.030 1.030 4.150 1.375 ;
        RECT  3.770 1.145 4.030 1.375 ;
        RECT  3.650 1.030 3.770 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.030 3.390 1.375 ;
        RECT  3.010 1.145 3.270 1.375 ;
        RECT  2.890 1.030 3.010 1.375 ;
        RECT  2.630 1.145 2.890 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.250 1.145 2.510 1.375 ;
        RECT  2.130 1.030 2.250 1.375 ;
        RECT  1.870 1.145 2.130 1.375 ;
        RECT  1.750 1.030 1.870 1.375 ;
        RECT  1.465 1.145 1.750 1.375 ;
        RECT  1.395 0.720 1.465 1.375 ;
        RECT  1.085 1.145 1.395 1.375 ;
        RECT  1.015 1.005 1.085 1.375 ;
        RECT  0.710 1.145 1.015 1.375 ;
        RECT  0.610 1.015 0.710 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.230 1.015 0.330 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.605 0.305 3.865 0.465 ;
        RECT  3.105 0.185 3.115 0.465 ;
        RECT  1.560 0.730 3.115 0.960 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        RECT  1.315 0.545 3.105 0.615 ;
        RECT  1.155 0.185 1.315 1.065 ;
        RECT  0.895 0.335 1.155 0.415 ;
        RECT  0.920 0.845 1.155 0.925 ;
        RECT  0.800 0.845 0.920 1.065 ;
        RECT  0.825 0.185 0.895 0.415 ;
        RECT  0.505 0.335 0.825 0.415 ;
        RECT  0.530 0.845 0.800 0.925 ;
        RECT  0.410 0.845 0.530 1.075 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.130 0.335 0.435 0.415 ;
        RECT  0.125 0.845 0.410 0.920 ;
        RECT  0.055 0.275 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.075 ;
    END
END CKBD20BWP40

MACRO CKBD24BWP40
    CLASS CORE ;
    FOREIGN CKBD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.440000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.155 0.305 4.465 0.465 ;
        RECT  4.095 0.185 4.155 0.465 ;
        RECT  4.085 0.185 4.095 0.945 ;
        RECT  3.775 0.305 4.085 0.945 ;
        RECT  3.745 0.185 3.775 0.945 ;
        RECT  3.705 0.185 3.745 0.465 ;
        RECT  1.780 0.715 3.745 0.945 ;
        RECT  3.395 0.305 3.705 0.465 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.246400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.155 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.170 -0.115 6.250 0.475 ;
        RECT  5.890 -0.115 6.170 0.115 ;
        RECT  5.770 -0.115 5.890 0.235 ;
        RECT  5.510 -0.115 5.770 0.115 ;
        RECT  5.390 -0.115 5.510 0.235 ;
        RECT  5.130 -0.115 5.390 0.115 ;
        RECT  5.010 -0.115 5.130 0.235 ;
        RECT  4.750 -0.115 5.010 0.115 ;
        RECT  4.630 -0.115 4.750 0.235 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.235 ;
        RECT  3.990 -0.115 4.250 0.115 ;
        RECT  3.870 -0.115 3.990 0.235 ;
        RECT  3.610 -0.115 3.870 0.115 ;
        RECT  3.490 -0.115 3.610 0.235 ;
        RECT  3.230 -0.115 3.490 0.115 ;
        RECT  3.110 -0.115 3.230 0.235 ;
        RECT  2.850 -0.115 3.110 0.115 ;
        RECT  2.730 -0.115 2.850 0.235 ;
        RECT  2.470 -0.115 2.730 0.115 ;
        RECT  2.350 -0.115 2.470 0.235 ;
        RECT  2.090 -0.115 2.350 0.115 ;
        RECT  1.970 -0.115 2.090 0.235 ;
        RECT  1.685 -0.115 1.970 0.115 ;
        RECT  1.615 -0.115 1.685 0.465 ;
        RECT  1.295 -0.115 1.615 0.115 ;
        RECT  1.225 -0.115 1.295 0.245 ;
        RECT  0.895 -0.115 1.225 0.115 ;
        RECT  0.825 -0.115 0.895 0.245 ;
        RECT  0.505 -0.115 0.825 0.115 ;
        RECT  0.435 -0.115 0.505 0.245 ;
        RECT  0.125 -0.115 0.435 0.115 ;
        RECT  0.055 -0.115 0.125 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.170 0.720 6.250 1.375 ;
        RECT  5.890 1.145 6.170 1.375 ;
        RECT  5.770 1.015 5.890 1.375 ;
        RECT  5.510 1.145 5.770 1.375 ;
        RECT  5.390 1.015 5.510 1.375 ;
        RECT  5.130 1.145 5.390 1.375 ;
        RECT  5.010 1.015 5.130 1.375 ;
        RECT  4.750 1.145 5.010 1.375 ;
        RECT  4.630 1.015 4.750 1.375 ;
        RECT  4.370 1.145 4.630 1.375 ;
        RECT  4.250 1.015 4.370 1.375 ;
        RECT  3.990 1.145 4.250 1.375 ;
        RECT  3.870 1.015 3.990 1.375 ;
        RECT  3.610 1.145 3.870 1.375 ;
        RECT  3.490 1.015 3.610 1.375 ;
        RECT  3.230 1.145 3.490 1.375 ;
        RECT  3.110 1.015 3.230 1.375 ;
        RECT  2.850 1.145 3.110 1.375 ;
        RECT  2.730 1.015 2.850 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 1.015 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 1.015 2.090 1.375 ;
        RECT  1.685 1.145 1.970 1.375 ;
        RECT  1.615 0.740 1.685 1.375 ;
        RECT  1.295 1.145 1.615 1.375 ;
        RECT  1.225 0.880 1.295 1.375 ;
        RECT  0.900 1.145 1.225 1.375 ;
        RECT  0.820 0.880 0.900 1.375 ;
        RECT  0.510 1.145 0.820 1.375 ;
        RECT  0.430 0.880 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.165 0.305 4.465 0.465 ;
        RECT  3.395 0.305 3.675 0.465 ;
        RECT  1.780 0.715 3.675 0.945 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        RECT  1.535 0.545 3.645 0.615 ;
        RECT  1.365 0.195 1.535 1.070 ;
        RECT  1.100 0.325 1.365 0.415 ;
        RECT  1.120 0.705 1.365 0.795 ;
        RECT  1.000 0.705 1.120 1.070 ;
        RECT  1.020 0.185 1.100 0.415 ;
        RECT  0.700 0.325 1.020 0.415 ;
        RECT  0.720 0.705 1.000 0.795 ;
        RECT  0.600 0.705 0.720 1.070 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.320 0.325 0.620 0.415 ;
        RECT  0.340 0.705 0.600 0.795 ;
        RECT  0.220 0.705 0.340 1.065 ;
        RECT  0.220 0.185 0.320 0.415 ;
    END
END CKBD24BWP40

MACRO CKBD2BWP40
    CLASS CORE ;
    FOREIGN CKBD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.152000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.385 0.805 0.875 ;
        RECT  0.555 0.385 0.735 0.455 ;
        RECT  0.555 0.775 0.735 0.875 ;
        RECT  0.465 0.185 0.555 0.455 ;
        RECT  0.465 0.775 0.555 1.065 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.245 0.640 ;
        RECT  0.035 0.485 0.105 0.775 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 -0.115 0.840 0.115 ;
        RECT  0.660 -0.115 0.780 0.265 ;
        RECT  0.340 -0.115 0.660 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.145 0.840 1.375 ;
        RECT  0.660 0.995 0.780 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.220 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.395 0.545 0.535 0.615 ;
        RECT  0.325 0.335 0.395 0.925 ;
        RECT  0.130 0.335 0.325 0.405 ;
        RECT  0.130 0.855 0.325 0.925 ;
        RECT  0.050 0.195 0.130 0.405 ;
        RECT  0.050 0.855 0.130 1.045 ;
    END
END CKBD2BWP40

MACRO CKBD3BWP40
    CLASS CORE ;
    FOREIGN CKBD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.185 0.945 0.490 ;
        RECT  0.875 0.700 0.945 1.045 ;
        RECT  0.855 0.185 0.875 1.045 ;
        RECT  0.665 0.355 0.855 0.820 ;
        RECT  0.545 0.355 0.665 0.475 ;
        RECT  0.545 0.700 0.665 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.280 ;
        RECT  0.360 -0.115 0.640 0.115 ;
        RECT  0.240 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 0.890 0.760 1.375 ;
        RECT  0.360 1.145 0.640 1.375 ;
        RECT  0.240 1.040 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.545 0.355 0.595 0.475 ;
        RECT  0.545 0.700 0.595 0.820 ;
        RECT  0.475 0.185 0.545 0.475 ;
        RECT  0.475 0.700 0.545 1.045 ;
        RECT  0.395 0.545 0.575 0.615 ;
        RECT  0.325 0.345 0.395 0.970 ;
        RECT  0.130 0.345 0.325 0.415 ;
        RECT  0.130 0.900 0.325 0.970 ;
        RECT  0.050 0.245 0.130 0.415 ;
        RECT  0.050 0.900 0.130 1.030 ;
    END
END CKBD3BWP40

MACRO CKBD4BWP40
    CLASS CORE ;
    FOREIGN CKBD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  1.055 0.700 1.125 1.045 ;
        RECT  1.015 0.355 1.055 0.465 ;
        RECT  1.015 0.700 1.055 0.820 ;
        RECT  0.805 0.355 1.015 0.820 ;
        RECT  0.725 0.355 0.805 0.465 ;
        RECT  0.725 0.700 0.805 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.280 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.475 ;
        RECT  0.950 -0.115 1.270 0.115 ;
        RECT  0.830 -0.115 0.950 0.280 ;
        RECT  0.530 -0.115 0.830 0.115 ;
        RECT  0.450 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.450 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.270 0.700 1.350 1.375 ;
        RECT  0.950 1.145 1.270 1.375 ;
        RECT  0.830 0.890 0.950 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.440 0.975 0.540 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.185 1.125 0.465 ;
        RECT  1.085 0.700 1.125 1.045 ;
        RECT  0.725 0.355 0.735 0.465 ;
        RECT  0.725 0.700 0.735 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  0.585 0.545 0.720 0.615 ;
        RECT  0.510 0.345 0.585 0.905 ;
        RECT  0.325 0.345 0.510 0.415 ;
        RECT  0.325 0.835 0.510 0.905 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.835 0.325 0.995 ;
    END
END CKBD4BWP40

MACRO CKBD5BWP40
    CLASS CORE ;
    FOREIGN CKBD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.340000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.155 0.355 1.415 0.465 ;
        RECT  1.155 0.700 1.415 0.820 ;
        RECT  1.105 0.355 1.155 0.820 ;
        RECT  1.085 0.355 1.105 1.045 ;
        RECT  1.015 0.185 1.085 1.045 ;
        RECT  0.945 0.355 1.015 0.820 ;
        RECT  0.695 0.355 0.945 0.465 ;
        RECT  0.695 0.700 0.945 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.063200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.385 0.635 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.320 0.280 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.510 -0.115 0.800 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.540 1.375 ;
        RECT  1.200 0.890 1.320 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.890 0.920 1.375 ;
        RECT  0.530 1.145 0.800 1.375 ;
        RECT  0.410 0.890 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.860 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.225 0.355 1.415 0.465 ;
        RECT  1.225 0.700 1.415 0.820 ;
        RECT  0.695 0.355 0.875 0.465 ;
        RECT  0.695 0.700 0.875 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        RECT  0.535 0.545 0.825 0.615 ;
        RECT  0.465 0.345 0.535 0.820 ;
        RECT  0.315 0.345 0.465 0.415 ;
        RECT  0.315 0.750 0.465 0.820 ;
        RECT  0.245 0.245 0.315 0.415 ;
        RECT  0.245 0.750 0.315 0.995 ;
    END
END CKBD5BWP40

MACRO CKBD6BWP40
    CLASS CORE ;
    FOREIGN CKBD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.384000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.155 0.355 1.455 0.465 ;
        RECT  1.155 0.700 1.455 0.820 ;
        RECT  1.145 0.355 1.155 0.820 ;
        RECT  1.125 0.355 1.145 1.045 ;
        RECT  1.055 0.185 1.125 1.045 ;
        RECT  0.945 0.355 1.055 0.820 ;
        RECT  0.725 0.355 0.945 0.465 ;
        RECT  0.725 0.700 0.945 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.385 0.635 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.465 ;
        RECT  1.360 -0.115 1.690 0.115 ;
        RECT  1.240 -0.115 1.360 0.280 ;
        RECT  0.960 -0.115 1.240 0.115 ;
        RECT  0.840 -0.115 0.960 0.280 ;
        RECT  0.540 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.540 0.270 ;
        RECT  0.140 -0.115 0.460 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.735 1.770 1.375 ;
        RECT  1.360 1.145 1.690 1.375 ;
        RECT  1.240 0.890 1.360 1.375 ;
        RECT  0.960 1.145 1.240 1.375 ;
        RECT  0.840 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.000 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.225 0.355 1.455 0.465 ;
        RECT  1.225 0.700 1.455 0.820 ;
        RECT  0.725 0.355 0.875 0.465 ;
        RECT  0.725 0.700 0.875 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  0.565 0.545 0.865 0.615 ;
        RECT  0.485 0.345 0.565 0.915 ;
        RECT  0.325 0.345 0.485 0.415 ;
        RECT  0.325 0.845 0.485 0.915 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.845 0.325 0.995 ;
    END
END CKBD6BWP40

MACRO CKBD8BWP40
    CLASS CORE ;
    FOREIGN CKBD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.512000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.765 0.305 2.055 0.465 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.655 0.185 1.715 0.950 ;
        RECT  1.365 0.305 1.655 0.950 ;
        RECT  1.325 0.305 1.365 0.465 ;
        RECT  0.825 0.720 1.365 0.950 ;
        RECT  1.235 0.185 1.325 0.465 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.092400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.300 0.625 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.115 2.380 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.960 -0.115 2.250 0.115 ;
        RECT  1.840 -0.115 1.960 0.235 ;
        RECT  1.560 -0.115 1.840 0.115 ;
        RECT  1.440 -0.115 1.560 0.235 ;
        RECT  1.160 -0.115 1.440 0.115 ;
        RECT  1.040 -0.115 1.160 0.235 ;
        RECT  0.730 -0.115 1.040 0.115 ;
        RECT  0.650 -0.115 0.730 0.465 ;
        RECT  0.360 -0.115 0.650 0.115 ;
        RECT  0.240 -0.115 0.360 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.145 2.380 1.375 ;
        RECT  2.250 0.700 2.330 1.375 ;
        RECT  1.960 1.145 2.250 1.375 ;
        RECT  1.840 1.020 1.960 1.375 ;
        RECT  1.560 1.145 1.840 1.375 ;
        RECT  1.440 1.020 1.560 1.375 ;
        RECT  1.160 1.145 1.440 1.375 ;
        RECT  1.040 1.020 1.160 1.375 ;
        RECT  0.730 1.145 1.040 1.375 ;
        RECT  0.650 0.700 0.730 1.375 ;
        RECT  0.360 1.145 0.650 1.375 ;
        RECT  0.240 1.015 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.785 0.305 2.055 0.465 ;
        RECT  1.235 0.185 1.295 0.465 ;
        RECT  0.825 0.720 1.295 0.950 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        RECT  0.535 0.545 1.215 0.615 ;
        RECT  0.445 0.185 0.535 1.055 ;
        RECT  0.125 0.335 0.445 0.415 ;
        RECT  0.125 0.850 0.445 0.930 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.850 0.125 1.035 ;
    END
END CKBD8BWP40

MACRO CKLHQD10BWP40
    CLASS CORE ;
    FOREIGN CKLHQD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.600000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.375 0.185 7.465 0.435 ;
        RECT  7.380 0.745 7.465 1.045 ;
        RECT  7.100 0.745 7.380 0.815 ;
        RECT  7.085 0.355 7.375 0.435 ;
        RECT  7.000 0.745 7.100 1.045 ;
        RECT  7.000 0.185 7.085 0.435 ;
        RECT  6.755 0.355 7.000 0.435 ;
        RECT  6.755 0.745 7.000 0.815 ;
        RECT  6.695 0.355 6.755 0.815 ;
        RECT  6.615 0.185 6.695 1.045 ;
        RECT  6.545 0.355 6.615 0.815 ;
        RECT  6.315 0.355 6.545 0.435 ;
        RECT  6.315 0.745 6.545 0.815 ;
        RECT  6.240 0.185 6.315 0.435 ;
        RECT  6.245 0.745 6.315 1.045 ;
        RECT  5.955 0.745 6.245 0.815 ;
        RECT  5.955 0.355 6.240 0.435 ;
        RECT  5.865 0.185 5.955 0.435 ;
        RECT  5.865 0.745 5.955 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.185800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.465 0.765 ;
        RECT  2.405 0.495 3.395 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.655 -0.115 7.700 0.115 ;
        RECT  7.570 -0.115 7.655 0.430 ;
        RECT  7.280 -0.115 7.570 0.115 ;
        RECT  7.190 -0.115 7.280 0.285 ;
        RECT  6.890 -0.115 7.190 0.115 ;
        RECT  6.805 -0.115 6.890 0.285 ;
        RECT  6.520 -0.115 6.805 0.115 ;
        RECT  6.430 -0.115 6.520 0.285 ;
        RECT  6.135 -0.115 6.430 0.115 ;
        RECT  6.050 -0.115 6.135 0.285 ;
        RECT  5.750 -0.115 6.050 0.115 ;
        RECT  5.680 -0.115 5.750 0.440 ;
        RECT  5.370 -0.115 5.680 0.115 ;
        RECT  5.250 -0.115 5.370 0.145 ;
        RECT  5.000 -0.115 5.250 0.115 ;
        RECT  4.870 -0.115 5.000 0.145 ;
        RECT  4.610 -0.115 4.870 0.115 ;
        RECT  4.490 -0.115 4.610 0.145 ;
        RECT  3.040 -0.115 4.490 0.115 ;
        RECT  2.900 -0.115 3.040 0.145 ;
        RECT  2.635 -0.115 2.900 0.115 ;
        RECT  2.520 -0.115 2.635 0.145 ;
        RECT  2.265 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.265 0.145 ;
        RECT  1.860 -0.115 2.140 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.260 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.665 1.145 7.700 1.375 ;
        RECT  7.570 0.720 7.665 1.375 ;
        RECT  7.285 1.145 7.570 1.375 ;
        RECT  7.190 0.965 7.285 1.375 ;
        RECT  6.900 1.145 7.190 1.375 ;
        RECT  6.805 0.965 6.900 1.375 ;
        RECT  6.525 1.145 6.805 1.375 ;
        RECT  6.430 0.965 6.525 1.375 ;
        RECT  6.135 1.145 6.430 1.375 ;
        RECT  6.050 0.965 6.135 1.375 ;
        RECT  5.770 1.145 6.050 1.375 ;
        RECT  5.650 1.005 5.770 1.375 ;
        RECT  5.350 1.145 5.650 1.375 ;
        RECT  5.275 0.990 5.350 1.375 ;
        RECT  4.970 1.145 5.275 1.375 ;
        RECT  4.895 0.990 4.970 1.375 ;
        RECT  4.590 1.145 4.895 1.375 ;
        RECT  4.470 1.130 4.590 1.375 ;
        RECT  4.215 1.145 4.470 1.375 ;
        RECT  4.085 1.130 4.215 1.375 ;
        RECT  3.830 1.145 4.085 1.375 ;
        RECT  3.710 1.130 3.830 1.375 ;
        RECT  1.885 1.145 3.710 1.375 ;
        RECT  1.815 0.745 1.885 1.375 ;
        RECT  1.540 1.145 1.815 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.375 0.185 7.465 0.435 ;
        RECT  7.380 0.745 7.465 1.045 ;
        RECT  7.100 0.745 7.380 0.815 ;
        RECT  7.085 0.355 7.375 0.435 ;
        RECT  7.000 0.745 7.100 1.045 ;
        RECT  7.000 0.185 7.085 0.435 ;
        RECT  6.825 0.355 7.000 0.435 ;
        RECT  6.825 0.745 7.000 0.815 ;
        RECT  6.315 0.355 6.475 0.435 ;
        RECT  6.315 0.745 6.475 0.815 ;
        RECT  6.240 0.185 6.315 0.435 ;
        RECT  6.245 0.745 6.315 1.045 ;
        RECT  5.955 0.745 6.245 0.815 ;
        RECT  5.955 0.355 6.240 0.435 ;
        RECT  5.865 0.185 5.955 0.435 ;
        RECT  5.865 0.745 5.955 1.045 ;
        RECT  5.785 0.540 6.285 0.620 ;
        RECT  5.715 0.540 5.785 0.920 ;
        RECT  2.295 0.850 5.715 0.920 ;
        RECT  5.540 0.355 5.610 0.780 ;
        RECT  5.535 0.355 5.540 0.445 ;
        RECT  4.820 0.710 5.540 0.780 ;
        RECT  5.465 0.195 5.535 0.445 ;
        RECT  5.350 0.520 5.460 0.640 ;
        RECT  5.280 0.215 5.350 0.640 ;
        RECT  1.330 0.215 5.280 0.285 ;
        RECT  2.295 0.355 5.180 0.425 ;
        RECT  4.750 0.545 4.820 0.780 ;
        RECT  2.330 0.990 4.805 1.060 ;
        RECT  3.690 0.545 4.750 0.620 ;
        RECT  2.205 0.355 2.295 0.920 ;
        RECT  2.005 0.385 2.075 1.035 ;
        RECT  1.965 0.385 2.005 0.640 ;
        RECT  1.730 0.520 1.965 0.640 ;
        RECT  1.660 0.875 1.725 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.195 0.800 0.800 ;
        RECT  0.620 0.195 0.730 0.265 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD10BWP40

MACRO CKLHQD12BWP40
    CLASS CORE ;
    FOREIGN CKLHQD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.752000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.790 0.185 7.885 0.435 ;
        RECT  7.795 0.745 7.885 1.045 ;
        RECT  7.505 0.745 7.795 0.835 ;
        RECT  7.505 0.355 7.790 0.435 ;
        RECT  7.415 0.185 7.505 0.435 ;
        RECT  7.420 0.745 7.505 1.045 ;
        RECT  7.140 0.745 7.420 0.815 ;
        RECT  7.125 0.355 7.415 0.435 ;
        RECT  7.040 0.745 7.140 1.045 ;
        RECT  7.040 0.185 7.125 0.435 ;
        RECT  7.035 0.355 7.040 0.435 ;
        RECT  7.035 0.745 7.040 0.815 ;
        RECT  6.735 0.355 7.035 0.815 ;
        RECT  6.685 0.185 6.735 1.045 ;
        RECT  6.655 0.185 6.685 0.435 ;
        RECT  6.660 0.745 6.685 1.045 ;
        RECT  6.355 0.745 6.660 0.815 ;
        RECT  6.355 0.355 6.655 0.435 ;
        RECT  6.280 0.185 6.355 0.435 ;
        RECT  6.285 0.745 6.355 1.045 ;
        RECT  5.995 0.745 6.285 0.815 ;
        RECT  5.995 0.355 6.280 0.435 ;
        RECT  5.905 0.185 5.995 0.435 ;
        RECT  5.905 0.745 5.995 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.181000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.465 0.765 ;
        RECT  2.405 0.495 3.395 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.075 -0.115 8.120 0.115 ;
        RECT  7.990 -0.115 8.075 0.430 ;
        RECT  7.690 -0.115 7.990 0.115 ;
        RECT  7.615 -0.115 7.690 0.285 ;
        RECT  7.320 -0.115 7.615 0.115 ;
        RECT  7.230 -0.115 7.320 0.285 ;
        RECT  6.930 -0.115 7.230 0.115 ;
        RECT  6.845 -0.115 6.930 0.285 ;
        RECT  6.560 -0.115 6.845 0.115 ;
        RECT  6.470 -0.115 6.560 0.285 ;
        RECT  6.175 -0.115 6.470 0.115 ;
        RECT  6.090 -0.115 6.175 0.285 ;
        RECT  5.750 -0.115 6.090 0.115 ;
        RECT  5.680 -0.115 5.750 0.440 ;
        RECT  5.370 -0.115 5.680 0.115 ;
        RECT  5.250 -0.115 5.370 0.145 ;
        RECT  5.000 -0.115 5.250 0.115 ;
        RECT  4.870 -0.115 5.000 0.145 ;
        RECT  4.610 -0.115 4.870 0.115 ;
        RECT  4.490 -0.115 4.610 0.145 ;
        RECT  3.040 -0.115 4.490 0.115 ;
        RECT  2.900 -0.115 3.040 0.145 ;
        RECT  2.635 -0.115 2.900 0.115 ;
        RECT  2.520 -0.115 2.635 0.145 ;
        RECT  2.265 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.265 0.145 ;
        RECT  1.860 -0.115 2.140 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.260 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.085 1.145 8.120 1.375 ;
        RECT  7.990 0.720 8.085 1.375 ;
        RECT  7.705 1.145 7.990 1.375 ;
        RECT  7.615 0.965 7.705 1.375 ;
        RECT  7.325 1.145 7.615 1.375 ;
        RECT  7.230 0.965 7.325 1.375 ;
        RECT  6.940 1.145 7.230 1.375 ;
        RECT  6.845 0.965 6.940 1.375 ;
        RECT  6.565 1.145 6.845 1.375 ;
        RECT  6.470 0.965 6.565 1.375 ;
        RECT  6.175 1.145 6.470 1.375 ;
        RECT  6.090 0.965 6.175 1.375 ;
        RECT  5.770 1.145 6.090 1.375 ;
        RECT  5.650 1.005 5.770 1.375 ;
        RECT  5.350 1.145 5.650 1.375 ;
        RECT  5.275 0.990 5.350 1.375 ;
        RECT  4.970 1.145 5.275 1.375 ;
        RECT  4.895 0.990 4.970 1.375 ;
        RECT  4.590 1.145 4.895 1.375 ;
        RECT  4.470 1.130 4.590 1.375 ;
        RECT  4.215 1.145 4.470 1.375 ;
        RECT  4.085 1.130 4.215 1.375 ;
        RECT  3.830 1.145 4.085 1.375 ;
        RECT  3.710 1.130 3.830 1.375 ;
        RECT  1.885 1.145 3.710 1.375 ;
        RECT  1.815 0.745 1.885 1.375 ;
        RECT  1.540 1.145 1.815 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.790 0.185 7.885 0.435 ;
        RECT  7.795 0.745 7.885 1.045 ;
        RECT  7.505 0.745 7.795 0.835 ;
        RECT  7.505 0.355 7.790 0.435 ;
        RECT  7.415 0.185 7.505 0.435 ;
        RECT  7.420 0.745 7.505 1.045 ;
        RECT  7.140 0.745 7.420 0.815 ;
        RECT  7.125 0.355 7.415 0.435 ;
        RECT  7.105 0.745 7.140 1.045 ;
        RECT  7.105 0.185 7.125 0.435 ;
        RECT  6.355 0.355 6.615 0.435 ;
        RECT  6.355 0.745 6.615 0.815 ;
        RECT  6.280 0.185 6.355 0.435 ;
        RECT  6.285 0.745 6.355 1.045 ;
        RECT  5.995 0.745 6.285 0.815 ;
        RECT  5.995 0.355 6.280 0.435 ;
        RECT  5.905 0.185 5.995 0.435 ;
        RECT  5.905 0.745 5.995 1.045 ;
        RECT  5.810 0.525 6.520 0.635 ;
        RECT  5.715 0.525 5.810 0.920 ;
        RECT  2.295 0.850 5.715 0.920 ;
        RECT  5.540 0.355 5.610 0.780 ;
        RECT  5.535 0.355 5.540 0.445 ;
        RECT  4.820 0.710 5.540 0.780 ;
        RECT  5.465 0.195 5.535 0.445 ;
        RECT  5.350 0.520 5.460 0.640 ;
        RECT  5.280 0.215 5.350 0.640 ;
        RECT  1.330 0.215 5.280 0.285 ;
        RECT  2.295 0.355 5.180 0.425 ;
        RECT  4.750 0.545 4.820 0.780 ;
        RECT  2.330 0.990 4.805 1.060 ;
        RECT  3.730 0.545 4.750 0.620 ;
        RECT  2.205 0.355 2.295 0.920 ;
        RECT  2.005 0.385 2.075 1.035 ;
        RECT  1.965 0.385 2.005 0.640 ;
        RECT  1.730 0.520 1.965 0.640 ;
        RECT  1.660 0.875 1.725 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.195 0.800 0.800 ;
        RECT  0.620 0.195 0.730 0.265 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD12BWP40

MACRO CKLHQD14BWP40
    CLASS CORE ;
    FOREIGN CKLHQD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.872000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.920 0.745 9.010 1.045 ;
        RECT  8.915 0.185 8.995 0.435 ;
        RECT  8.625 0.745 8.920 0.835 ;
        RECT  8.625 0.355 8.915 0.435 ;
        RECT  8.530 0.185 8.625 0.435 ;
        RECT  8.535 0.745 8.625 1.045 ;
        RECT  8.245 0.745 8.535 0.835 ;
        RECT  8.245 0.355 8.530 0.435 ;
        RECT  8.155 0.185 8.245 0.435 ;
        RECT  8.160 0.745 8.245 1.045 ;
        RECT  8.015 0.745 8.160 0.815 ;
        RECT  8.015 0.355 8.155 0.435 ;
        RECT  7.880 0.355 8.015 0.815 ;
        RECT  7.865 0.355 7.880 1.045 ;
        RECT  7.780 0.185 7.865 1.045 ;
        RECT  7.665 0.355 7.780 0.815 ;
        RECT  7.475 0.355 7.665 0.435 ;
        RECT  7.475 0.745 7.665 0.815 ;
        RECT  7.395 0.185 7.475 0.435 ;
        RECT  7.400 0.745 7.475 1.045 ;
        RECT  7.095 0.745 7.400 0.815 ;
        RECT  7.095 0.355 7.395 0.435 ;
        RECT  7.020 0.185 7.095 0.435 ;
        RECT  7.025 0.745 7.095 1.045 ;
        RECT  6.700 0.745 7.025 0.815 ;
        RECT  6.700 0.355 7.020 0.435 ;
        RECT  6.610 0.185 6.700 0.435 ;
        RECT  6.610 0.745 6.700 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.205800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.495 3.745 0.765 ;
        RECT  2.405 0.495 3.675 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.185 -0.115 9.240 0.115 ;
        RECT  9.110 -0.115 9.185 0.430 ;
        RECT  8.815 -0.115 9.110 0.115 ;
        RECT  8.715 -0.115 8.815 0.285 ;
        RECT  8.430 -0.115 8.715 0.115 ;
        RECT  8.355 -0.115 8.430 0.285 ;
        RECT  8.060 -0.115 8.355 0.115 ;
        RECT  7.970 -0.115 8.060 0.285 ;
        RECT  7.670 -0.115 7.970 0.115 ;
        RECT  7.585 -0.115 7.670 0.285 ;
        RECT  7.300 -0.115 7.585 0.115 ;
        RECT  7.210 -0.115 7.300 0.285 ;
        RECT  6.880 -0.115 7.210 0.115 ;
        RECT  6.795 -0.115 6.880 0.285 ;
        RECT  6.455 -0.115 6.795 0.115 ;
        RECT  6.385 -0.115 6.455 0.440 ;
        RECT  6.075 -0.115 6.385 0.115 ;
        RECT  5.915 -0.115 6.075 0.145 ;
        RECT  5.680 -0.115 5.915 0.115 ;
        RECT  5.555 -0.115 5.680 0.145 ;
        RECT  5.300 -0.115 5.555 0.115 ;
        RECT  5.175 -0.115 5.300 0.145 ;
        RECT  4.915 -0.115 5.175 0.115 ;
        RECT  4.795 -0.115 4.915 0.145 ;
        RECT  3.020 -0.115 4.795 0.115 ;
        RECT  2.900 -0.115 3.020 0.145 ;
        RECT  2.660 -0.115 2.900 0.115 ;
        RECT  2.520 -0.115 2.660 0.145 ;
        RECT  2.280 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.280 0.145 ;
        RECT  1.860 -0.115 2.140 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.185 1.145 9.240 1.375 ;
        RECT  9.105 0.720 9.185 1.375 ;
        RECT  8.810 1.145 9.105 1.375 ;
        RECT  8.725 0.965 8.810 1.375 ;
        RECT  8.445 1.145 8.725 1.375 ;
        RECT  8.355 0.965 8.445 1.375 ;
        RECT  8.065 1.145 8.355 1.375 ;
        RECT  7.970 0.965 8.065 1.375 ;
        RECT  7.680 1.145 7.970 1.375 ;
        RECT  7.585 0.965 7.680 1.375 ;
        RECT  7.305 1.145 7.585 1.375 ;
        RECT  7.210 0.965 7.305 1.375 ;
        RECT  6.880 1.145 7.210 1.375 ;
        RECT  6.795 0.965 6.880 1.375 ;
        RECT  6.460 1.145 6.795 1.375 ;
        RECT  6.370 1.005 6.460 1.375 ;
        RECT  6.040 1.145 6.370 1.375 ;
        RECT  5.955 0.990 6.040 1.375 ;
        RECT  5.655 1.145 5.955 1.375 ;
        RECT  5.580 0.990 5.655 1.375 ;
        RECT  5.285 1.145 5.580 1.375 ;
        RECT  5.120 1.130 5.285 1.375 ;
        RECT  4.880 1.145 5.120 1.375 ;
        RECT  4.740 1.130 4.880 1.375 ;
        RECT  4.475 1.145 4.740 1.375 ;
        RECT  4.355 1.130 4.475 1.375 ;
        RECT  4.095 1.145 4.355 1.375 ;
        RECT  3.975 1.130 4.095 1.375 ;
        RECT  1.935 1.145 3.975 1.375 ;
        RECT  1.865 0.745 1.935 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.920 0.745 9.010 1.045 ;
        RECT  8.915 0.185 8.995 0.435 ;
        RECT  8.625 0.745 8.920 0.835 ;
        RECT  8.625 0.355 8.915 0.435 ;
        RECT  8.530 0.185 8.625 0.435 ;
        RECT  8.535 0.745 8.625 1.045 ;
        RECT  8.245 0.745 8.535 0.835 ;
        RECT  8.245 0.355 8.530 0.435 ;
        RECT  8.155 0.185 8.245 0.435 ;
        RECT  8.160 0.745 8.245 1.045 ;
        RECT  8.085 0.745 8.160 0.815 ;
        RECT  8.085 0.355 8.155 0.435 ;
        RECT  7.475 0.355 7.595 0.435 ;
        RECT  7.475 0.745 7.595 0.815 ;
        RECT  7.395 0.185 7.475 0.435 ;
        RECT  7.400 0.745 7.475 1.045 ;
        RECT  7.095 0.745 7.400 0.815 ;
        RECT  7.095 0.355 7.395 0.435 ;
        RECT  7.020 0.185 7.095 0.435 ;
        RECT  7.025 0.745 7.095 1.045 ;
        RECT  6.700 0.745 7.025 0.815 ;
        RECT  6.700 0.355 7.020 0.435 ;
        RECT  6.610 0.185 6.700 0.435 ;
        RECT  6.610 0.745 6.700 1.045 ;
        RECT  6.490 0.525 7.535 0.635 ;
        RECT  6.420 0.525 6.490 0.920 ;
        RECT  2.335 0.850 6.420 0.920 ;
        RECT  6.225 0.355 6.295 0.780 ;
        RECT  6.220 0.355 6.225 0.445 ;
        RECT  5.430 0.710 6.225 0.780 ;
        RECT  6.150 0.195 6.220 0.445 ;
        RECT  6.035 0.520 6.145 0.640 ;
        RECT  5.965 0.215 6.035 0.640 ;
        RECT  1.330 0.215 5.965 0.285 ;
        RECT  2.335 0.355 5.865 0.425 ;
        RECT  2.415 0.990 5.490 1.060 ;
        RECT  5.360 0.545 5.430 0.780 ;
        RECT  4.155 0.545 5.360 0.615 ;
        RECT  2.245 0.355 2.335 0.920 ;
        RECT  2.055 0.375 2.125 1.035 ;
        RECT  1.960 0.375 2.055 0.445 ;
        RECT  1.730 0.520 2.055 0.640 ;
        RECT  1.660 0.880 1.740 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.810 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.730 0.185 0.810 0.800 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD14BWP40

MACRO CKLHQD16BWP40
    CLASS CORE ;
    FOREIGN CKLHQD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.000000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.040 0.185 10.125 0.435 ;
        RECT  10.045 0.745 10.125 1.045 ;
        RECT  9.750 0.745 10.045 0.835 ;
        RECT  9.735 0.355 10.040 0.435 ;
        RECT  9.660 0.745 9.750 1.045 ;
        RECT  9.655 0.185 9.735 0.435 ;
        RECT  9.365 0.745 9.660 0.835 ;
        RECT  9.365 0.355 9.655 0.435 ;
        RECT  9.270 0.185 9.365 0.435 ;
        RECT  9.275 0.745 9.365 1.045 ;
        RECT  8.985 0.745 9.275 0.835 ;
        RECT  8.985 0.355 9.270 0.435 ;
        RECT  8.895 0.185 8.985 0.435 ;
        RECT  8.900 0.745 8.985 1.045 ;
        RECT  8.855 0.745 8.900 0.815 ;
        RECT  8.855 0.355 8.895 0.435 ;
        RECT  8.620 0.355 8.855 0.815 ;
        RECT  8.605 0.355 8.620 1.045 ;
        RECT  8.520 0.185 8.605 1.045 ;
        RECT  8.505 0.355 8.520 0.815 ;
        RECT  8.215 0.355 8.505 0.435 ;
        RECT  8.215 0.745 8.505 0.815 ;
        RECT  8.135 0.185 8.215 0.435 ;
        RECT  8.140 0.745 8.215 1.045 ;
        RECT  7.835 0.745 8.140 0.815 ;
        RECT  7.835 0.355 8.135 0.435 ;
        RECT  7.760 0.185 7.835 0.435 ;
        RECT  7.765 0.745 7.835 1.045 ;
        RECT  7.425 0.745 7.765 0.815 ;
        RECT  7.425 0.355 7.760 0.435 ;
        RECT  7.335 0.185 7.425 0.435 ;
        RECT  7.335 0.745 7.425 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.249400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.495 4.165 0.765 ;
        RECT  2.500 0.495 4.095 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.305 -0.115 10.360 0.115 ;
        RECT  10.230 -0.115 10.305 0.420 ;
        RECT  9.940 -0.115 10.230 0.115 ;
        RECT  9.850 -0.115 9.940 0.285 ;
        RECT  9.555 -0.115 9.850 0.115 ;
        RECT  9.455 -0.115 9.555 0.285 ;
        RECT  9.170 -0.115 9.455 0.115 ;
        RECT  9.095 -0.115 9.170 0.285 ;
        RECT  8.800 -0.115 9.095 0.115 ;
        RECT  8.710 -0.115 8.800 0.285 ;
        RECT  8.410 -0.115 8.710 0.115 ;
        RECT  8.325 -0.115 8.410 0.285 ;
        RECT  8.040 -0.115 8.325 0.115 ;
        RECT  7.950 -0.115 8.040 0.285 ;
        RECT  7.625 -0.115 7.950 0.115 ;
        RECT  7.540 -0.115 7.625 0.285 ;
        RECT  7.200 -0.115 7.540 0.115 ;
        RECT  7.130 -0.115 7.200 0.440 ;
        RECT  6.800 -0.115 7.130 0.115 ;
        RECT  6.660 -0.115 6.800 0.145 ;
        RECT  6.430 -0.115 6.660 0.115 ;
        RECT  6.300 -0.115 6.430 0.145 ;
        RECT  6.050 -0.115 6.300 0.115 ;
        RECT  5.920 -0.115 6.050 0.145 ;
        RECT  5.670 -0.115 5.920 0.115 ;
        RECT  5.545 -0.115 5.670 0.145 ;
        RECT  3.460 -0.115 5.545 0.115 ;
        RECT  3.320 -0.115 3.460 0.145 ;
        RECT  3.080 -0.115 3.320 0.115 ;
        RECT  2.960 -0.115 3.080 0.145 ;
        RECT  2.720 -0.115 2.960 0.115 ;
        RECT  2.580 -0.115 2.720 0.145 ;
        RECT  2.310 -0.115 2.580 0.115 ;
        RECT  2.170 -0.115 2.310 0.145 ;
        RECT  1.860 -0.115 2.170 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.305 1.145 10.360 1.375 ;
        RECT  10.225 0.720 10.305 1.375 ;
        RECT  9.935 1.145 10.225 1.375 ;
        RECT  9.850 0.965 9.935 1.375 ;
        RECT  9.550 1.145 9.850 1.375 ;
        RECT  9.465 0.965 9.550 1.375 ;
        RECT  9.185 1.145 9.465 1.375 ;
        RECT  9.095 0.965 9.185 1.375 ;
        RECT  8.805 1.145 9.095 1.375 ;
        RECT  8.710 0.965 8.805 1.375 ;
        RECT  8.420 1.145 8.710 1.375 ;
        RECT  8.325 0.965 8.420 1.375 ;
        RECT  8.045 1.145 8.325 1.375 ;
        RECT  7.950 0.965 8.045 1.375 ;
        RECT  7.625 1.145 7.950 1.375 ;
        RECT  7.540 0.965 7.625 1.375 ;
        RECT  7.205 1.145 7.540 1.375 ;
        RECT  7.115 1.005 7.205 1.375 ;
        RECT  6.775 1.145 7.115 1.375 ;
        RECT  6.700 0.990 6.775 1.375 ;
        RECT  6.400 1.145 6.700 1.375 ;
        RECT  6.325 0.990 6.400 1.375 ;
        RECT  6.030 1.145 6.325 1.375 ;
        RECT  5.885 1.130 6.030 1.375 ;
        RECT  5.645 1.145 5.885 1.375 ;
        RECT  5.485 1.130 5.645 1.375 ;
        RECT  5.240 1.145 5.485 1.375 ;
        RECT  5.070 1.130 5.240 1.375 ;
        RECT  4.845 1.145 5.070 1.375 ;
        RECT  4.720 1.130 4.845 1.375 ;
        RECT  4.460 1.145 4.720 1.375 ;
        RECT  4.340 1.130 4.460 1.375 ;
        RECT  1.935 1.145 4.340 1.375 ;
        RECT  1.865 0.740 1.935 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.040 0.185 10.125 0.435 ;
        RECT  10.045 0.745 10.125 1.045 ;
        RECT  9.750 0.745 10.045 0.835 ;
        RECT  9.735 0.355 10.040 0.435 ;
        RECT  9.660 0.745 9.750 1.045 ;
        RECT  9.655 0.185 9.735 0.435 ;
        RECT  9.365 0.745 9.660 0.835 ;
        RECT  9.365 0.355 9.655 0.435 ;
        RECT  9.270 0.185 9.365 0.435 ;
        RECT  9.275 0.745 9.365 1.045 ;
        RECT  8.985 0.745 9.275 0.835 ;
        RECT  8.985 0.355 9.270 0.435 ;
        RECT  8.925 0.185 8.985 0.435 ;
        RECT  8.925 0.745 8.985 1.045 ;
        RECT  8.215 0.355 8.435 0.435 ;
        RECT  8.215 0.745 8.435 0.815 ;
        RECT  8.135 0.185 8.215 0.435 ;
        RECT  8.140 0.745 8.215 1.045 ;
        RECT  7.835 0.745 8.140 0.815 ;
        RECT  7.835 0.355 8.135 0.435 ;
        RECT  7.760 0.185 7.835 0.435 ;
        RECT  7.765 0.745 7.835 1.045 ;
        RECT  7.425 0.745 7.765 0.815 ;
        RECT  7.425 0.355 7.760 0.435 ;
        RECT  7.335 0.185 7.425 0.435 ;
        RECT  7.335 0.745 7.425 1.045 ;
        RECT  7.235 0.545 8.310 0.615 ;
        RECT  7.165 0.545 7.235 0.920 ;
        RECT  2.335 0.850 7.165 0.920 ;
        RECT  6.970 0.355 7.040 0.780 ;
        RECT  6.965 0.355 6.970 0.445 ;
        RECT  6.000 0.710 6.970 0.780 ;
        RECT  6.895 0.195 6.965 0.445 ;
        RECT  6.780 0.520 6.890 0.640 ;
        RECT  6.710 0.215 6.780 0.640 ;
        RECT  1.330 0.215 6.710 0.285 ;
        RECT  2.335 0.355 6.610 0.425 ;
        RECT  2.400 0.990 6.235 1.060 ;
        RECT  5.930 0.545 6.000 0.780 ;
        RECT  4.475 0.545 5.930 0.615 ;
        RECT  2.245 0.355 2.335 0.920 ;
        RECT  2.055 0.375 2.125 1.035 ;
        RECT  1.960 0.375 2.055 0.445 ;
        RECT  1.730 0.520 2.055 0.640 ;
        RECT  1.660 0.880 1.740 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.810 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.730 0.185 0.810 0.800 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD16BWP40

MACRO CKLHQD18BWP40
    CLASS CORE ;
    FOREIGN CKLHQD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.096000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.600 0.185 10.685 0.435 ;
        RECT  10.600 0.745 10.685 1.045 ;
        RECT  10.305 0.355 10.600 0.435 ;
        RECT  10.305 0.745 10.600 0.835 ;
        RECT  10.220 0.185 10.305 0.435 ;
        RECT  10.225 0.745 10.305 1.045 ;
        RECT  9.930 0.745 10.225 0.835 ;
        RECT  9.915 0.355 10.220 0.435 ;
        RECT  9.840 0.745 9.930 1.045 ;
        RECT  9.835 0.185 9.915 0.435 ;
        RECT  9.545 0.745 9.840 0.835 ;
        RECT  9.545 0.355 9.835 0.435 ;
        RECT  9.450 0.185 9.545 0.435 ;
        RECT  9.455 0.745 9.545 1.045 ;
        RECT  9.165 0.745 9.455 0.835 ;
        RECT  9.165 0.355 9.450 0.435 ;
        RECT  9.135 0.185 9.165 0.435 ;
        RECT  9.135 0.745 9.165 1.045 ;
        RECT  9.080 0.185 9.135 1.045 ;
        RECT  9.075 0.185 9.080 0.815 ;
        RECT  8.855 0.355 9.075 0.815 ;
        RECT  8.785 0.355 8.855 0.435 ;
        RECT  8.800 0.745 8.855 0.815 ;
        RECT  8.700 0.745 8.800 1.045 ;
        RECT  8.700 0.185 8.785 0.435 ;
        RECT  8.395 0.355 8.700 0.435 ;
        RECT  8.395 0.745 8.700 0.815 ;
        RECT  8.315 0.185 8.395 0.435 ;
        RECT  8.320 0.745 8.395 1.045 ;
        RECT  8.015 0.745 8.320 0.815 ;
        RECT  8.015 0.355 8.315 0.435 ;
        RECT  7.940 0.185 8.015 0.435 ;
        RECT  7.920 0.745 8.015 1.045 ;
        RECT  7.625 0.355 7.940 0.435 ;
        RECT  7.625 0.745 7.920 0.815 ;
        RECT  7.535 0.185 7.625 0.435 ;
        RECT  7.535 0.745 7.625 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.273800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.305 0.765 ;
        RECT  2.500 0.495 4.235 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.865 -0.115 10.920 0.115 ;
        RECT  10.790 -0.115 10.865 0.420 ;
        RECT  10.500 -0.115 10.790 0.115 ;
        RECT  10.410 -0.115 10.500 0.285 ;
        RECT  10.120 -0.115 10.410 0.115 ;
        RECT  10.030 -0.115 10.120 0.285 ;
        RECT  9.735 -0.115 10.030 0.115 ;
        RECT  9.635 -0.115 9.735 0.285 ;
        RECT  9.350 -0.115 9.635 0.115 ;
        RECT  9.275 -0.115 9.350 0.285 ;
        RECT  8.980 -0.115 9.275 0.115 ;
        RECT  8.890 -0.115 8.980 0.285 ;
        RECT  8.590 -0.115 8.890 0.115 ;
        RECT  8.505 -0.115 8.590 0.285 ;
        RECT  8.220 -0.115 8.505 0.115 ;
        RECT  8.130 -0.115 8.220 0.285 ;
        RECT  7.805 -0.115 8.130 0.115 ;
        RECT  7.720 -0.115 7.805 0.285 ;
        RECT  7.400 -0.115 7.720 0.115 ;
        RECT  7.330 -0.115 7.400 0.440 ;
        RECT  7.000 -0.115 7.330 0.115 ;
        RECT  6.860 -0.115 7.000 0.145 ;
        RECT  6.630 -0.115 6.860 0.115 ;
        RECT  6.500 -0.115 6.630 0.145 ;
        RECT  6.250 -0.115 6.500 0.115 ;
        RECT  6.120 -0.115 6.250 0.145 ;
        RECT  5.870 -0.115 6.120 0.115 ;
        RECT  5.745 -0.115 5.870 0.145 ;
        RECT  3.460 -0.115 5.745 0.115 ;
        RECT  3.320 -0.115 3.460 0.145 ;
        RECT  3.080 -0.115 3.320 0.115 ;
        RECT  2.960 -0.115 3.080 0.145 ;
        RECT  2.720 -0.115 2.960 0.115 ;
        RECT  2.580 -0.115 2.720 0.145 ;
        RECT  2.310 -0.115 2.580 0.115 ;
        RECT  2.170 -0.115 2.310 0.145 ;
        RECT  1.860 -0.115 2.170 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.865 1.145 10.920 1.375 ;
        RECT  10.775 0.720 10.865 1.375 ;
        RECT  10.485 1.145 10.775 1.375 ;
        RECT  10.410 0.965 10.485 1.375 ;
        RECT  10.115 1.145 10.410 1.375 ;
        RECT  10.030 0.965 10.115 1.375 ;
        RECT  9.730 1.145 10.030 1.375 ;
        RECT  9.645 0.965 9.730 1.375 ;
        RECT  9.365 1.145 9.645 1.375 ;
        RECT  9.275 0.965 9.365 1.375 ;
        RECT  8.985 1.145 9.275 1.375 ;
        RECT  8.890 0.965 8.985 1.375 ;
        RECT  8.600 1.145 8.890 1.375 ;
        RECT  8.505 0.965 8.600 1.375 ;
        RECT  8.225 1.145 8.505 1.375 ;
        RECT  8.130 0.965 8.225 1.375 ;
        RECT  7.820 1.145 8.130 1.375 ;
        RECT  7.720 0.965 7.820 1.375 ;
        RECT  7.405 1.145 7.720 1.375 ;
        RECT  7.315 1.005 7.405 1.375 ;
        RECT  6.975 1.145 7.315 1.375 ;
        RECT  6.900 0.990 6.975 1.375 ;
        RECT  6.600 1.145 6.900 1.375 ;
        RECT  6.525 0.990 6.600 1.375 ;
        RECT  6.230 1.145 6.525 1.375 ;
        RECT  6.085 1.130 6.230 1.375 ;
        RECT  5.845 1.145 6.085 1.375 ;
        RECT  5.685 1.130 5.845 1.375 ;
        RECT  5.440 1.145 5.685 1.375 ;
        RECT  5.270 1.130 5.440 1.375 ;
        RECT  5.045 1.145 5.270 1.375 ;
        RECT  4.920 1.130 5.045 1.375 ;
        RECT  4.660 1.145 4.920 1.375 ;
        RECT  4.535 1.130 4.660 1.375 ;
        RECT  1.935 1.145 4.535 1.375 ;
        RECT  1.865 0.740 1.935 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.600 0.185 10.685 0.435 ;
        RECT  10.600 0.745 10.685 1.045 ;
        RECT  10.305 0.355 10.600 0.435 ;
        RECT  10.305 0.745 10.600 0.835 ;
        RECT  10.220 0.185 10.305 0.435 ;
        RECT  10.225 0.745 10.305 1.045 ;
        RECT  9.930 0.745 10.225 0.835 ;
        RECT  9.915 0.355 10.220 0.435 ;
        RECT  9.840 0.745 9.930 1.045 ;
        RECT  9.835 0.185 9.915 0.435 ;
        RECT  9.545 0.745 9.840 0.835 ;
        RECT  9.545 0.355 9.835 0.435 ;
        RECT  9.450 0.185 9.545 0.435 ;
        RECT  9.455 0.745 9.545 1.045 ;
        RECT  9.205 0.745 9.455 0.835 ;
        RECT  9.205 0.355 9.450 0.435 ;
        RECT  8.700 0.185 8.785 0.435 ;
        RECT  8.700 0.745 8.785 1.045 ;
        RECT  8.395 0.355 8.700 0.435 ;
        RECT  8.395 0.745 8.700 0.815 ;
        RECT  8.315 0.185 8.395 0.435 ;
        RECT  8.320 0.745 8.395 1.045 ;
        RECT  8.015 0.745 8.320 0.815 ;
        RECT  8.015 0.355 8.315 0.435 ;
        RECT  7.940 0.185 8.015 0.435 ;
        RECT  7.920 0.745 8.015 1.045 ;
        RECT  7.625 0.355 7.940 0.435 ;
        RECT  7.625 0.745 7.920 0.815 ;
        RECT  7.535 0.185 7.625 0.435 ;
        RECT  7.535 0.745 7.625 1.045 ;
        RECT  7.435 0.525 8.565 0.635 ;
        RECT  7.365 0.525 7.435 0.920 ;
        RECT  2.335 0.850 7.365 0.920 ;
        RECT  7.170 0.355 7.240 0.780 ;
        RECT  7.165 0.355 7.170 0.445 ;
        RECT  6.200 0.710 7.170 0.780 ;
        RECT  7.095 0.195 7.165 0.445 ;
        RECT  6.980 0.520 7.090 0.640 ;
        RECT  6.910 0.215 6.980 0.640 ;
        RECT  1.330 0.215 6.910 0.285 ;
        RECT  2.335 0.355 6.810 0.425 ;
        RECT  2.400 0.990 6.435 1.060 ;
        RECT  6.130 0.545 6.200 0.780 ;
        RECT  4.485 0.545 6.130 0.615 ;
        RECT  2.245 0.355 2.335 0.920 ;
        RECT  2.055 0.375 2.125 1.035 ;
        RECT  1.960 0.375 2.055 0.445 ;
        RECT  1.730 0.520 2.055 0.640 ;
        RECT  1.660 0.880 1.740 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.810 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.730 0.185 0.810 0.800 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD18BWP40

MACRO CKLHQD1BWP40
    CLASS CORE ;
    FOREIGN CKLHQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.185 3.045 1.045 ;
        RECT  2.955 0.185 2.975 0.465 ;
        RECT  2.955 0.745 2.975 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.046400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.495 1.925 0.640 ;
        RECT  1.715 0.495 1.805 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 3.080 0.115 ;
        RECT  2.770 -0.115 2.840 0.440 ;
        RECT  2.440 -0.115 2.770 0.115 ;
        RECT  2.310 -0.115 2.440 0.125 ;
        RECT  2.090 -0.115 2.310 0.115 ;
        RECT  1.970 -0.115 2.090 0.125 ;
        RECT  1.670 -0.115 1.970 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.270 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.145 3.080 1.375 ;
        RECT  2.740 1.005 2.860 1.375 ;
        RECT  2.480 1.145 2.740 1.375 ;
        RECT  2.360 1.000 2.480 1.375 ;
        RECT  1.720 1.145 2.360 1.375 ;
        RECT  1.600 1.000 1.720 1.375 ;
        RECT  1.150 1.145 1.600 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.875 0.520 2.895 0.640 ;
        RECT  2.805 0.520 2.875 0.920 ;
        RECT  2.065 0.850 2.805 0.920 ;
        RECT  2.615 0.195 2.685 0.780 ;
        RECT  2.585 0.195 2.615 0.450 ;
        RECT  2.325 0.710 2.615 0.780 ;
        RECT  2.505 0.525 2.535 0.640 ;
        RECT  2.435 0.195 2.505 0.640 ;
        RECT  1.330 0.195 2.435 0.265 ;
        RECT  2.255 0.520 2.325 0.780 ;
        RECT  2.065 0.355 2.260 0.425 ;
        RECT  1.995 0.355 2.065 1.035 ;
        RECT  1.645 0.355 1.890 0.425 ;
        RECT  1.815 0.860 1.885 1.035 ;
        RECT  1.645 0.860 1.815 0.930 ;
        RECT  1.575 0.355 1.645 0.930 ;
        RECT  1.540 0.520 1.575 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.345 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.195 1.330 0.810 ;
        RECT  1.180 0.195 1.260 0.265 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.195 0.800 0.800 ;
        RECT  0.620 0.195 0.730 0.265 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD1BWP40

MACRO CKLHQD20BWP40
    CLASS CORE ;
    FOREIGN CKLHQD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.232000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.020 0.185 11.105 0.435 ;
        RECT  11.020 0.745 11.105 1.045 ;
        RECT  10.725 0.355 11.020 0.435 ;
        RECT  10.725 0.745 11.020 0.835 ;
        RECT  10.640 0.185 10.725 0.435 ;
        RECT  10.640 0.745 10.725 1.045 ;
        RECT  10.345 0.355 10.640 0.435 ;
        RECT  10.345 0.745 10.640 0.835 ;
        RECT  10.260 0.185 10.345 0.435 ;
        RECT  10.265 0.745 10.345 1.045 ;
        RECT  9.970 0.745 10.265 0.835 ;
        RECT  9.955 0.355 10.260 0.435 ;
        RECT  9.880 0.745 9.970 1.045 ;
        RECT  9.875 0.185 9.955 0.435 ;
        RECT  9.585 0.745 9.880 0.835 ;
        RECT  9.585 0.355 9.875 0.435 ;
        RECT  9.490 0.185 9.585 0.435 ;
        RECT  9.495 0.745 9.585 1.045 ;
        RECT  9.415 0.745 9.495 0.835 ;
        RECT  9.415 0.355 9.490 0.435 ;
        RECT  9.205 0.355 9.415 0.835 ;
        RECT  9.120 0.185 9.205 1.045 ;
        RECT  9.115 0.185 9.120 0.815 ;
        RECT  9.065 0.355 9.115 0.815 ;
        RECT  8.825 0.355 9.065 0.435 ;
        RECT  8.840 0.745 9.065 0.815 ;
        RECT  8.740 0.745 8.840 1.045 ;
        RECT  8.740 0.185 8.825 0.435 ;
        RECT  8.435 0.355 8.740 0.435 ;
        RECT  8.435 0.745 8.740 0.815 ;
        RECT  8.355 0.185 8.435 0.435 ;
        RECT  8.360 0.745 8.435 1.045 ;
        RECT  8.025 0.745 8.360 0.815 ;
        RECT  8.025 0.355 8.355 0.435 ;
        RECT  7.950 0.185 8.025 0.435 ;
        RECT  7.955 0.745 8.025 1.045 ;
        RECT  7.625 0.745 7.955 0.815 ;
        RECT  7.625 0.355 7.950 0.435 ;
        RECT  7.535 0.185 7.625 0.435 ;
        RECT  7.535 0.745 7.625 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.271400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 0.495 4.315 0.765 ;
        RECT  2.500 0.495 4.225 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.285 -0.115 11.340 0.115 ;
        RECT  11.210 -0.115 11.285 0.430 ;
        RECT  10.920 -0.115 11.210 0.115 ;
        RECT  10.830 -0.115 10.920 0.285 ;
        RECT  10.540 -0.115 10.830 0.115 ;
        RECT  10.450 -0.115 10.540 0.285 ;
        RECT  10.160 -0.115 10.450 0.115 ;
        RECT  10.070 -0.115 10.160 0.285 ;
        RECT  9.775 -0.115 10.070 0.115 ;
        RECT  9.675 -0.115 9.775 0.285 ;
        RECT  9.390 -0.115 9.675 0.115 ;
        RECT  9.315 -0.115 9.390 0.285 ;
        RECT  9.020 -0.115 9.315 0.115 ;
        RECT  8.930 -0.115 9.020 0.285 ;
        RECT  8.630 -0.115 8.930 0.115 ;
        RECT  8.545 -0.115 8.630 0.285 ;
        RECT  8.260 -0.115 8.545 0.115 ;
        RECT  8.170 -0.115 8.260 0.285 ;
        RECT  7.825 -0.115 8.170 0.115 ;
        RECT  7.740 -0.115 7.825 0.285 ;
        RECT  7.400 -0.115 7.740 0.115 ;
        RECT  7.330 -0.115 7.400 0.440 ;
        RECT  7.000 -0.115 7.330 0.115 ;
        RECT  6.860 -0.115 7.000 0.145 ;
        RECT  6.630 -0.115 6.860 0.115 ;
        RECT  6.500 -0.115 6.630 0.145 ;
        RECT  6.250 -0.115 6.500 0.115 ;
        RECT  6.120 -0.115 6.250 0.145 ;
        RECT  5.870 -0.115 6.120 0.115 ;
        RECT  5.745 -0.115 5.870 0.145 ;
        RECT  3.460 -0.115 5.745 0.115 ;
        RECT  3.320 -0.115 3.460 0.145 ;
        RECT  3.080 -0.115 3.320 0.115 ;
        RECT  2.960 -0.115 3.080 0.145 ;
        RECT  2.720 -0.115 2.960 0.115 ;
        RECT  2.580 -0.115 2.720 0.145 ;
        RECT  2.310 -0.115 2.580 0.115 ;
        RECT  2.170 -0.115 2.310 0.145 ;
        RECT  1.860 -0.115 2.170 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.285 1.145 11.340 1.375 ;
        RECT  11.195 0.720 11.285 1.375 ;
        RECT  10.905 1.145 11.195 1.375 ;
        RECT  10.830 0.965 10.905 1.375 ;
        RECT  10.525 1.145 10.830 1.375 ;
        RECT  10.450 0.965 10.525 1.375 ;
        RECT  10.155 1.145 10.450 1.375 ;
        RECT  10.070 0.965 10.155 1.375 ;
        RECT  9.770 1.145 10.070 1.375 ;
        RECT  9.685 0.965 9.770 1.375 ;
        RECT  9.405 1.145 9.685 1.375 ;
        RECT  9.315 0.965 9.405 1.375 ;
        RECT  9.025 1.145 9.315 1.375 ;
        RECT  8.930 0.965 9.025 1.375 ;
        RECT  8.640 1.145 8.930 1.375 ;
        RECT  8.545 0.965 8.640 1.375 ;
        RECT  8.265 1.145 8.545 1.375 ;
        RECT  8.170 0.965 8.265 1.375 ;
        RECT  7.825 1.145 8.170 1.375 ;
        RECT  7.740 0.965 7.825 1.375 ;
        RECT  7.405 1.145 7.740 1.375 ;
        RECT  7.315 1.005 7.405 1.375 ;
        RECT  6.975 1.145 7.315 1.375 ;
        RECT  6.900 0.990 6.975 1.375 ;
        RECT  6.600 1.145 6.900 1.375 ;
        RECT  6.525 0.990 6.600 1.375 ;
        RECT  6.230 1.145 6.525 1.375 ;
        RECT  6.085 1.130 6.230 1.375 ;
        RECT  5.845 1.145 6.085 1.375 ;
        RECT  5.685 1.130 5.845 1.375 ;
        RECT  5.440 1.145 5.685 1.375 ;
        RECT  5.270 1.130 5.440 1.375 ;
        RECT  5.045 1.145 5.270 1.375 ;
        RECT  4.920 1.130 5.045 1.375 ;
        RECT  4.660 1.145 4.920 1.375 ;
        RECT  4.535 1.130 4.660 1.375 ;
        RECT  1.935 1.145 4.535 1.375 ;
        RECT  1.865 0.745 1.935 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.020 0.185 11.105 0.435 ;
        RECT  11.020 0.745 11.105 1.045 ;
        RECT  10.725 0.355 11.020 0.435 ;
        RECT  10.725 0.745 11.020 0.835 ;
        RECT  10.640 0.185 10.725 0.435 ;
        RECT  10.640 0.745 10.725 1.045 ;
        RECT  10.345 0.355 10.640 0.435 ;
        RECT  10.345 0.745 10.640 0.835 ;
        RECT  10.260 0.185 10.345 0.435 ;
        RECT  10.265 0.745 10.345 1.045 ;
        RECT  9.970 0.745 10.265 0.835 ;
        RECT  9.955 0.355 10.260 0.435 ;
        RECT  9.880 0.745 9.970 1.045 ;
        RECT  9.875 0.185 9.955 0.435 ;
        RECT  9.585 0.745 9.880 0.835 ;
        RECT  9.585 0.355 9.875 0.435 ;
        RECT  9.490 0.185 9.585 0.435 ;
        RECT  9.495 0.745 9.585 1.045 ;
        RECT  9.485 0.745 9.495 0.835 ;
        RECT  9.485 0.355 9.490 0.435 ;
        RECT  8.825 0.355 8.995 0.435 ;
        RECT  8.840 0.745 8.995 0.815 ;
        RECT  8.740 0.745 8.840 1.045 ;
        RECT  8.740 0.185 8.825 0.435 ;
        RECT  8.435 0.355 8.740 0.435 ;
        RECT  8.435 0.745 8.740 0.815 ;
        RECT  8.355 0.185 8.435 0.435 ;
        RECT  8.360 0.745 8.435 1.045 ;
        RECT  8.025 0.745 8.360 0.815 ;
        RECT  8.025 0.355 8.355 0.435 ;
        RECT  7.950 0.185 8.025 0.435 ;
        RECT  7.955 0.745 8.025 1.045 ;
        RECT  7.625 0.745 7.955 0.815 ;
        RECT  7.625 0.355 7.950 0.435 ;
        RECT  7.535 0.185 7.625 0.435 ;
        RECT  7.535 0.745 7.625 1.045 ;
        RECT  7.435 0.525 8.840 0.635 ;
        RECT  7.365 0.525 7.435 0.920 ;
        RECT  2.335 0.850 7.365 0.920 ;
        RECT  7.170 0.355 7.240 0.780 ;
        RECT  7.165 0.355 7.170 0.445 ;
        RECT  6.200 0.710 7.170 0.780 ;
        RECT  7.090 0.195 7.165 0.445 ;
        RECT  6.980 0.520 7.090 0.640 ;
        RECT  6.910 0.215 6.980 0.640 ;
        RECT  1.330 0.215 6.910 0.285 ;
        RECT  2.335 0.355 6.810 0.425 ;
        RECT  2.400 0.990 6.435 1.060 ;
        RECT  6.130 0.545 6.200 0.780 ;
        RECT  4.445 0.545 6.130 0.615 ;
        RECT  2.245 0.355 2.335 0.920 ;
        RECT  2.055 0.375 2.125 1.035 ;
        RECT  1.960 0.375 2.055 0.445 ;
        RECT  1.730 0.520 2.055 0.640 ;
        RECT  1.660 0.880 1.740 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.810 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.730 0.185 0.810 0.800 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD20BWP40

MACRO CKLHQD24BWP40
    CLASS CORE ;
    FOREIGN CKLHQD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.440000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.840 0.185 12.925 0.435 ;
        RECT  12.835 0.745 12.925 1.045 ;
        RECT  12.540 0.355 12.840 0.435 ;
        RECT  12.545 0.745 12.835 0.835 ;
        RECT  12.460 0.745 12.545 1.045 ;
        RECT  12.460 0.185 12.540 0.435 ;
        RECT  12.185 0.355 12.460 0.435 ;
        RECT  12.185 0.745 12.460 0.835 ;
        RECT  12.080 0.185 12.185 0.435 ;
        RECT  12.080 0.745 12.185 1.045 ;
        RECT  11.785 0.355 12.080 0.435 ;
        RECT  11.785 0.745 12.080 0.835 ;
        RECT  11.695 0.185 11.785 0.435 ;
        RECT  11.695 0.745 11.785 1.045 ;
        RECT  11.405 0.355 11.695 0.435 ;
        RECT  11.405 0.745 11.695 0.835 ;
        RECT  11.320 0.185 11.405 0.435 ;
        RECT  11.325 0.745 11.405 1.045 ;
        RECT  11.030 0.745 11.325 0.835 ;
        RECT  11.015 0.355 11.320 0.435 ;
        RECT  10.940 0.745 11.030 1.045 ;
        RECT  10.935 0.185 11.015 0.435 ;
        RECT  10.815 0.745 10.940 0.835 ;
        RECT  10.815 0.355 10.935 0.435 ;
        RECT  10.645 0.355 10.815 0.835 ;
        RECT  10.550 0.185 10.645 1.045 ;
        RECT  10.535 0.355 10.550 1.045 ;
        RECT  10.465 0.355 10.535 0.835 ;
        RECT  10.265 0.355 10.465 0.435 ;
        RECT  10.265 0.745 10.465 0.835 ;
        RECT  10.175 0.185 10.265 0.435 ;
        RECT  10.155 0.745 10.265 1.045 ;
        RECT  9.885 0.355 10.175 0.435 ;
        RECT  9.875 0.745 10.155 0.815 ;
        RECT  9.800 0.185 9.885 0.435 ;
        RECT  9.800 0.745 9.875 1.045 ;
        RECT  9.495 0.355 9.800 0.435 ;
        RECT  9.525 0.745 9.800 0.815 ;
        RECT  9.420 0.745 9.525 1.045 ;
        RECT  9.415 0.185 9.495 0.435 ;
        RECT  9.115 0.745 9.420 0.815 ;
        RECT  9.115 0.355 9.415 0.435 ;
        RECT  9.040 0.185 9.115 0.435 ;
        RECT  9.035 0.745 9.115 1.045 ;
        RECT  8.755 0.355 9.040 0.435 ;
        RECT  8.755 0.745 9.035 0.815 ;
        RECT  8.665 0.185 8.755 0.435 ;
        RECT  8.665 0.745 8.755 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.322600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.495 4.725 0.765 ;
        RECT  2.500 0.495 4.655 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.105 -0.115 13.160 0.115 ;
        RECT  13.030 -0.115 13.105 0.450 ;
        RECT  12.735 -0.115 13.030 0.115 ;
        RECT  12.645 -0.115 12.735 0.285 ;
        RECT  12.355 -0.115 12.645 0.115 ;
        RECT  12.265 -0.115 12.355 0.285 ;
        RECT  11.980 -0.115 12.265 0.115 ;
        RECT  11.890 -0.115 11.980 0.285 ;
        RECT  11.600 -0.115 11.890 0.115 ;
        RECT  11.510 -0.115 11.600 0.285 ;
        RECT  11.220 -0.115 11.510 0.115 ;
        RECT  11.130 -0.115 11.220 0.285 ;
        RECT  10.835 -0.115 11.130 0.115 ;
        RECT  10.735 -0.115 10.835 0.285 ;
        RECT  10.450 -0.115 10.735 0.115 ;
        RECT  10.375 -0.115 10.450 0.285 ;
        RECT  10.080 -0.115 10.375 0.115 ;
        RECT  9.990 -0.115 10.080 0.285 ;
        RECT  9.690 -0.115 9.990 0.115 ;
        RECT  9.605 -0.115 9.690 0.285 ;
        RECT  9.320 -0.115 9.605 0.115 ;
        RECT  9.230 -0.115 9.320 0.285 ;
        RECT  8.935 -0.115 9.230 0.115 ;
        RECT  8.850 -0.115 8.935 0.285 ;
        RECT  8.550 -0.115 8.850 0.115 ;
        RECT  8.480 -0.115 8.550 0.440 ;
        RECT  8.115 -0.115 8.480 0.115 ;
        RECT  8.045 -0.115 8.115 0.270 ;
        RECT  7.760 -0.115 8.045 0.115 ;
        RECT  7.640 -0.115 7.760 0.145 ;
        RECT  7.385 -0.115 7.640 0.115 ;
        RECT  7.260 -0.115 7.385 0.145 ;
        RECT  7.010 -0.115 7.260 0.115 ;
        RECT  6.880 -0.115 7.010 0.145 ;
        RECT  6.630 -0.115 6.880 0.115 ;
        RECT  6.505 -0.115 6.630 0.145 ;
        RECT  6.240 -0.115 6.505 0.115 ;
        RECT  6.120 -0.115 6.240 0.145 ;
        RECT  5.860 -0.115 6.120 0.115 ;
        RECT  5.740 -0.115 5.860 0.145 ;
        RECT  3.460 -0.115 5.740 0.115 ;
        RECT  3.320 -0.115 3.460 0.145 ;
        RECT  3.080 -0.115 3.320 0.115 ;
        RECT  2.960 -0.115 3.080 0.145 ;
        RECT  2.720 -0.115 2.960 0.115 ;
        RECT  2.580 -0.115 2.720 0.145 ;
        RECT  2.310 -0.115 2.580 0.115 ;
        RECT  2.170 -0.115 2.310 0.145 ;
        RECT  1.860 -0.115 2.170 0.115 ;
        RECT  1.740 -0.115 1.860 0.125 ;
        RECT  1.500 -0.115 1.740 0.115 ;
        RECT  1.380 -0.115 1.500 0.145 ;
        RECT  1.095 -0.115 1.380 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.105 1.145 13.160 1.375 ;
        RECT  13.025 0.720 13.105 1.375 ;
        RECT  12.725 1.145 13.025 1.375 ;
        RECT  12.655 0.965 12.725 1.375 ;
        RECT  12.345 1.145 12.655 1.375 ;
        RECT  12.270 0.965 12.345 1.375 ;
        RECT  11.965 1.145 12.270 1.375 ;
        RECT  11.890 0.965 11.965 1.375 ;
        RECT  11.585 1.145 11.890 1.375 ;
        RECT  11.510 0.965 11.585 1.375 ;
        RECT  11.215 1.145 11.510 1.375 ;
        RECT  11.130 0.965 11.215 1.375 ;
        RECT  10.830 1.145 11.130 1.375 ;
        RECT  10.745 0.965 10.830 1.375 ;
        RECT  10.465 1.145 10.745 1.375 ;
        RECT  10.375 0.965 10.465 1.375 ;
        RECT  10.085 1.145 10.375 1.375 ;
        RECT  9.990 0.965 10.085 1.375 ;
        RECT  9.700 1.145 9.990 1.375 ;
        RECT  9.605 0.965 9.700 1.375 ;
        RECT  9.325 1.145 9.605 1.375 ;
        RECT  9.230 0.965 9.325 1.375 ;
        RECT  8.935 1.145 9.230 1.375 ;
        RECT  8.850 0.965 8.935 1.375 ;
        RECT  8.570 1.145 8.850 1.375 ;
        RECT  8.450 1.005 8.570 1.375 ;
        RECT  8.120 1.145 8.450 1.375 ;
        RECT  8.045 0.995 8.120 1.375 ;
        RECT  7.740 1.145 8.045 1.375 ;
        RECT  7.665 0.995 7.740 1.375 ;
        RECT  7.360 1.145 7.665 1.375 ;
        RECT  7.280 0.995 7.360 1.375 ;
        RECT  6.990 1.145 7.280 1.375 ;
        RECT  6.845 1.130 6.990 1.375 ;
        RECT  6.605 1.145 6.845 1.375 ;
        RECT  6.445 1.130 6.605 1.375 ;
        RECT  6.200 1.145 6.445 1.375 ;
        RECT  6.030 1.130 6.200 1.375 ;
        RECT  5.805 1.145 6.030 1.375 ;
        RECT  5.680 1.130 5.805 1.375 ;
        RECT  5.420 1.145 5.680 1.375 ;
        RECT  5.295 1.130 5.420 1.375 ;
        RECT  5.040 1.145 5.295 1.375 ;
        RECT  4.920 1.130 5.040 1.375 ;
        RECT  1.935 1.145 4.920 1.375 ;
        RECT  1.865 0.745 1.935 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.420 1.020 1.540 1.375 ;
        RECT  1.150 1.145 1.420 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.585 0.525 10.290 0.635 ;
        RECT  8.515 0.525 8.585 0.920 ;
        RECT  2.335 0.850 8.515 0.920 ;
        RECT  8.270 0.195 8.340 0.765 ;
        RECT  8.230 0.195 8.270 0.465 ;
        RECT  6.960 0.695 8.270 0.765 ;
        RECT  7.935 0.390 8.230 0.465 ;
        RECT  7.740 0.545 8.080 0.615 ;
        RECT  7.850 0.195 7.935 0.465 ;
        RECT  7.670 0.215 7.740 0.615 ;
        RECT  1.330 0.215 7.670 0.285 ;
        RECT  2.335 0.355 7.570 0.425 ;
        RECT  2.400 0.990 7.195 1.060 ;
        RECT  6.890 0.545 6.960 0.765 ;
        RECT  4.910 0.545 6.890 0.615 ;
        RECT  2.245 0.355 2.335 0.920 ;
        RECT  2.055 0.375 2.125 1.035 ;
        RECT  1.960 0.375 2.055 0.445 ;
        RECT  1.730 0.520 2.055 0.640 ;
        RECT  1.660 0.880 1.740 0.950 ;
        RECT  1.590 0.365 1.660 0.950 ;
        RECT  0.875 0.880 1.590 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.810 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.730 0.185 0.810 0.800 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
        RECT  11.015 0.355 11.320 0.435 ;
        RECT  10.940 0.745 11.030 1.045 ;
        RECT  10.935 0.185 11.015 0.435 ;
        RECT  10.885 0.745 10.940 0.835 ;
        RECT  10.885 0.355 10.935 0.435 ;
        RECT  10.265 0.355 10.395 0.435 ;
        RECT  10.265 0.745 10.395 0.835 ;
        RECT  10.175 0.185 10.265 0.435 ;
        RECT  10.155 0.745 10.265 1.045 ;
        RECT  9.885 0.355 10.175 0.435 ;
        RECT  9.875 0.745 10.155 0.815 ;
        RECT  9.800 0.185 9.885 0.435 ;
        RECT  9.800 0.745 9.875 1.045 ;
        RECT  9.495 0.355 9.800 0.435 ;
        RECT  9.525 0.745 9.800 0.815 ;
        RECT  9.420 0.745 9.525 1.045 ;
        RECT  9.415 0.185 9.495 0.435 ;
        RECT  9.115 0.745 9.420 0.815 ;
        RECT  9.115 0.355 9.415 0.435 ;
        RECT  9.040 0.185 9.115 0.435 ;
        RECT  9.035 0.745 9.115 1.045 ;
        RECT  8.755 0.355 9.040 0.435 ;
        RECT  8.755 0.745 9.035 0.815 ;
        RECT  8.665 0.185 8.755 0.435 ;
        RECT  8.665 0.745 8.755 1.045 ;
        RECT  12.840 0.185 12.925 0.435 ;
        RECT  12.835 0.745 12.925 1.045 ;
        RECT  12.540 0.355 12.840 0.435 ;
        RECT  12.545 0.745 12.835 0.835 ;
        RECT  12.460 0.745 12.545 1.045 ;
        RECT  12.460 0.185 12.540 0.435 ;
        RECT  12.185 0.355 12.460 0.435 ;
        RECT  12.185 0.745 12.460 0.835 ;
        RECT  12.080 0.185 12.185 0.435 ;
        RECT  12.080 0.745 12.185 1.045 ;
        RECT  11.785 0.355 12.080 0.435 ;
        RECT  11.785 0.745 12.080 0.835 ;
        RECT  11.695 0.185 11.785 0.435 ;
        RECT  11.695 0.745 11.785 1.045 ;
        RECT  11.405 0.355 11.695 0.435 ;
        RECT  11.405 0.745 11.695 0.835 ;
        RECT  11.320 0.185 11.405 0.435 ;
        RECT  11.325 0.745 11.405 1.045 ;
        RECT  11.030 0.745 11.325 0.835 ;
    END
END CKLHQD24BWP40

MACRO CKLHQD2BWP40
    CLASS CORE ;
    FOREIGN CKLHQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.555 0.355 3.605 0.815 ;
        RECT  3.535 0.185 3.555 1.045 ;
        RECT  3.465 0.185 3.535 0.435 ;
        RECT  3.465 0.745 3.535 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.069800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.495 1.925 0.640 ;
        RECT  1.715 0.495 1.805 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.735 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.735 0.285 ;
        RECT  3.350 -0.115 3.650 0.115 ;
        RECT  3.280 -0.115 3.350 0.440 ;
        RECT  2.995 -0.115 3.280 0.115 ;
        RECT  2.870 -0.115 2.995 0.145 ;
        RECT  2.080 -0.115 2.870 0.115 ;
        RECT  1.950 -0.115 2.080 0.145 ;
        RECT  1.670 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.275 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.655 0.865 3.730 1.375 ;
        RECT  3.350 1.145 3.655 1.375 ;
        RECT  3.275 1.005 3.350 1.375 ;
        RECT  2.715 1.145 3.275 1.375 ;
        RECT  2.575 1.130 2.715 1.375 ;
        RECT  1.720 1.145 2.575 1.375 ;
        RECT  1.600 1.000 1.720 1.375 ;
        RECT  1.150 1.145 1.600 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.385 0.525 3.465 0.635 ;
        RECT  3.315 0.525 3.385 0.920 ;
        RECT  2.115 0.850 3.315 0.920 ;
        RECT  3.125 0.195 3.195 0.780 ;
        RECT  3.085 0.195 3.125 0.450 ;
        RECT  2.650 0.710 3.125 0.780 ;
        RECT  3.015 0.520 3.045 0.640 ;
        RECT  2.945 0.215 3.015 0.640 ;
        RECT  1.330 0.215 2.945 0.285 ;
        RECT  2.000 0.990 2.910 1.060 ;
        RECT  2.115 0.355 2.800 0.425 ;
        RECT  2.580 0.520 2.650 0.780 ;
        RECT  2.025 0.355 2.115 0.920 ;
        RECT  1.645 0.355 1.890 0.425 ;
        RECT  1.815 0.860 1.885 1.035 ;
        RECT  1.645 0.860 1.815 0.930 ;
        RECT  1.575 0.355 1.645 0.930 ;
        RECT  1.540 0.520 1.575 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.365 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.195 0.800 0.800 ;
        RECT  0.620 0.195 0.730 0.265 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD2BWP40

MACRO CKLHQD3BWP40
    CLASS CORE ;
    FOREIGN CKLHQD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 0.435 ;
        RECT  3.815 0.745 3.885 1.045 ;
        RECT  3.795 0.185 3.815 1.045 ;
        RECT  3.790 0.185 3.795 0.815 ;
        RECT  3.605 0.365 3.790 0.815 ;
        RECT  3.505 0.365 3.605 0.435 ;
        RECT  3.505 0.745 3.605 0.815 ;
        RECT  3.395 0.185 3.505 0.435 ;
        RECT  3.415 0.745 3.505 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.069800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.495 1.925 0.640 ;
        RECT  1.715 0.495 1.805 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.685 -0.115 3.920 0.115 ;
        RECT  3.600 -0.115 3.685 0.285 ;
        RECT  3.300 -0.115 3.600 0.115 ;
        RECT  3.230 -0.115 3.300 0.440 ;
        RECT  2.945 -0.115 3.230 0.115 ;
        RECT  2.820 -0.115 2.945 0.145 ;
        RECT  2.080 -0.115 2.820 0.115 ;
        RECT  1.950 -0.115 2.080 0.145 ;
        RECT  1.670 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.275 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 1.145 3.920 1.375 ;
        RECT  3.580 0.910 3.700 1.375 ;
        RECT  3.300 1.145 3.580 1.375 ;
        RECT  3.225 1.005 3.300 1.375 ;
        RECT  2.715 1.145 3.225 1.375 ;
        RECT  2.575 1.130 2.715 1.375 ;
        RECT  1.720 1.145 2.575 1.375 ;
        RECT  1.600 1.000 1.720 1.375 ;
        RECT  1.150 1.145 1.600 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.335 0.525 3.435 0.635 ;
        RECT  3.265 0.525 3.335 0.920 ;
        RECT  2.115 0.850 3.265 0.920 ;
        RECT  3.075 0.195 3.145 0.780 ;
        RECT  3.035 0.195 3.075 0.450 ;
        RECT  2.650 0.710 3.075 0.780 ;
        RECT  2.965 0.525 2.995 0.640 ;
        RECT  2.895 0.215 2.965 0.640 ;
        RECT  2.000 0.990 2.910 1.060 ;
        RECT  1.330 0.215 2.895 0.285 ;
        RECT  2.115 0.355 2.750 0.425 ;
        RECT  2.580 0.520 2.650 0.780 ;
        RECT  2.025 0.355 2.115 0.920 ;
        RECT  1.645 0.355 1.890 0.425 ;
        RECT  1.815 0.860 1.885 1.035 ;
        RECT  1.645 0.860 1.815 0.930 ;
        RECT  1.575 0.355 1.645 0.930 ;
        RECT  1.540 0.520 1.575 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.365 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.195 0.800 0.800 ;
        RECT  0.620 0.195 0.730 0.265 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD3BWP40

MACRO CKLHQD4BWP40
    CLASS CORE ;
    FOREIGN CKLHQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.185 4.925 0.435 ;
        RECT  4.835 0.745 4.925 1.045 ;
        RECT  4.795 0.355 4.850 0.435 ;
        RECT  4.795 0.745 4.835 0.815 ;
        RECT  4.585 0.355 4.795 0.815 ;
        RECT  4.565 0.355 4.585 0.435 ;
        RECT  4.565 0.745 4.585 0.815 ;
        RECT  4.475 0.185 4.565 0.435 ;
        RECT  4.475 0.745 4.565 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.117400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 2.765 0.765 ;
        RECT  2.175 0.495 2.695 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.045 -0.115 5.125 0.475 ;
        RECT  4.745 -0.115 5.045 0.115 ;
        RECT  4.660 -0.115 4.745 0.285 ;
        RECT  4.360 -0.115 4.660 0.115 ;
        RECT  4.290 -0.115 4.360 0.440 ;
        RECT  4.020 -0.115 4.290 0.115 ;
        RECT  3.870 -0.115 4.020 0.145 ;
        RECT  3.625 -0.115 3.870 0.115 ;
        RECT  3.515 -0.115 3.625 0.145 ;
        RECT  2.470 -0.115 3.515 0.115 ;
        RECT  2.330 -0.115 2.470 0.145 ;
        RECT  2.090 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.090 0.145 ;
        RECT  1.670 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.265 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.145 1.145 5.180 1.375 ;
        RECT  5.025 0.720 5.145 1.375 ;
        RECT  4.760 1.145 5.025 1.375 ;
        RECT  4.640 0.910 4.760 1.375 ;
        RECT  4.355 1.145 4.640 1.375 ;
        RECT  4.285 1.005 4.355 1.375 ;
        RECT  4.190 1.145 4.285 1.375 ;
        RECT  4.090 0.990 4.190 1.375 ;
        RECT  3.800 1.145 4.090 1.375 ;
        RECT  3.725 1.000 3.800 1.375 ;
        RECT  3.420 1.145 3.725 1.375 ;
        RECT  3.300 1.130 3.420 1.375 ;
        RECT  3.045 1.145 3.300 1.375 ;
        RECT  2.920 1.130 3.045 1.375 ;
        RECT  1.695 1.145 2.920 1.375 ;
        RECT  1.620 0.740 1.695 1.375 ;
        RECT  1.150 1.145 1.620 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.185 4.925 0.435 ;
        RECT  4.865 0.745 4.925 1.045 ;
        RECT  4.475 0.185 4.515 0.435 ;
        RECT  4.475 0.745 4.515 1.045 ;
        RECT  4.395 0.525 4.475 0.635 ;
        RECT  4.325 0.525 4.395 0.920 ;
        RECT  2.085 0.850 4.325 0.920 ;
        RECT  4.135 0.195 4.205 0.780 ;
        RECT  4.105 0.195 4.135 0.450 ;
        RECT  3.635 0.710 4.135 0.780 ;
        RECT  4.025 0.525 4.055 0.640 ;
        RECT  3.955 0.215 4.025 0.640 ;
        RECT  1.330 0.215 3.955 0.285 ;
        RECT  2.085 0.355 3.820 0.425 ;
        RECT  3.565 0.540 3.635 0.780 ;
        RECT  2.120 0.990 3.635 1.060 ;
        RECT  3.055 0.540 3.565 0.615 ;
        RECT  1.995 0.355 2.085 0.920 ;
        RECT  1.815 0.380 1.885 1.035 ;
        RECT  1.770 0.380 1.815 0.450 ;
        RECT  1.540 0.520 1.815 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.365 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.185 0.800 0.800 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD4BWP40

MACRO CKLHQD5BWP40
    CLASS CORE ;
    FOREIGN CKLHQD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.364000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.325 0.185 5.410 0.435 ;
        RECT  5.330 0.745 5.405 1.045 ;
        RECT  5.075 0.745 5.330 0.815 ;
        RECT  5.075 0.355 5.325 0.435 ;
        RECT  5.025 0.355 5.075 0.815 ;
        RECT  4.950 0.185 5.025 1.045 ;
        RECT  4.935 0.355 4.950 1.045 ;
        RECT  4.865 0.355 4.935 0.815 ;
        RECT  4.645 0.355 4.865 0.435 ;
        RECT  4.645 0.745 4.865 0.815 ;
        RECT  4.555 0.185 4.645 0.435 ;
        RECT  4.555 0.745 4.645 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.117400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 2.765 0.765 ;
        RECT  2.175 0.495 2.695 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.230 -0.115 5.460 0.115 ;
        RECT  5.140 -0.115 5.230 0.285 ;
        RECT  4.845 -0.115 5.140 0.115 ;
        RECT  4.760 -0.115 4.845 0.285 ;
        RECT  4.360 -0.115 4.760 0.115 ;
        RECT  4.290 -0.115 4.360 0.440 ;
        RECT  4.020 -0.115 4.290 0.115 ;
        RECT  3.870 -0.115 4.020 0.145 ;
        RECT  3.625 -0.115 3.870 0.115 ;
        RECT  3.515 -0.115 3.625 0.145 ;
        RECT  2.470 -0.115 3.515 0.115 ;
        RECT  2.330 -0.115 2.470 0.145 ;
        RECT  2.090 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.090 0.145 ;
        RECT  1.670 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.280 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.240 1.145 5.460 1.375 ;
        RECT  5.120 0.910 5.240 1.375 ;
        RECT  4.860 1.145 5.120 1.375 ;
        RECT  4.740 0.910 4.860 1.375 ;
        RECT  4.355 1.145 4.740 1.375 ;
        RECT  4.285 1.005 4.355 1.375 ;
        RECT  4.190 1.145 4.285 1.375 ;
        RECT  4.090 0.990 4.190 1.375 ;
        RECT  3.800 1.145 4.090 1.375 ;
        RECT  3.725 1.000 3.800 1.375 ;
        RECT  3.420 1.145 3.725 1.375 ;
        RECT  3.300 1.130 3.420 1.375 ;
        RECT  3.045 1.145 3.300 1.375 ;
        RECT  2.920 1.130 3.045 1.375 ;
        RECT  1.695 1.145 2.920 1.375 ;
        RECT  1.625 0.735 1.695 1.375 ;
        RECT  1.150 1.145 1.625 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.325 0.185 5.410 0.435 ;
        RECT  5.330 0.745 5.405 1.045 ;
        RECT  5.145 0.745 5.330 0.815 ;
        RECT  5.145 0.355 5.325 0.435 ;
        RECT  4.645 0.355 4.795 0.435 ;
        RECT  4.645 0.745 4.795 0.815 ;
        RECT  4.555 0.185 4.645 0.435 ;
        RECT  4.555 0.745 4.645 1.045 ;
        RECT  4.395 0.525 4.590 0.635 ;
        RECT  4.325 0.525 4.395 0.920 ;
        RECT  2.085 0.850 4.325 0.920 ;
        RECT  4.135 0.195 4.205 0.780 ;
        RECT  4.105 0.195 4.135 0.450 ;
        RECT  3.660 0.710 4.135 0.780 ;
        RECT  4.025 0.525 4.055 0.640 ;
        RECT  3.955 0.215 4.025 0.640 ;
        RECT  1.330 0.215 3.955 0.285 ;
        RECT  2.085 0.355 3.820 0.425 ;
        RECT  3.590 0.545 3.660 0.780 ;
        RECT  2.120 0.990 3.635 1.060 ;
        RECT  3.060 0.545 3.590 0.615 ;
        RECT  1.995 0.355 2.085 0.920 ;
        RECT  1.815 0.380 1.885 1.035 ;
        RECT  1.770 0.380 1.815 0.450 ;
        RECT  1.540 0.520 1.815 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.365 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.185 0.800 0.800 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD5BWP40

MACRO CKLHQD6BWP40
    CLASS CORE ;
    FOREIGN CKLHQD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.235 0.185 5.335 0.465 ;
        RECT  5.240 0.745 5.335 1.045 ;
        RECT  5.075 0.745 5.240 0.815 ;
        RECT  5.075 0.355 5.235 0.465 ;
        RECT  4.935 0.355 5.075 0.815 ;
        RECT  4.865 0.185 4.935 1.045 ;
        RECT  4.860 0.185 4.865 0.455 ;
        RECT  4.845 0.745 4.865 1.045 ;
        RECT  4.575 0.355 4.860 0.455 ;
        RECT  4.575 0.745 4.845 0.815 ;
        RECT  4.485 0.185 4.575 0.455 ;
        RECT  4.485 0.745 4.575 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.115000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.485 0.765 ;
        RECT  2.175 0.495 2.415 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 -0.115 5.600 0.115 ;
        RECT  5.425 -0.115 5.515 0.435 ;
        RECT  5.140 -0.115 5.425 0.115 ;
        RECT  5.050 -0.115 5.140 0.285 ;
        RECT  4.755 -0.115 5.050 0.115 ;
        RECT  4.670 -0.115 4.755 0.285 ;
        RECT  4.360 -0.115 4.670 0.115 ;
        RECT  4.290 -0.115 4.360 0.440 ;
        RECT  4.020 -0.115 4.290 0.115 ;
        RECT  3.870 -0.115 4.020 0.145 ;
        RECT  3.625 -0.115 3.870 0.115 ;
        RECT  3.515 -0.115 3.625 0.145 ;
        RECT  2.470 -0.115 3.515 0.115 ;
        RECT  2.330 -0.115 2.470 0.145 ;
        RECT  2.090 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.090 0.145 ;
        RECT  1.670 -0.115 1.950 0.115 ;
        RECT  1.550 -0.115 1.670 0.125 ;
        RECT  1.095 -0.115 1.550 0.115 ;
        RECT  1.025 -0.115 1.095 0.265 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 1.145 5.600 1.375 ;
        RECT  5.430 0.720 5.515 1.375 ;
        RECT  5.150 1.145 5.430 1.375 ;
        RECT  5.030 0.910 5.150 1.375 ;
        RECT  4.770 1.145 5.030 1.375 ;
        RECT  4.650 0.910 4.770 1.375 ;
        RECT  4.355 1.145 4.650 1.375 ;
        RECT  4.285 1.005 4.355 1.375 ;
        RECT  4.190 1.145 4.285 1.375 ;
        RECT  4.090 0.990 4.190 1.375 ;
        RECT  3.800 1.145 4.090 1.375 ;
        RECT  3.725 1.000 3.800 1.375 ;
        RECT  3.420 1.145 3.725 1.375 ;
        RECT  3.300 1.130 3.420 1.375 ;
        RECT  3.045 1.145 3.300 1.375 ;
        RECT  2.920 1.130 3.045 1.375 ;
        RECT  1.720 1.145 2.920 1.375 ;
        RECT  1.600 1.000 1.720 1.375 ;
        RECT  1.150 1.145 1.600 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.235 0.185 5.335 0.465 ;
        RECT  5.240 0.745 5.335 1.045 ;
        RECT  5.145 0.745 5.240 0.815 ;
        RECT  5.145 0.355 5.235 0.465 ;
        RECT  4.575 0.355 4.795 0.455 ;
        RECT  4.575 0.745 4.795 0.815 ;
        RECT  4.485 0.185 4.575 0.455 ;
        RECT  4.485 0.745 4.575 1.045 ;
        RECT  4.405 0.540 4.665 0.615 ;
        RECT  4.325 0.540 4.405 0.920 ;
        RECT  2.085 0.850 4.325 0.920 ;
        RECT  4.135 0.195 4.205 0.780 ;
        RECT  4.105 0.195 4.135 0.450 ;
        RECT  3.585 0.710 4.135 0.780 ;
        RECT  4.025 0.520 4.055 0.640 ;
        RECT  3.955 0.215 4.025 0.640 ;
        RECT  1.330 0.215 3.955 0.285 ;
        RECT  2.085 0.355 3.820 0.425 ;
        RECT  2.120 0.990 3.635 1.060 ;
        RECT  3.515 0.520 3.585 0.780 ;
        RECT  1.995 0.355 2.085 0.920 ;
        RECT  1.815 0.380 1.885 1.035 ;
        RECT  1.770 0.380 1.815 0.450 ;
        RECT  1.540 0.520 1.815 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.365 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.260 0.215 1.330 0.810 ;
        RECT  1.180 0.215 1.260 0.285 ;
        RECT  0.985 0.740 1.260 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.915 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.185 0.800 0.800 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD6BWP40

MACRO CKLHQD8BWP40
    CLASS CORE ;
    FOREIGN CKLHQD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 0.745 5.940 1.045 ;
        RECT  5.840 0.185 5.925 0.435 ;
        RECT  5.535 0.355 5.840 0.435 ;
        RECT  5.535 0.745 5.840 0.815 ;
        RECT  5.455 0.185 5.535 0.435 ;
        RECT  5.460 0.745 5.535 1.045 ;
        RECT  5.355 0.745 5.460 0.815 ;
        RECT  5.355 0.355 5.455 0.435 ;
        RECT  5.155 0.355 5.355 0.815 ;
        RECT  5.080 0.185 5.155 1.045 ;
        RECT  5.075 0.355 5.080 1.045 ;
        RECT  5.005 0.355 5.075 0.815 ;
        RECT  4.795 0.355 5.005 0.435 ;
        RECT  4.795 0.745 5.005 0.815 ;
        RECT  4.705 0.185 4.795 0.435 ;
        RECT  4.705 0.745 4.795 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.405 0.905 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.137800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.625 0.765 ;
        RECT  2.195 0.495 2.555 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.115 -0.115 6.160 0.115 ;
        RECT  6.030 -0.115 6.115 0.400 ;
        RECT  5.730 -0.115 6.030 0.115 ;
        RECT  5.645 -0.115 5.730 0.285 ;
        RECT  5.360 -0.115 5.645 0.115 ;
        RECT  5.270 -0.115 5.360 0.285 ;
        RECT  4.975 -0.115 5.270 0.115 ;
        RECT  4.890 -0.115 4.975 0.285 ;
        RECT  4.590 -0.115 4.890 0.115 ;
        RECT  4.520 -0.115 4.590 0.440 ;
        RECT  4.235 -0.115 4.520 0.115 ;
        RECT  4.090 -0.115 4.235 0.145 ;
        RECT  3.975 -0.115 4.090 0.115 ;
        RECT  3.845 -0.115 3.975 0.145 ;
        RECT  3.595 -0.115 3.845 0.115 ;
        RECT  3.465 -0.115 3.595 0.145 ;
        RECT  3.200 -0.115 3.465 0.115 ;
        RECT  3.070 -0.115 3.200 0.145 ;
        RECT  2.455 -0.115 3.070 0.115 ;
        RECT  2.325 -0.115 2.455 0.145 ;
        RECT  2.075 -0.115 2.325 0.115 ;
        RECT  1.945 -0.115 2.075 0.145 ;
        RECT  1.660 -0.115 1.945 0.115 ;
        RECT  1.540 -0.115 1.660 0.125 ;
        RECT  1.095 -0.115 1.540 0.115 ;
        RECT  1.025 -0.115 1.095 0.290 ;
        RECT  0.320 -0.115 1.025 0.115 ;
        RECT  0.240 -0.115 0.320 0.265 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.110 1.145 6.160 1.375 ;
        RECT  6.035 0.720 6.110 1.375 ;
        RECT  5.750 1.145 6.035 1.375 ;
        RECT  5.630 0.910 5.750 1.375 ;
        RECT  5.370 1.145 5.630 1.375 ;
        RECT  5.250 0.910 5.370 1.375 ;
        RECT  4.990 1.145 5.250 1.375 ;
        RECT  4.870 0.910 4.990 1.375 ;
        RECT  4.590 1.145 4.870 1.375 ;
        RECT  4.515 1.005 4.590 1.375 ;
        RECT  4.420 1.145 4.515 1.375 ;
        RECT  4.320 0.990 4.420 1.375 ;
        RECT  4.010 1.145 4.320 1.375 ;
        RECT  3.935 1.005 4.010 1.375 ;
        RECT  3.650 1.145 3.935 1.375 ;
        RECT  3.530 1.130 3.650 1.375 ;
        RECT  3.275 1.145 3.530 1.375 ;
        RECT  3.150 1.130 3.275 1.375 ;
        RECT  1.750 1.145 3.150 1.375 ;
        RECT  1.630 1.000 1.750 1.375 ;
        RECT  1.150 1.145 1.630 1.375 ;
        RECT  1.030 1.020 1.150 1.375 ;
        RECT  0.130 1.145 1.030 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.840 0.745 5.940 1.045 ;
        RECT  5.840 0.185 5.925 0.435 ;
        RECT  5.535 0.355 5.840 0.435 ;
        RECT  5.535 0.745 5.840 0.815 ;
        RECT  5.455 0.185 5.535 0.435 ;
        RECT  5.460 0.745 5.535 1.045 ;
        RECT  5.425 0.745 5.460 0.815 ;
        RECT  5.425 0.355 5.455 0.435 ;
        RECT  4.795 0.355 4.935 0.435 ;
        RECT  4.795 0.745 4.935 0.815 ;
        RECT  4.705 0.185 4.795 0.435 ;
        RECT  4.705 0.745 4.795 1.045 ;
        RECT  4.625 0.525 4.705 0.635 ;
        RECT  4.555 0.525 4.625 0.920 ;
        RECT  2.125 0.850 4.555 0.920 ;
        RECT  4.375 0.195 4.445 0.780 ;
        RECT  4.335 0.195 4.375 0.450 ;
        RECT  3.755 0.710 4.375 0.780 ;
        RECT  4.255 0.520 4.295 0.640 ;
        RECT  4.160 0.215 4.255 0.640 ;
        RECT  1.320 0.215 4.160 0.285 ;
        RECT  2.195 0.990 3.840 1.060 ;
        RECT  2.125 0.355 3.780 0.425 ;
        RECT  3.685 0.520 3.755 0.780 ;
        RECT  2.035 0.355 2.125 0.920 ;
        RECT  1.845 0.355 1.915 1.035 ;
        RECT  1.770 0.355 1.845 0.640 ;
        RECT  1.540 0.520 1.770 0.640 ;
        RECT  1.470 0.885 1.505 1.025 ;
        RECT  1.400 0.355 1.470 1.025 ;
        RECT  0.875 0.880 1.400 0.950 ;
        RECT  1.250 0.215 1.320 0.810 ;
        RECT  1.180 0.215 1.250 0.285 ;
        RECT  0.985 0.740 1.250 0.810 ;
        RECT  1.110 0.370 1.180 0.640 ;
        RECT  0.800 0.370 1.110 0.440 ;
        RECT  0.905 0.520 0.985 0.810 ;
        RECT  0.805 0.880 0.875 1.065 ;
        RECT  0.545 0.995 0.805 1.065 ;
        RECT  0.730 0.185 0.800 0.800 ;
        RECT  0.620 0.185 0.730 0.255 ;
        RECT  0.715 0.730 0.730 0.800 ;
        RECT  0.645 0.730 0.715 0.905 ;
        RECT  0.550 0.345 0.630 0.640 ;
        RECT  0.545 0.570 0.550 0.640 ;
        RECT  0.475 0.570 0.545 1.065 ;
        RECT  0.470 0.195 0.530 0.265 ;
        RECT  0.400 0.195 0.470 0.415 ;
        RECT  0.125 0.345 0.400 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END CKLHQD8BWP40

MACRO CKLNQD10BWP40
    CLASS CORE ;
    FOREIGN CKLNQD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.616000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.235 0.185 5.325 0.485 ;
        RECT  5.215 0.755 5.325 1.060 ;
        RECT  4.925 0.350 5.235 0.485 ;
        RECT  4.925 0.755 5.215 0.920 ;
        RECT  4.840 0.185 4.925 0.485 ;
        RECT  4.840 0.755 4.925 1.060 ;
        RECT  4.655 0.350 4.840 0.485 ;
        RECT  4.655 0.755 4.840 0.920 ;
        RECT  4.545 0.350 4.655 0.920 ;
        RECT  4.540 0.350 4.545 1.060 ;
        RECT  4.465 0.185 4.540 1.060 ;
        RECT  4.455 0.350 4.465 1.060 ;
        RECT  4.445 0.350 4.455 0.920 ;
        RECT  4.160 0.350 4.445 0.455 ;
        RECT  4.160 0.755 4.445 0.920 ;
        RECT  4.080 0.185 4.160 0.455 ;
        RECT  4.080 0.755 4.160 1.045 ;
        RECT  3.780 0.350 4.080 0.455 ;
        RECT  3.780 0.755 4.080 0.910 ;
        RECT  3.705 0.185 3.780 0.455 ;
        RECT  3.705 0.755 3.780 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.097400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.125 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.530 -0.115 5.600 0.115 ;
        RECT  5.445 -0.115 5.530 0.460 ;
        RECT  5.125 -0.115 5.445 0.115 ;
        RECT  5.015 -0.115 5.125 0.270 ;
        RECT  4.745 -0.115 5.015 0.115 ;
        RECT  4.635 -0.115 4.745 0.270 ;
        RECT  4.365 -0.115 4.635 0.115 ;
        RECT  4.255 -0.115 4.365 0.270 ;
        RECT  3.975 -0.115 4.255 0.115 ;
        RECT  3.880 -0.115 3.975 0.245 ;
        RECT  3.590 -0.115 3.880 0.115 ;
        RECT  3.515 -0.115 3.590 0.260 ;
        RECT  3.255 -0.115 3.515 0.115 ;
        RECT  3.095 -0.115 3.255 0.140 ;
        RECT  2.000 -0.115 3.095 0.115 ;
        RECT  1.880 -0.115 2.000 0.120 ;
        RECT  1.595 -0.115 1.880 0.115 ;
        RECT  1.480 -0.115 1.595 0.145 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.540 1.145 5.600 1.375 ;
        RECT  5.455 0.720 5.540 1.375 ;
        RECT  5.115 1.145 5.455 1.375 ;
        RECT  5.030 1.005 5.115 1.375 ;
        RECT  4.745 1.145 5.030 1.375 ;
        RECT  4.645 1.005 4.745 1.375 ;
        RECT  4.350 1.145 4.645 1.375 ;
        RECT  4.275 1.005 4.350 1.375 ;
        RECT  3.975 1.145 4.275 1.375 ;
        RECT  3.885 0.985 3.975 1.375 ;
        RECT  3.600 1.145 3.885 1.375 ;
        RECT  3.500 0.850 3.600 1.375 ;
        RECT  3.205 1.145 3.500 1.375 ;
        RECT  3.130 0.850 3.205 1.375 ;
        RECT  2.825 1.145 3.130 1.375 ;
        RECT  2.750 0.865 2.825 1.375 ;
        RECT  2.435 1.145 2.750 1.375 ;
        RECT  2.355 0.865 2.435 1.375 ;
        RECT  1.960 1.145 2.355 1.375 ;
        RECT  1.840 0.985 1.960 1.375 ;
        RECT  1.580 1.145 1.840 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.235 0.185 5.325 0.485 ;
        RECT  5.215 0.755 5.325 1.060 ;
        RECT  4.925 0.350 5.235 0.485 ;
        RECT  4.925 0.755 5.215 0.920 ;
        RECT  4.840 0.185 4.925 0.485 ;
        RECT  4.840 0.755 4.925 1.060 ;
        RECT  4.725 0.350 4.840 0.485 ;
        RECT  4.725 0.755 4.840 0.920 ;
        RECT  4.160 0.350 4.375 0.455 ;
        RECT  4.160 0.755 4.375 0.920 ;
        RECT  4.080 0.185 4.160 0.455 ;
        RECT  4.080 0.755 4.160 1.045 ;
        RECT  3.780 0.350 4.080 0.455 ;
        RECT  3.780 0.755 4.080 0.910 ;
        RECT  3.705 0.185 3.780 0.455 ;
        RECT  3.705 0.755 3.780 1.040 ;
        RECT  3.625 0.545 4.210 0.615 ;
        RECT  3.555 0.350 3.625 0.765 ;
        RECT  2.445 0.350 3.555 0.420 ;
        RECT  3.400 0.695 3.555 0.765 ;
        RECT  2.540 0.210 3.430 0.280 ;
        RECT  3.315 0.695 3.400 1.075 ;
        RECT  3.025 0.695 3.315 0.765 ;
        RECT  2.305 0.545 3.305 0.615 ;
        RECT  2.940 0.695 3.025 1.075 ;
        RECT  2.650 0.695 2.940 0.765 ;
        RECT  2.540 0.695 2.650 1.075 ;
        RECT  2.375 0.300 2.445 0.420 ;
        RECT  2.235 0.215 2.305 0.615 ;
        RECT  1.390 0.215 2.235 0.285 ;
        RECT  1.895 0.355 2.155 0.425 ;
        RECT  2.065 0.845 2.135 1.050 ;
        RECT  1.895 0.845 2.065 0.915 ;
        RECT  1.825 0.355 1.895 0.915 ;
        RECT  1.800 0.520 1.825 0.655 ;
        RECT  1.730 0.355 1.755 0.465 ;
        RECT  1.660 0.355 1.730 1.040 ;
        RECT  0.895 0.880 1.660 0.950 ;
        RECT  1.320 0.215 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD10BWP40

MACRO CKLNQD12BWP40
    CLASS CORE ;
    FOREIGN CKLNQD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.395 0.755 6.495 1.060 ;
        RECT  6.395 0.185 6.480 0.455 ;
        RECT  6.110 0.350 6.395 0.455 ;
        RECT  6.125 0.755 6.395 0.915 ;
        RECT  6.010 0.755 6.125 1.060 ;
        RECT  6.020 0.185 6.110 0.455 ;
        RECT  5.725 0.350 6.020 0.455 ;
        RECT  5.725 0.755 6.010 0.920 ;
        RECT  5.640 0.185 5.725 0.455 ;
        RECT  5.635 0.755 5.725 1.060 ;
        RECT  5.495 0.350 5.640 0.455 ;
        RECT  5.495 0.755 5.635 0.920 ;
        RECT  5.345 0.350 5.495 0.920 ;
        RECT  5.340 0.350 5.345 1.060 ;
        RECT  5.265 0.185 5.340 1.060 ;
        RECT  5.255 0.350 5.265 1.060 ;
        RECT  5.145 0.350 5.255 0.920 ;
        RECT  4.960 0.350 5.145 0.455 ;
        RECT  4.960 0.755 5.145 0.920 ;
        RECT  4.880 0.185 4.960 0.455 ;
        RECT  4.880 0.755 4.960 1.045 ;
        RECT  4.580 0.350 4.880 0.455 ;
        RECT  4.580 0.755 4.880 0.910 ;
        RECT  4.505 0.185 4.580 0.455 ;
        RECT  4.505 0.755 4.580 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.121000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.670 -0.115 6.720 0.115 ;
        RECT  6.585 -0.115 6.670 0.460 ;
        RECT  6.305 -0.115 6.585 0.115 ;
        RECT  6.195 -0.115 6.305 0.270 ;
        RECT  5.925 -0.115 6.195 0.115 ;
        RECT  5.815 -0.115 5.925 0.270 ;
        RECT  5.545 -0.115 5.815 0.115 ;
        RECT  5.435 -0.115 5.545 0.270 ;
        RECT  5.165 -0.115 5.435 0.115 ;
        RECT  5.055 -0.115 5.165 0.270 ;
        RECT  4.775 -0.115 5.055 0.115 ;
        RECT  4.680 -0.115 4.775 0.245 ;
        RECT  4.390 -0.115 4.680 0.115 ;
        RECT  4.315 -0.115 4.390 0.260 ;
        RECT  4.055 -0.115 4.315 0.115 ;
        RECT  3.895 -0.115 4.055 0.140 ;
        RECT  3.650 -0.115 3.895 0.115 ;
        RECT  3.530 -0.115 3.650 0.140 ;
        RECT  2.240 -0.115 3.530 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.235 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.145 6.720 1.375 ;
        RECT  6.585 0.720 6.670 1.375 ;
        RECT  6.290 1.145 6.585 1.375 ;
        RECT  6.210 1.005 6.290 1.375 ;
        RECT  5.915 1.145 6.210 1.375 ;
        RECT  5.830 1.005 5.915 1.375 ;
        RECT  5.545 1.145 5.830 1.375 ;
        RECT  5.445 1.005 5.545 1.375 ;
        RECT  5.150 1.145 5.445 1.375 ;
        RECT  5.075 1.005 5.150 1.375 ;
        RECT  4.775 1.145 5.075 1.375 ;
        RECT  4.685 0.985 4.775 1.375 ;
        RECT  4.400 1.145 4.685 1.375 ;
        RECT  4.300 0.850 4.400 1.375 ;
        RECT  4.005 1.145 4.300 1.375 ;
        RECT  3.930 0.850 4.005 1.375 ;
        RECT  3.635 1.145 3.930 1.375 ;
        RECT  3.550 0.865 3.635 1.375 ;
        RECT  3.450 1.145 3.550 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.865 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.395 0.755 6.495 1.060 ;
        RECT  6.395 0.185 6.480 0.455 ;
        RECT  6.110 0.350 6.395 0.455 ;
        RECT  6.125 0.755 6.395 0.915 ;
        RECT  6.010 0.755 6.125 1.060 ;
        RECT  6.020 0.185 6.110 0.455 ;
        RECT  5.725 0.350 6.020 0.455 ;
        RECT  5.725 0.755 6.010 0.920 ;
        RECT  5.640 0.185 5.725 0.455 ;
        RECT  5.635 0.755 5.725 1.060 ;
        RECT  5.565 0.350 5.640 0.455 ;
        RECT  5.565 0.755 5.635 0.920 ;
        RECT  4.960 0.350 5.075 0.455 ;
        RECT  4.960 0.755 5.075 0.920 ;
        RECT  4.880 0.185 4.960 0.455 ;
        RECT  4.880 0.755 4.960 1.045 ;
        RECT  4.580 0.350 4.880 0.455 ;
        RECT  4.580 0.755 4.880 0.910 ;
        RECT  4.505 0.185 4.580 0.455 ;
        RECT  4.505 0.755 4.580 1.040 ;
        RECT  4.425 0.535 4.945 0.625 ;
        RECT  4.355 0.350 4.425 0.765 ;
        RECT  2.685 0.350 4.355 0.420 ;
        RECT  4.200 0.695 4.355 0.765 ;
        RECT  2.780 0.210 4.230 0.280 ;
        RECT  4.115 0.695 4.200 1.075 ;
        RECT  2.545 0.545 4.115 0.615 ;
        RECT  3.825 0.695 4.115 0.765 ;
        RECT  3.735 0.695 3.825 1.075 ;
        RECT  3.265 0.695 3.735 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.745 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.675 0.215 1.745 0.390 ;
        RECT  1.390 0.320 1.675 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD12BWP40

MACRO CKLNQD14BWP40
    CLASS CORE ;
    FOREIGN CKLNQD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.140 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.840000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.775 0.185 6.870 0.455 ;
        RECT  6.775 0.755 6.870 1.060 ;
        RECT  6.480 0.350 6.775 0.455 ;
        RECT  6.495 0.755 6.775 0.915 ;
        RECT  6.395 0.755 6.495 1.060 ;
        RECT  6.395 0.185 6.480 0.455 ;
        RECT  6.110 0.350 6.395 0.455 ;
        RECT  6.110 0.755 6.395 0.915 ;
        RECT  6.020 0.185 6.110 0.455 ;
        RECT  6.010 0.755 6.110 1.060 ;
        RECT  5.775 0.350 6.020 0.455 ;
        RECT  5.775 0.755 6.010 0.920 ;
        RECT  5.725 0.350 5.775 0.920 ;
        RECT  5.640 0.185 5.725 1.060 ;
        RECT  5.635 0.350 5.640 1.060 ;
        RECT  5.425 0.350 5.635 0.920 ;
        RECT  5.340 0.350 5.425 0.455 ;
        RECT  5.345 0.755 5.425 0.920 ;
        RECT  5.255 0.755 5.345 1.060 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  4.960 0.350 5.265 0.455 ;
        RECT  4.960 0.755 5.255 0.920 ;
        RECT  4.880 0.185 4.960 0.455 ;
        RECT  4.880 0.755 4.960 1.035 ;
        RECT  4.580 0.350 4.880 0.455 ;
        RECT  4.580 0.755 4.880 0.910 ;
        RECT  4.505 0.185 4.580 0.455 ;
        RECT  4.505 0.755 4.580 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.122600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.060 -0.115 7.140 0.115 ;
        RECT  6.975 -0.115 7.060 0.460 ;
        RECT  6.685 -0.115 6.975 0.115 ;
        RECT  6.575 -0.115 6.685 0.270 ;
        RECT  6.305 -0.115 6.575 0.115 ;
        RECT  6.195 -0.115 6.305 0.270 ;
        RECT  5.925 -0.115 6.195 0.115 ;
        RECT  5.815 -0.115 5.925 0.270 ;
        RECT  5.545 -0.115 5.815 0.115 ;
        RECT  5.435 -0.115 5.545 0.270 ;
        RECT  5.165 -0.115 5.435 0.115 ;
        RECT  5.055 -0.115 5.165 0.270 ;
        RECT  4.775 -0.115 5.055 0.115 ;
        RECT  4.680 -0.115 4.775 0.245 ;
        RECT  4.390 -0.115 4.680 0.115 ;
        RECT  4.315 -0.115 4.390 0.260 ;
        RECT  4.055 -0.115 4.315 0.115 ;
        RECT  3.895 -0.115 4.055 0.140 ;
        RECT  3.650 -0.115 3.895 0.115 ;
        RECT  3.530 -0.115 3.650 0.140 ;
        RECT  2.240 -0.115 3.530 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.240 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.060 1.145 7.140 1.375 ;
        RECT  6.975 0.720 7.060 1.375 ;
        RECT  6.685 1.145 6.975 1.375 ;
        RECT  6.595 1.005 6.685 1.375 ;
        RECT  6.290 1.145 6.595 1.375 ;
        RECT  6.210 1.005 6.290 1.375 ;
        RECT  5.915 1.145 6.210 1.375 ;
        RECT  5.830 1.005 5.915 1.375 ;
        RECT  5.545 1.145 5.830 1.375 ;
        RECT  5.445 1.005 5.545 1.375 ;
        RECT  5.150 1.145 5.445 1.375 ;
        RECT  5.075 1.005 5.150 1.375 ;
        RECT  4.775 1.145 5.075 1.375 ;
        RECT  4.685 0.985 4.775 1.375 ;
        RECT  4.400 1.145 4.685 1.375 ;
        RECT  4.300 0.850 4.400 1.375 ;
        RECT  4.005 1.145 4.300 1.375 ;
        RECT  3.930 0.850 4.005 1.375 ;
        RECT  3.635 1.145 3.930 1.375 ;
        RECT  3.550 0.865 3.635 1.375 ;
        RECT  3.450 1.145 3.550 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.865 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.775 0.185 6.870 0.455 ;
        RECT  6.775 0.755 6.870 1.060 ;
        RECT  6.480 0.350 6.775 0.455 ;
        RECT  6.495 0.755 6.775 0.915 ;
        RECT  6.395 0.755 6.495 1.060 ;
        RECT  6.395 0.185 6.480 0.455 ;
        RECT  6.110 0.350 6.395 0.455 ;
        RECT  6.110 0.755 6.395 0.915 ;
        RECT  6.020 0.185 6.110 0.455 ;
        RECT  6.010 0.755 6.110 1.060 ;
        RECT  5.845 0.350 6.020 0.455 ;
        RECT  5.845 0.755 6.010 0.920 ;
        RECT  5.340 0.350 5.355 0.455 ;
        RECT  5.345 0.755 5.355 0.920 ;
        RECT  5.255 0.755 5.345 1.060 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  4.960 0.350 5.265 0.455 ;
        RECT  4.960 0.755 5.255 0.920 ;
        RECT  4.880 0.185 4.960 0.455 ;
        RECT  4.880 0.755 4.960 1.035 ;
        RECT  4.580 0.350 4.880 0.455 ;
        RECT  4.580 0.755 4.880 0.910 ;
        RECT  4.505 0.185 4.580 0.455 ;
        RECT  4.505 0.755 4.580 1.040 ;
        RECT  4.425 0.535 5.265 0.625 ;
        RECT  4.355 0.350 4.425 0.765 ;
        RECT  2.685 0.350 4.355 0.420 ;
        RECT  4.200 0.695 4.355 0.765 ;
        RECT  2.780 0.210 4.230 0.280 ;
        RECT  4.115 0.695 4.200 1.075 ;
        RECT  2.545 0.545 4.115 0.615 ;
        RECT  3.825 0.695 4.115 0.765 ;
        RECT  3.735 0.695 3.825 1.075 ;
        RECT  3.265 0.695 3.735 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.745 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.675 0.215 1.745 0.390 ;
        RECT  1.390 0.320 1.675 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD14BWP40

MACRO CKLNQD16BWP40
    CLASS CORE ;
    FOREIGN CKLNQD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.920 0.185 8.015 0.455 ;
        RECT  7.915 0.755 8.010 1.060 ;
        RECT  7.630 0.350 7.920 0.455 ;
        RECT  7.630 0.755 7.915 0.915 ;
        RECT  7.535 0.185 7.630 0.455 ;
        RECT  7.535 0.755 7.630 1.060 ;
        RECT  7.240 0.350 7.535 0.455 ;
        RECT  7.255 0.755 7.535 0.915 ;
        RECT  7.155 0.755 7.255 1.060 ;
        RECT  7.155 0.185 7.240 0.455 ;
        RECT  6.895 0.350 7.155 0.455 ;
        RECT  6.895 0.755 7.155 0.915 ;
        RECT  6.870 0.350 6.895 0.915 ;
        RECT  6.780 0.185 6.870 1.060 ;
        RECT  6.755 0.350 6.780 1.060 ;
        RECT  6.545 0.350 6.755 0.920 ;
        RECT  6.485 0.350 6.545 0.455 ;
        RECT  6.485 0.755 6.545 0.920 ;
        RECT  6.400 0.185 6.485 0.455 ;
        RECT  6.400 0.755 6.485 1.060 ;
        RECT  6.100 0.350 6.400 0.455 ;
        RECT  6.105 0.755 6.400 0.920 ;
        RECT  6.015 0.755 6.105 1.060 ;
        RECT  6.025 0.185 6.100 0.455 ;
        RECT  5.720 0.350 6.025 0.455 ;
        RECT  5.720 0.755 6.015 0.920 ;
        RECT  5.640 0.185 5.720 0.455 ;
        RECT  5.640 0.755 5.720 1.035 ;
        RECT  5.340 0.350 5.640 0.455 ;
        RECT  5.340 0.755 5.640 0.910 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  5.265 0.755 5.340 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.169000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.195 -0.115 8.260 0.115 ;
        RECT  8.110 -0.115 8.195 0.460 ;
        RECT  7.825 -0.115 8.110 0.115 ;
        RECT  7.715 -0.115 7.825 0.270 ;
        RECT  7.445 -0.115 7.715 0.115 ;
        RECT  7.335 -0.115 7.445 0.270 ;
        RECT  7.065 -0.115 7.335 0.115 ;
        RECT  6.955 -0.115 7.065 0.270 ;
        RECT  6.685 -0.115 6.955 0.115 ;
        RECT  6.575 -0.115 6.685 0.270 ;
        RECT  6.305 -0.115 6.575 0.115 ;
        RECT  6.195 -0.115 6.305 0.270 ;
        RECT  5.925 -0.115 6.195 0.115 ;
        RECT  5.815 -0.115 5.925 0.270 ;
        RECT  5.535 -0.115 5.815 0.115 ;
        RECT  5.440 -0.115 5.535 0.245 ;
        RECT  5.150 -0.115 5.440 0.115 ;
        RECT  5.075 -0.115 5.150 0.260 ;
        RECT  4.815 -0.115 5.075 0.115 ;
        RECT  4.655 -0.115 4.815 0.140 ;
        RECT  4.410 -0.115 4.655 0.115 ;
        RECT  4.290 -0.115 4.410 0.140 ;
        RECT  4.030 -0.115 4.290 0.115 ;
        RECT  3.910 -0.115 4.030 0.140 ;
        RECT  2.240 -0.115 3.910 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.235 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.195 1.145 8.260 1.375 ;
        RECT  8.110 0.720 8.195 1.375 ;
        RECT  7.825 1.145 8.110 1.375 ;
        RECT  7.715 1.010 7.825 1.375 ;
        RECT  7.445 1.145 7.715 1.375 ;
        RECT  7.335 1.005 7.445 1.375 ;
        RECT  7.050 1.145 7.335 1.375 ;
        RECT  6.970 1.005 7.050 1.375 ;
        RECT  6.675 1.145 6.970 1.375 ;
        RECT  6.590 1.005 6.675 1.375 ;
        RECT  6.305 1.145 6.590 1.375 ;
        RECT  6.205 1.005 6.305 1.375 ;
        RECT  5.910 1.145 6.205 1.375 ;
        RECT  5.835 1.005 5.910 1.375 ;
        RECT  5.535 1.145 5.835 1.375 ;
        RECT  5.445 0.985 5.535 1.375 ;
        RECT  5.160 1.145 5.445 1.375 ;
        RECT  5.060 0.850 5.160 1.375 ;
        RECT  4.765 1.145 5.060 1.375 ;
        RECT  4.690 0.850 4.765 1.375 ;
        RECT  4.395 1.145 4.690 1.375 ;
        RECT  4.310 0.865 4.395 1.375 ;
        RECT  4.015 1.145 4.310 1.375 ;
        RECT  3.935 0.865 4.015 1.375 ;
        RECT  3.835 1.145 3.935 1.375 ;
        RECT  3.740 0.920 3.835 1.375 ;
        RECT  3.450 1.145 3.740 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.865 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.920 0.185 8.015 0.455 ;
        RECT  7.915 0.755 8.010 1.060 ;
        RECT  7.630 0.350 7.920 0.455 ;
        RECT  7.630 0.755 7.915 0.915 ;
        RECT  7.535 0.185 7.630 0.455 ;
        RECT  7.535 0.755 7.630 1.060 ;
        RECT  7.240 0.350 7.535 0.455 ;
        RECT  7.255 0.755 7.535 0.915 ;
        RECT  7.155 0.755 7.255 1.060 ;
        RECT  7.155 0.185 7.240 0.455 ;
        RECT  6.965 0.350 7.155 0.455 ;
        RECT  6.965 0.755 7.155 0.915 ;
        RECT  6.400 0.185 6.475 0.455 ;
        RECT  6.400 0.755 6.475 1.060 ;
        RECT  6.100 0.350 6.400 0.455 ;
        RECT  6.105 0.755 6.400 0.920 ;
        RECT  6.015 0.755 6.105 1.060 ;
        RECT  6.025 0.185 6.100 0.455 ;
        RECT  5.720 0.350 6.025 0.455 ;
        RECT  5.720 0.755 6.015 0.920 ;
        RECT  5.640 0.185 5.720 0.455 ;
        RECT  5.640 0.755 5.720 1.035 ;
        RECT  5.340 0.350 5.640 0.455 ;
        RECT  5.340 0.755 5.640 0.910 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  5.265 0.755 5.340 1.040 ;
        RECT  5.185 0.535 6.355 0.625 ;
        RECT  5.115 0.350 5.185 0.765 ;
        RECT  2.685 0.350 5.115 0.420 ;
        RECT  4.960 0.695 5.115 0.765 ;
        RECT  2.780 0.210 4.990 0.280 ;
        RECT  4.875 0.695 4.960 1.075 ;
        RECT  2.545 0.545 4.905 0.615 ;
        RECT  4.585 0.695 4.875 0.765 ;
        RECT  4.495 0.695 4.585 1.075 ;
        RECT  4.210 0.695 4.495 0.765 ;
        RECT  4.110 0.695 4.210 1.075 ;
        RECT  3.650 0.695 4.110 0.765 ;
        RECT  3.560 0.695 3.650 1.075 ;
        RECT  3.265 0.695 3.560 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.745 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.675 0.215 1.745 0.390 ;
        RECT  1.390 0.320 1.675 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD16BWP40

MACRO CKLNQD18BWP40
    CLASS CORE ;
    FOREIGN CKLNQD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.080000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.295 0.185 8.390 0.455 ;
        RECT  8.295 0.755 8.385 1.060 ;
        RECT  8.015 0.350 8.295 0.455 ;
        RECT  8.010 0.755 8.295 0.915 ;
        RECT  7.920 0.185 8.015 0.455 ;
        RECT  7.915 0.755 8.010 1.060 ;
        RECT  7.630 0.350 7.920 0.455 ;
        RECT  7.630 0.755 7.915 0.915 ;
        RECT  7.535 0.185 7.630 0.455 ;
        RECT  7.535 0.755 7.630 1.060 ;
        RECT  7.240 0.350 7.535 0.455 ;
        RECT  7.255 0.755 7.535 0.915 ;
        RECT  7.175 0.755 7.255 1.060 ;
        RECT  7.175 0.185 7.240 0.455 ;
        RECT  7.155 0.185 7.175 1.060 ;
        RECT  6.870 0.350 7.155 0.915 ;
        RECT  6.825 0.185 6.870 1.060 ;
        RECT  6.780 0.185 6.825 0.455 ;
        RECT  6.770 0.755 6.825 1.060 ;
        RECT  6.485 0.350 6.780 0.455 ;
        RECT  6.485 0.755 6.770 0.920 ;
        RECT  6.400 0.185 6.485 0.455 ;
        RECT  6.400 0.755 6.485 1.060 ;
        RECT  6.100 0.350 6.400 0.455 ;
        RECT  6.105 0.755 6.400 0.920 ;
        RECT  6.015 0.755 6.105 1.060 ;
        RECT  6.025 0.185 6.100 0.455 ;
        RECT  5.720 0.350 6.025 0.455 ;
        RECT  5.720 0.755 6.015 0.920 ;
        RECT  5.640 0.185 5.720 0.455 ;
        RECT  5.640 0.755 5.720 1.035 ;
        RECT  5.340 0.350 5.640 0.455 ;
        RECT  5.340 0.755 5.640 0.910 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  5.265 0.755 5.340 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.169000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.615 -0.115 8.680 0.115 ;
        RECT  8.530 -0.115 8.615 0.460 ;
        RECT  8.210 -0.115 8.530 0.115 ;
        RECT  8.095 -0.115 8.210 0.270 ;
        RECT  7.825 -0.115 8.095 0.115 ;
        RECT  7.715 -0.115 7.825 0.270 ;
        RECT  7.445 -0.115 7.715 0.115 ;
        RECT  7.335 -0.115 7.445 0.270 ;
        RECT  7.065 -0.115 7.335 0.115 ;
        RECT  6.955 -0.115 7.065 0.270 ;
        RECT  6.685 -0.115 6.955 0.115 ;
        RECT  6.575 -0.115 6.685 0.270 ;
        RECT  6.305 -0.115 6.575 0.115 ;
        RECT  6.195 -0.115 6.305 0.270 ;
        RECT  5.925 -0.115 6.195 0.115 ;
        RECT  5.815 -0.115 5.925 0.270 ;
        RECT  5.535 -0.115 5.815 0.115 ;
        RECT  5.440 -0.115 5.535 0.245 ;
        RECT  5.150 -0.115 5.440 0.115 ;
        RECT  5.075 -0.115 5.150 0.260 ;
        RECT  4.815 -0.115 5.075 0.115 ;
        RECT  4.655 -0.115 4.815 0.140 ;
        RECT  4.410 -0.115 4.655 0.115 ;
        RECT  4.290 -0.115 4.410 0.140 ;
        RECT  4.030 -0.115 4.290 0.115 ;
        RECT  3.910 -0.115 4.030 0.140 ;
        RECT  2.240 -0.115 3.910 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.240 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.615 1.145 8.680 1.375 ;
        RECT  8.530 0.720 8.615 1.375 ;
        RECT  8.205 1.145 8.530 1.375 ;
        RECT  8.095 1.010 8.205 1.375 ;
        RECT  7.825 1.145 8.095 1.375 ;
        RECT  7.715 1.010 7.825 1.375 ;
        RECT  7.445 1.145 7.715 1.375 ;
        RECT  7.335 1.005 7.445 1.375 ;
        RECT  7.050 1.145 7.335 1.375 ;
        RECT  6.970 1.005 7.050 1.375 ;
        RECT  6.675 1.145 6.970 1.375 ;
        RECT  6.590 1.005 6.675 1.375 ;
        RECT  6.305 1.145 6.590 1.375 ;
        RECT  6.205 1.005 6.305 1.375 ;
        RECT  5.910 1.145 6.205 1.375 ;
        RECT  5.835 1.005 5.910 1.375 ;
        RECT  5.535 1.145 5.835 1.375 ;
        RECT  5.445 0.985 5.535 1.375 ;
        RECT  5.160 1.145 5.445 1.375 ;
        RECT  5.060 0.840 5.160 1.375 ;
        RECT  4.765 1.145 5.060 1.375 ;
        RECT  4.690 0.860 4.765 1.375 ;
        RECT  4.395 1.145 4.690 1.375 ;
        RECT  4.310 0.865 4.395 1.375 ;
        RECT  4.015 1.145 4.310 1.375 ;
        RECT  3.935 0.865 4.015 1.375 ;
        RECT  3.835 1.145 3.935 1.375 ;
        RECT  3.740 1.005 3.835 1.375 ;
        RECT  3.450 1.145 3.740 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.845 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.295 0.185 8.390 0.455 ;
        RECT  8.295 0.755 8.385 1.060 ;
        RECT  8.015 0.350 8.295 0.455 ;
        RECT  8.010 0.755 8.295 0.915 ;
        RECT  7.920 0.185 8.015 0.455 ;
        RECT  7.915 0.755 8.010 1.060 ;
        RECT  7.630 0.350 7.920 0.455 ;
        RECT  7.630 0.755 7.915 0.915 ;
        RECT  7.535 0.185 7.630 0.455 ;
        RECT  7.535 0.755 7.630 1.060 ;
        RECT  7.245 0.350 7.535 0.455 ;
        RECT  7.255 0.755 7.535 0.915 ;
        RECT  7.245 0.755 7.255 1.060 ;
        RECT  6.485 0.350 6.755 0.455 ;
        RECT  6.485 0.755 6.755 0.920 ;
        RECT  6.400 0.185 6.485 0.455 ;
        RECT  6.400 0.755 6.485 1.060 ;
        RECT  6.100 0.350 6.400 0.455 ;
        RECT  6.105 0.755 6.400 0.920 ;
        RECT  6.015 0.755 6.105 1.060 ;
        RECT  6.025 0.185 6.100 0.455 ;
        RECT  5.720 0.350 6.025 0.455 ;
        RECT  5.720 0.755 6.015 0.920 ;
        RECT  5.640 0.185 5.720 0.455 ;
        RECT  5.640 0.755 5.720 1.035 ;
        RECT  5.340 0.350 5.640 0.455 ;
        RECT  5.340 0.755 5.640 0.910 ;
        RECT  5.265 0.185 5.340 0.455 ;
        RECT  5.265 0.755 5.340 1.040 ;
        RECT  5.185 0.535 6.710 0.625 ;
        RECT  5.115 0.350 5.185 0.765 ;
        RECT  2.685 0.350 5.115 0.420 ;
        RECT  4.960 0.695 5.115 0.765 ;
        RECT  2.780 0.210 4.990 0.280 ;
        RECT  4.875 0.695 4.960 1.075 ;
        RECT  2.545 0.545 4.880 0.615 ;
        RECT  4.585 0.695 4.875 0.765 ;
        RECT  4.495 0.695 4.585 1.075 ;
        RECT  4.210 0.695 4.495 0.765 ;
        RECT  4.110 0.695 4.210 1.075 ;
        RECT  3.650 0.695 4.110 0.765 ;
        RECT  3.560 0.695 3.650 1.075 ;
        RECT  3.265 0.695 3.560 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.745 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.675 0.215 1.745 0.390 ;
        RECT  1.390 0.320 1.675 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD18BWP40

MACRO CKLNQD1BWP40
    CLASS CORE ;
    FOREIGN CKLNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.116000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.215 3.185 1.045 ;
        RECT  3.095 0.215 3.115 0.385 ;
        RECT  3.095 0.760 3.115 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.069000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.520 2.465 0.645 ;
        RECT  2.370 0.520 2.445 0.790 ;
        RECT  2.095 0.720 2.370 0.790 ;
        RECT  1.995 0.495 2.095 0.790 ;
        RECT  1.785 0.495 1.995 0.650 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.950 -0.115 3.220 0.115 ;
        RECT  2.880 -0.115 2.950 0.440 ;
        RECT  2.160 -0.115 2.880 0.115 ;
        RECT  2.020 -0.115 2.160 0.135 ;
        RECT  1.810 -0.115 2.020 0.115 ;
        RECT  1.690 -0.115 1.810 0.135 ;
        RECT  1.200 -0.115 1.690 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.145 3.220 1.375 ;
        RECT  2.860 0.885 2.940 1.375 ;
        RECT  2.335 1.145 2.860 1.375 ;
        RECT  2.265 0.865 2.335 1.375 ;
        RECT  1.770 1.145 2.265 1.375 ;
        RECT  1.650 0.985 1.770 1.375 ;
        RECT  1.170 1.145 1.650 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.980 0.520 3.005 0.640 ;
        RECT  2.910 0.520 2.980 0.815 ;
        RECT  2.605 0.745 2.910 0.815 ;
        RECT  2.730 0.205 2.800 0.640 ;
        RECT  2.275 0.205 2.730 0.275 ;
        RECT  2.605 0.965 2.730 1.075 ;
        RECT  2.535 0.345 2.605 1.075 ;
        RECT  2.405 0.345 2.535 0.415 ;
        RECT  2.455 0.955 2.535 1.075 ;
        RECT  2.195 0.205 2.275 0.650 ;
        RECT  1.390 0.205 2.195 0.275 ;
        RECT  1.710 0.355 1.970 0.425 ;
        RECT  1.875 0.845 1.945 1.050 ;
        RECT  1.710 0.845 1.875 0.915 ;
        RECT  1.640 0.355 1.710 0.915 ;
        RECT  1.610 0.520 1.640 0.655 ;
        RECT  1.540 0.345 1.570 0.455 ;
        RECT  1.470 0.345 1.540 1.040 ;
        RECT  0.895 0.880 1.470 0.950 ;
        RECT  1.320 0.205 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.640 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD1BWP40

MACRO CKLNQD20BWP40
    CLASS CORE ;
    FOREIGN CKLNQD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.200000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.870 0.185 8.980 0.455 ;
        RECT  8.875 0.755 8.975 1.060 ;
        RECT  8.585 0.755 8.875 0.915 ;
        RECT  8.590 0.350 8.870 0.455 ;
        RECT  8.495 0.185 8.590 0.455 ;
        RECT  8.495 0.755 8.585 1.060 ;
        RECT  8.215 0.350 8.495 0.455 ;
        RECT  8.210 0.755 8.495 0.915 ;
        RECT  8.120 0.185 8.215 0.455 ;
        RECT  8.115 0.755 8.210 1.060 ;
        RECT  7.830 0.350 8.120 0.455 ;
        RECT  7.830 0.755 8.115 0.915 ;
        RECT  7.735 0.185 7.830 0.455 ;
        RECT  7.735 0.755 7.830 1.060 ;
        RECT  7.455 0.350 7.735 0.455 ;
        RECT  7.455 0.755 7.735 0.915 ;
        RECT  7.440 0.350 7.455 1.060 ;
        RECT  7.355 0.185 7.440 1.060 ;
        RECT  7.105 0.350 7.355 0.915 ;
        RECT  7.070 0.350 7.105 0.455 ;
        RECT  7.070 0.755 7.105 0.915 ;
        RECT  6.980 0.185 7.070 0.455 ;
        RECT  6.970 0.755 7.070 1.060 ;
        RECT  6.685 0.350 6.980 0.455 ;
        RECT  6.685 0.755 6.970 0.920 ;
        RECT  6.600 0.185 6.685 0.455 ;
        RECT  6.600 0.755 6.685 1.060 ;
        RECT  6.300 0.350 6.600 0.455 ;
        RECT  6.305 0.755 6.600 0.920 ;
        RECT  6.215 0.755 6.305 1.060 ;
        RECT  6.225 0.185 6.300 0.455 ;
        RECT  5.920 0.350 6.225 0.455 ;
        RECT  5.920 0.755 6.215 0.920 ;
        RECT  5.840 0.185 5.920 0.455 ;
        RECT  5.840 0.755 5.920 1.035 ;
        RECT  5.540 0.350 5.840 0.455 ;
        RECT  5.540 0.755 5.840 0.910 ;
        RECT  5.465 0.185 5.540 0.455 ;
        RECT  5.465 0.755 5.540 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.192200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.175 -0.115 9.240 0.115 ;
        RECT  9.090 -0.115 9.175 0.460 ;
        RECT  8.785 -0.115 9.090 0.115 ;
        RECT  8.675 -0.115 8.785 0.270 ;
        RECT  8.410 -0.115 8.675 0.115 ;
        RECT  8.295 -0.115 8.410 0.270 ;
        RECT  8.025 -0.115 8.295 0.115 ;
        RECT  7.915 -0.115 8.025 0.270 ;
        RECT  7.645 -0.115 7.915 0.115 ;
        RECT  7.535 -0.115 7.645 0.270 ;
        RECT  7.265 -0.115 7.535 0.115 ;
        RECT  7.155 -0.115 7.265 0.270 ;
        RECT  6.885 -0.115 7.155 0.115 ;
        RECT  6.775 -0.115 6.885 0.270 ;
        RECT  6.505 -0.115 6.775 0.115 ;
        RECT  6.395 -0.115 6.505 0.270 ;
        RECT  6.125 -0.115 6.395 0.115 ;
        RECT  6.015 -0.115 6.125 0.270 ;
        RECT  5.735 -0.115 6.015 0.115 ;
        RECT  5.640 -0.115 5.735 0.245 ;
        RECT  5.350 -0.115 5.640 0.115 ;
        RECT  5.275 -0.115 5.350 0.260 ;
        RECT  5.015 -0.115 5.275 0.115 ;
        RECT  4.855 -0.115 5.015 0.140 ;
        RECT  4.610 -0.115 4.855 0.115 ;
        RECT  4.490 -0.115 4.610 0.140 ;
        RECT  4.230 -0.115 4.490 0.115 ;
        RECT  4.110 -0.115 4.230 0.140 ;
        RECT  2.240 -0.115 4.110 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.235 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.175 1.145 9.240 1.375 ;
        RECT  9.090 0.720 9.175 1.375 ;
        RECT  8.785 1.145 9.090 1.375 ;
        RECT  8.675 1.010 8.785 1.375 ;
        RECT  8.405 1.145 8.675 1.375 ;
        RECT  8.295 1.010 8.405 1.375 ;
        RECT  8.025 1.145 8.295 1.375 ;
        RECT  7.915 1.010 8.025 1.375 ;
        RECT  7.645 1.145 7.915 1.375 ;
        RECT  7.535 1.005 7.645 1.375 ;
        RECT  7.250 1.145 7.535 1.375 ;
        RECT  7.170 1.005 7.250 1.375 ;
        RECT  6.875 1.145 7.170 1.375 ;
        RECT  6.790 1.005 6.875 1.375 ;
        RECT  6.505 1.145 6.790 1.375 ;
        RECT  6.405 1.005 6.505 1.375 ;
        RECT  6.110 1.145 6.405 1.375 ;
        RECT  6.035 1.005 6.110 1.375 ;
        RECT  5.735 1.145 6.035 1.375 ;
        RECT  5.645 0.985 5.735 1.375 ;
        RECT  5.360 1.145 5.645 1.375 ;
        RECT  5.260 0.850 5.360 1.375 ;
        RECT  4.965 1.145 5.260 1.375 ;
        RECT  4.890 0.850 4.965 1.375 ;
        RECT  4.595 1.145 4.890 1.375 ;
        RECT  4.510 0.865 4.595 1.375 ;
        RECT  4.215 1.145 4.510 1.375 ;
        RECT  4.135 0.865 4.215 1.375 ;
        RECT  3.835 1.145 4.135 1.375 ;
        RECT  3.740 0.865 3.835 1.375 ;
        RECT  3.450 1.145 3.740 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.865 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.870 0.185 8.980 0.455 ;
        RECT  8.875 0.755 8.975 1.060 ;
        RECT  8.585 0.755 8.875 0.915 ;
        RECT  8.590 0.350 8.870 0.455 ;
        RECT  8.495 0.185 8.590 0.455 ;
        RECT  8.495 0.755 8.585 1.060 ;
        RECT  8.215 0.350 8.495 0.455 ;
        RECT  8.210 0.755 8.495 0.915 ;
        RECT  8.120 0.185 8.215 0.455 ;
        RECT  8.115 0.755 8.210 1.060 ;
        RECT  7.830 0.350 8.120 0.455 ;
        RECT  7.830 0.755 8.115 0.915 ;
        RECT  7.735 0.185 7.830 0.455 ;
        RECT  7.735 0.755 7.830 1.060 ;
        RECT  7.525 0.350 7.735 0.455 ;
        RECT  7.525 0.755 7.735 0.915 ;
        RECT  6.980 0.185 7.035 0.455 ;
        RECT  6.970 0.755 7.035 1.060 ;
        RECT  6.685 0.350 6.980 0.455 ;
        RECT  6.685 0.755 6.970 0.920 ;
        RECT  6.600 0.185 6.685 0.455 ;
        RECT  6.600 0.755 6.685 1.060 ;
        RECT  6.300 0.350 6.600 0.455 ;
        RECT  6.305 0.755 6.600 0.920 ;
        RECT  6.215 0.755 6.305 1.060 ;
        RECT  6.225 0.185 6.300 0.455 ;
        RECT  5.920 0.350 6.225 0.455 ;
        RECT  5.920 0.755 6.215 0.920 ;
        RECT  5.840 0.185 5.920 0.455 ;
        RECT  5.840 0.755 5.920 1.035 ;
        RECT  5.540 0.350 5.840 0.455 ;
        RECT  5.540 0.755 5.840 0.910 ;
        RECT  5.465 0.185 5.540 0.455 ;
        RECT  5.465 0.755 5.540 1.040 ;
        RECT  5.385 0.535 6.765 0.625 ;
        RECT  5.315 0.350 5.385 0.765 ;
        RECT  2.685 0.350 5.315 0.420 ;
        RECT  5.160 0.695 5.315 0.765 ;
        RECT  2.780 0.210 5.190 0.280 ;
        RECT  5.075 0.695 5.160 1.075 ;
        RECT  4.785 0.695 5.075 0.765 ;
        RECT  2.545 0.545 5.065 0.615 ;
        RECT  4.695 0.695 4.785 1.075 ;
        RECT  4.410 0.695 4.695 0.765 ;
        RECT  4.310 0.695 4.410 1.075 ;
        RECT  4.020 0.695 4.310 0.765 ;
        RECT  3.940 0.695 4.020 1.075 ;
        RECT  3.650 0.695 3.940 0.765 ;
        RECT  3.560 0.695 3.650 1.075 ;
        RECT  3.265 0.695 3.560 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.740 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.670 0.215 1.740 0.390 ;
        RECT  1.390 0.320 1.670 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD20BWP40

MACRO CKLNQD24BWP40
    CLASS CORE ;
    FOREIGN CKLNQD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.348000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.255 0.185 9.355 0.455 ;
        RECT  9.245 0.755 9.345 1.060 ;
        RECT  8.980 0.350 9.255 0.455 ;
        RECT  8.975 0.755 9.245 0.925 ;
        RECT  8.870 0.185 8.980 0.455 ;
        RECT  8.855 0.755 8.975 1.060 ;
        RECT  8.590 0.350 8.870 0.455 ;
        RECT  8.585 0.755 8.855 0.915 ;
        RECT  8.495 0.185 8.590 0.455 ;
        RECT  8.495 0.755 8.585 1.060 ;
        RECT  8.215 0.350 8.495 0.455 ;
        RECT  8.225 0.755 8.495 0.915 ;
        RECT  8.115 0.755 8.225 1.060 ;
        RECT  8.120 0.185 8.215 0.455 ;
        RECT  7.830 0.350 8.120 0.455 ;
        RECT  7.830 0.755 8.115 0.915 ;
        RECT  7.735 0.185 7.830 0.455 ;
        RECT  7.735 0.755 7.830 1.060 ;
        RECT  7.595 0.350 7.735 0.455 ;
        RECT  7.595 0.755 7.735 0.915 ;
        RECT  7.455 0.350 7.595 0.915 ;
        RECT  7.440 0.350 7.455 1.060 ;
        RECT  7.355 0.185 7.440 1.060 ;
        RECT  7.245 0.350 7.355 0.915 ;
        RECT  7.070 0.350 7.245 0.455 ;
        RECT  7.070 0.755 7.245 0.915 ;
        RECT  6.980 0.185 7.070 0.455 ;
        RECT  6.970 0.755 7.070 1.060 ;
        RECT  6.685 0.350 6.980 0.455 ;
        RECT  6.685 0.755 6.970 0.920 ;
        RECT  6.600 0.185 6.685 0.455 ;
        RECT  6.600 0.755 6.685 1.060 ;
        RECT  6.300 0.350 6.600 0.455 ;
        RECT  6.305 0.755 6.600 0.920 ;
        RECT  6.195 0.755 6.305 1.060 ;
        RECT  6.225 0.185 6.300 0.455 ;
        RECT  5.920 0.350 6.225 0.455 ;
        RECT  5.920 0.755 6.195 0.920 ;
        RECT  5.840 0.185 5.920 0.455 ;
        RECT  5.840 0.755 5.920 1.035 ;
        RECT  5.540 0.350 5.840 0.455 ;
        RECT  5.540 0.755 5.840 0.910 ;
        RECT  5.465 0.185 5.540 0.455 ;
        RECT  5.465 0.755 5.540 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.189400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 0.495 2.365 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.595 -0.115 9.660 0.115 ;
        RECT  9.505 -0.115 9.595 0.460 ;
        RECT  9.165 -0.115 9.505 0.115 ;
        RECT  9.055 -0.115 9.165 0.270 ;
        RECT  8.785 -0.115 9.055 0.115 ;
        RECT  8.675 -0.115 8.785 0.270 ;
        RECT  8.410 -0.115 8.675 0.115 ;
        RECT  8.295 -0.115 8.410 0.270 ;
        RECT  8.025 -0.115 8.295 0.115 ;
        RECT  7.915 -0.115 8.025 0.270 ;
        RECT  7.645 -0.115 7.915 0.115 ;
        RECT  7.535 -0.115 7.645 0.270 ;
        RECT  7.265 -0.115 7.535 0.115 ;
        RECT  7.155 -0.115 7.265 0.270 ;
        RECT  6.885 -0.115 7.155 0.115 ;
        RECT  6.775 -0.115 6.885 0.270 ;
        RECT  6.505 -0.115 6.775 0.115 ;
        RECT  6.395 -0.115 6.505 0.270 ;
        RECT  6.125 -0.115 6.395 0.115 ;
        RECT  6.015 -0.115 6.125 0.270 ;
        RECT  5.735 -0.115 6.015 0.115 ;
        RECT  5.640 -0.115 5.735 0.245 ;
        RECT  5.350 -0.115 5.640 0.115 ;
        RECT  5.275 -0.115 5.350 0.260 ;
        RECT  5.015 -0.115 5.275 0.115 ;
        RECT  4.855 -0.115 5.015 0.140 ;
        RECT  4.610 -0.115 4.855 0.115 ;
        RECT  4.490 -0.115 4.610 0.140 ;
        RECT  4.230 -0.115 4.490 0.115 ;
        RECT  4.110 -0.115 4.230 0.140 ;
        RECT  2.240 -0.115 4.110 0.115 ;
        RECT  2.120 -0.115 2.240 0.120 ;
        RECT  1.595 -0.115 2.120 0.115 ;
        RECT  1.480 -0.115 1.595 0.250 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.595 1.145 9.660 1.375 ;
        RECT  9.510 0.720 9.595 1.375 ;
        RECT  9.165 1.145 9.510 1.375 ;
        RECT  9.055 1.010 9.165 1.375 ;
        RECT  8.785 1.145 9.055 1.375 ;
        RECT  8.675 1.010 8.785 1.375 ;
        RECT  8.405 1.145 8.675 1.375 ;
        RECT  8.295 1.010 8.405 1.375 ;
        RECT  8.025 1.145 8.295 1.375 ;
        RECT  7.915 1.010 8.025 1.375 ;
        RECT  7.645 1.145 7.915 1.375 ;
        RECT  7.535 1.005 7.645 1.375 ;
        RECT  7.250 1.145 7.535 1.375 ;
        RECT  7.170 1.005 7.250 1.375 ;
        RECT  6.875 1.145 7.170 1.375 ;
        RECT  6.790 1.005 6.875 1.375 ;
        RECT  6.505 1.145 6.790 1.375 ;
        RECT  6.405 1.005 6.505 1.375 ;
        RECT  6.110 1.145 6.405 1.375 ;
        RECT  6.035 1.005 6.110 1.375 ;
        RECT  5.735 1.145 6.035 1.375 ;
        RECT  5.645 0.985 5.735 1.375 ;
        RECT  5.360 1.145 5.645 1.375 ;
        RECT  5.260 0.860 5.360 1.375 ;
        RECT  4.965 1.145 5.260 1.375 ;
        RECT  4.890 0.860 4.965 1.375 ;
        RECT  4.595 1.145 4.890 1.375 ;
        RECT  4.510 0.865 4.595 1.375 ;
        RECT  4.215 1.145 4.510 1.375 ;
        RECT  4.135 0.865 4.215 1.375 ;
        RECT  3.835 1.145 4.135 1.375 ;
        RECT  3.740 0.865 3.835 1.375 ;
        RECT  3.450 1.145 3.740 1.375 ;
        RECT  3.365 0.865 3.450 1.375 ;
        RECT  3.065 1.145 3.365 1.375 ;
        RECT  2.990 0.865 3.065 1.375 ;
        RECT  2.675 1.145 2.990 1.375 ;
        RECT  2.595 0.880 2.675 1.375 ;
        RECT  2.200 1.145 2.595 1.375 ;
        RECT  2.080 0.985 2.200 1.375 ;
        RECT  1.580 1.145 2.080 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.255 0.185 9.355 0.455 ;
        RECT  9.245 0.755 9.345 1.060 ;
        RECT  8.980 0.350 9.255 0.455 ;
        RECT  8.975 0.755 9.245 0.925 ;
        RECT  8.870 0.185 8.980 0.455 ;
        RECT  8.855 0.755 8.975 1.060 ;
        RECT  8.590 0.350 8.870 0.455 ;
        RECT  8.585 0.755 8.855 0.915 ;
        RECT  8.495 0.185 8.590 0.455 ;
        RECT  8.495 0.755 8.585 1.060 ;
        RECT  8.215 0.350 8.495 0.455 ;
        RECT  8.225 0.755 8.495 0.915 ;
        RECT  8.115 0.755 8.225 1.060 ;
        RECT  8.120 0.185 8.215 0.455 ;
        RECT  7.830 0.350 8.120 0.455 ;
        RECT  7.830 0.755 8.115 0.915 ;
        RECT  7.735 0.185 7.830 0.455 ;
        RECT  7.735 0.755 7.830 1.060 ;
        RECT  7.665 0.350 7.735 0.455 ;
        RECT  7.665 0.755 7.735 0.915 ;
        RECT  7.070 0.350 7.175 0.455 ;
        RECT  7.070 0.755 7.175 0.915 ;
        RECT  6.980 0.185 7.070 0.455 ;
        RECT  6.970 0.755 7.070 1.060 ;
        RECT  6.685 0.350 6.980 0.455 ;
        RECT  6.685 0.755 6.970 0.920 ;
        RECT  6.600 0.185 6.685 0.455 ;
        RECT  6.600 0.755 6.685 1.060 ;
        RECT  6.300 0.350 6.600 0.455 ;
        RECT  6.305 0.755 6.600 0.920 ;
        RECT  6.195 0.755 6.305 1.060 ;
        RECT  6.225 0.185 6.300 0.455 ;
        RECT  5.920 0.350 6.225 0.455 ;
        RECT  5.920 0.755 6.195 0.920 ;
        RECT  5.840 0.185 5.920 0.455 ;
        RECT  5.840 0.755 5.920 1.035 ;
        RECT  5.540 0.350 5.840 0.455 ;
        RECT  5.540 0.755 5.840 0.910 ;
        RECT  5.465 0.185 5.540 0.455 ;
        RECT  5.465 0.755 5.540 1.040 ;
        RECT  5.385 0.535 6.945 0.625 ;
        RECT  5.315 0.350 5.385 0.765 ;
        RECT  2.685 0.350 5.315 0.420 ;
        RECT  5.160 0.695 5.315 0.765 ;
        RECT  2.780 0.210 5.190 0.280 ;
        RECT  5.075 0.695 5.160 1.075 ;
        RECT  4.785 0.695 5.075 0.765 ;
        RECT  2.545 0.545 5.065 0.615 ;
        RECT  4.695 0.695 4.785 1.075 ;
        RECT  4.410 0.695 4.695 0.765 ;
        RECT  4.310 0.695 4.410 1.075 ;
        RECT  4.020 0.695 4.310 0.765 ;
        RECT  3.940 0.695 4.020 1.075 ;
        RECT  3.650 0.695 3.940 0.765 ;
        RECT  3.560 0.695 3.650 1.075 ;
        RECT  3.265 0.695 3.560 0.765 ;
        RECT  3.180 0.695 3.265 1.075 ;
        RECT  2.890 0.695 3.180 0.765 ;
        RECT  2.780 0.695 2.890 1.075 ;
        RECT  2.615 0.300 2.685 0.420 ;
        RECT  2.475 0.215 2.545 0.615 ;
        RECT  1.745 0.215 2.475 0.285 ;
        RECT  2.135 0.355 2.395 0.425 ;
        RECT  2.305 0.845 2.375 1.050 ;
        RECT  2.135 0.845 2.305 0.915 ;
        RECT  2.065 0.355 2.135 0.915 ;
        RECT  2.040 0.520 2.065 0.655 ;
        RECT  1.970 0.355 1.995 0.465 ;
        RECT  1.900 0.355 1.970 1.040 ;
        RECT  0.895 0.880 1.900 0.950 ;
        RECT  1.390 0.740 1.790 0.810 ;
        RECT  1.675 0.215 1.745 0.390 ;
        RECT  1.390 0.320 1.675 0.390 ;
        RECT  1.320 0.320 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD24BWP40

MACRO CKLNQD2BWP40
    CLASS CORE ;
    FOREIGN CKLNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.135 0.355 3.185 0.820 ;
        RECT  3.115 0.215 3.135 1.045 ;
        RECT  3.045 0.215 3.115 0.425 ;
        RECT  3.045 0.745 3.115 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.068600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.520 2.465 0.645 ;
        RECT  2.370 0.520 2.445 0.790 ;
        RECT  2.065 0.720 2.370 0.790 ;
        RECT  1.995 0.495 2.065 0.790 ;
        RECT  1.785 0.495 1.995 0.650 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.115 3.360 0.115 ;
        RECT  3.225 -0.115 3.305 0.285 ;
        RECT  2.930 -0.115 3.225 0.115 ;
        RECT  2.860 -0.115 2.930 0.440 ;
        RECT  2.160 -0.115 2.860 0.115 ;
        RECT  2.020 -0.115 2.160 0.135 ;
        RECT  1.810 -0.115 2.020 0.115 ;
        RECT  1.690 -0.115 1.810 0.135 ;
        RECT  1.200 -0.115 1.690 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.315 1.145 3.360 1.375 ;
        RECT  3.215 0.925 3.315 1.375 ;
        RECT  2.920 1.145 3.215 1.375 ;
        RECT  2.845 0.880 2.920 1.375 ;
        RECT  2.335 1.145 2.845 1.375 ;
        RECT  2.265 0.865 2.335 1.375 ;
        RECT  1.770 1.145 2.265 1.375 ;
        RECT  1.650 1.030 1.770 1.375 ;
        RECT  1.170 1.145 1.650 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.960 0.520 3.045 0.640 ;
        RECT  2.890 0.520 2.960 0.810 ;
        RECT  2.605 0.740 2.890 0.810 ;
        RECT  2.710 0.205 2.780 0.640 ;
        RECT  2.605 0.965 2.730 1.075 ;
        RECT  2.275 0.205 2.710 0.275 ;
        RECT  2.535 0.345 2.605 1.075 ;
        RECT  2.405 0.345 2.535 0.415 ;
        RECT  2.455 0.955 2.535 1.075 ;
        RECT  2.195 0.205 2.275 0.650 ;
        RECT  1.390 0.205 2.195 0.275 ;
        RECT  1.710 0.355 1.970 0.425 ;
        RECT  1.875 0.870 1.945 1.075 ;
        RECT  1.710 0.870 1.875 0.940 ;
        RECT  1.640 0.355 1.710 0.940 ;
        RECT  1.610 0.520 1.640 0.655 ;
        RECT  1.540 0.345 1.570 0.455 ;
        RECT  1.470 0.345 1.540 1.040 ;
        RECT  0.895 0.880 1.470 0.950 ;
        RECT  1.320 0.205 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.640 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD2BWP40

MACRO CKLNQD3BWP40
    CLASS CORE ;
    FOREIGN CKLNQD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.252000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.735 3.605 1.045 ;
        RECT  3.465 0.185 3.535 0.455 ;
        RECT  3.395 0.735 3.515 0.820 ;
        RECT  3.395 0.355 3.465 0.455 ;
        RECT  3.185 0.355 3.395 0.820 ;
        RECT  3.120 0.355 3.185 0.455 ;
        RECT  3.135 0.735 3.185 0.820 ;
        RECT  3.045 0.735 3.135 1.045 ;
        RECT  3.030 0.185 3.120 0.455 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.067000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.445 0.520 2.465 0.645 ;
        RECT  2.370 0.520 2.445 0.775 ;
        RECT  2.065 0.705 2.370 0.775 ;
        RECT  1.995 0.495 2.065 0.775 ;
        RECT  1.785 0.495 1.995 0.650 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.350 -0.115 3.640 0.115 ;
        RECT  3.255 -0.115 3.350 0.240 ;
        RECT  2.930 -0.115 3.255 0.115 ;
        RECT  2.860 -0.115 2.930 0.440 ;
        RECT  2.160 -0.115 2.860 0.115 ;
        RECT  2.020 -0.115 2.160 0.135 ;
        RECT  1.810 -0.115 2.020 0.115 ;
        RECT  1.690 -0.115 1.810 0.135 ;
        RECT  1.200 -0.115 1.690 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.340 1.145 3.640 1.375 ;
        RECT  3.220 0.910 3.340 1.375 ;
        RECT  2.940 1.145 3.220 1.375 ;
        RECT  2.820 0.910 2.940 1.375 ;
        RECT  2.340 1.145 2.820 1.375 ;
        RECT  2.265 0.845 2.340 1.375 ;
        RECT  1.770 1.145 2.265 1.375 ;
        RECT  1.650 0.985 1.770 1.375 ;
        RECT  1.170 1.145 1.650 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.960 0.535 3.070 0.640 ;
        RECT  2.890 0.535 2.960 0.820 ;
        RECT  2.605 0.750 2.890 0.820 ;
        RECT  2.710 0.205 2.780 0.640 ;
        RECT  2.605 0.965 2.730 1.075 ;
        RECT  2.275 0.205 2.710 0.275 ;
        RECT  2.535 0.345 2.605 1.075 ;
        RECT  2.405 0.345 2.535 0.415 ;
        RECT  2.455 0.955 2.535 1.075 ;
        RECT  2.195 0.205 2.275 0.635 ;
        RECT  1.390 0.205 2.195 0.275 ;
        RECT  1.710 0.355 1.970 0.425 ;
        RECT  1.875 0.845 1.945 1.050 ;
        RECT  1.710 0.845 1.875 0.915 ;
        RECT  1.640 0.355 1.710 0.915 ;
        RECT  1.610 0.520 1.640 0.655 ;
        RECT  1.540 0.345 1.570 0.455 ;
        RECT  1.470 0.345 1.540 1.040 ;
        RECT  0.895 0.880 1.470 0.950 ;
        RECT  1.320 0.205 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.640 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD3BWP40

MACRO CKLNQD4BWP40
    CLASS CORE ;
    FOREIGN CKLNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.880 0.185 3.960 0.455 ;
        RECT  3.875 0.755 3.960 1.035 ;
        RECT  3.815 0.350 3.880 0.455 ;
        RECT  3.815 0.755 3.875 0.910 ;
        RECT  3.605 0.350 3.815 0.910 ;
        RECT  3.580 0.350 3.605 0.455 ;
        RECT  3.580 0.755 3.605 0.910 ;
        RECT  3.505 0.185 3.580 0.455 ;
        RECT  3.505 0.755 3.580 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.073000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.125 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 -0.115 4.200 0.115 ;
        RECT  4.055 -0.115 4.145 0.465 ;
        RECT  3.775 -0.115 4.055 0.115 ;
        RECT  3.680 -0.115 3.775 0.245 ;
        RECT  3.390 -0.115 3.680 0.115 ;
        RECT  3.315 -0.115 3.390 0.260 ;
        RECT  3.050 -0.115 3.315 0.115 ;
        RECT  2.910 -0.115 3.050 0.140 ;
        RECT  2.000 -0.115 2.910 0.115 ;
        RECT  1.880 -0.115 2.000 0.120 ;
        RECT  1.595 -0.115 1.880 0.115 ;
        RECT  1.480 -0.115 1.595 0.145 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.155 1.145 4.200 1.375 ;
        RECT  4.065 0.715 4.155 1.375 ;
        RECT  3.775 1.145 4.065 1.375 ;
        RECT  3.685 0.985 3.775 1.375 ;
        RECT  3.385 1.145 3.685 1.375 ;
        RECT  3.315 0.845 3.385 1.375 ;
        RECT  3.005 1.145 3.315 1.375 ;
        RECT  2.930 0.865 3.005 1.375 ;
        RECT  2.825 1.145 2.930 1.375 ;
        RECT  2.750 0.925 2.825 1.375 ;
        RECT  2.425 1.145 2.750 1.375 ;
        RECT  2.345 0.875 2.425 1.375 ;
        RECT  1.960 1.145 2.345 1.375 ;
        RECT  1.840 0.985 1.960 1.375 ;
        RECT  1.580 1.145 1.840 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.185 3.960 0.455 ;
        RECT  3.885 0.755 3.960 1.035 ;
        RECT  3.505 0.185 3.535 0.455 ;
        RECT  3.505 0.755 3.535 1.040 ;
        RECT  3.425 0.545 3.535 0.635 ;
        RECT  3.355 0.350 3.425 0.765 ;
        RECT  2.535 0.350 3.355 0.420 ;
        RECT  3.215 0.695 3.355 0.765 ;
        RECT  2.450 0.210 3.230 0.280 ;
        RECT  3.105 0.695 3.215 1.075 ;
        RECT  2.305 0.545 3.205 0.615 ;
        RECT  2.655 0.695 3.105 0.765 ;
        RECT  2.545 0.695 2.655 1.075 ;
        RECT  2.375 0.210 2.450 0.345 ;
        RECT  2.235 0.215 2.305 0.615 ;
        RECT  1.390 0.215 2.235 0.285 ;
        RECT  1.895 0.355 2.155 0.425 ;
        RECT  2.065 0.845 2.135 1.050 ;
        RECT  1.895 0.845 2.065 0.915 ;
        RECT  1.825 0.355 1.895 0.915 ;
        RECT  1.800 0.520 1.825 0.655 ;
        RECT  1.730 0.355 1.755 0.465 ;
        RECT  1.660 0.355 1.730 1.040 ;
        RECT  0.895 0.880 1.660 0.950 ;
        RECT  1.320 0.215 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD4BWP40

MACRO CKLNQD5BWP40
    CLASS CORE ;
    FOREIGN CKLNQD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.384000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 0.185 4.445 0.380 ;
        RECT  4.340 0.755 4.445 1.060 ;
        RECT  3.960 0.310 4.350 0.380 ;
        RECT  3.960 0.755 4.340 0.920 ;
        RECT  3.955 0.185 3.960 0.380 ;
        RECT  3.955 0.755 3.960 1.035 ;
        RECT  3.880 0.185 3.955 1.035 ;
        RECT  3.745 0.310 3.880 0.910 ;
        RECT  3.580 0.310 3.745 0.380 ;
        RECT  3.580 0.755 3.745 0.910 ;
        RECT  3.505 0.185 3.580 0.380 ;
        RECT  3.505 0.755 3.580 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.073000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.125 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.165 -0.115 4.480 0.115 ;
        RECT  4.055 -0.115 4.165 0.240 ;
        RECT  3.775 -0.115 4.055 0.115 ;
        RECT  3.680 -0.115 3.775 0.235 ;
        RECT  3.390 -0.115 3.680 0.115 ;
        RECT  3.315 -0.115 3.390 0.260 ;
        RECT  3.050 -0.115 3.315 0.115 ;
        RECT  2.910 -0.115 3.050 0.140 ;
        RECT  2.000 -0.115 2.910 0.115 ;
        RECT  1.880 -0.115 2.000 0.120 ;
        RECT  1.595 -0.115 1.880 0.115 ;
        RECT  1.480 -0.115 1.595 0.145 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.480 1.375 ;
        RECT  4.075 1.005 4.150 1.375 ;
        RECT  3.775 1.145 4.075 1.375 ;
        RECT  3.685 0.985 3.775 1.375 ;
        RECT  3.400 1.145 3.685 1.375 ;
        RECT  3.300 0.850 3.400 1.375 ;
        RECT  3.005 1.145 3.300 1.375 ;
        RECT  2.930 0.850 3.005 1.375 ;
        RECT  2.825 1.145 2.930 1.375 ;
        RECT  2.750 0.980 2.825 1.375 ;
        RECT  2.425 1.145 2.750 1.375 ;
        RECT  2.345 0.875 2.425 1.375 ;
        RECT  1.960 1.145 2.345 1.375 ;
        RECT  1.840 0.985 1.960 1.375 ;
        RECT  1.580 1.145 1.840 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.185 4.445 0.380 ;
        RECT  4.340 0.755 4.445 1.060 ;
        RECT  4.025 0.310 4.350 0.380 ;
        RECT  4.025 0.755 4.340 0.920 ;
        RECT  3.580 0.310 3.675 0.380 ;
        RECT  3.580 0.755 3.675 0.910 ;
        RECT  3.505 0.185 3.580 0.380 ;
        RECT  3.505 0.755 3.580 1.040 ;
        RECT  3.425 0.535 3.535 0.625 ;
        RECT  3.355 0.350 3.425 0.765 ;
        RECT  2.535 0.350 3.355 0.420 ;
        RECT  3.215 0.695 3.355 0.765 ;
        RECT  2.450 0.210 3.230 0.280 ;
        RECT  3.105 0.695 3.215 1.075 ;
        RECT  2.305 0.545 3.205 0.615 ;
        RECT  2.655 0.695 3.105 0.765 ;
        RECT  2.545 0.695 2.655 1.075 ;
        RECT  2.375 0.210 2.450 0.345 ;
        RECT  2.235 0.215 2.305 0.615 ;
        RECT  1.390 0.215 2.235 0.285 ;
        RECT  1.895 0.355 2.155 0.425 ;
        RECT  2.065 0.845 2.135 1.050 ;
        RECT  1.895 0.845 2.065 0.915 ;
        RECT  1.825 0.355 1.895 0.915 ;
        RECT  1.800 0.520 1.825 0.655 ;
        RECT  1.730 0.355 1.755 0.465 ;
        RECT  1.660 0.355 1.730 1.040 ;
        RECT  0.895 0.880 1.660 0.950 ;
        RECT  1.320 0.215 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD5BWP40

MACRO CKLNQD6BWP40
    CLASS CORE ;
    FOREIGN CKLNQD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.255 0.755 4.345 1.060 ;
        RECT  4.265 0.185 4.340 0.380 ;
        RECT  4.095 0.300 4.265 0.380 ;
        RECT  4.095 0.755 4.255 0.920 ;
        RECT  3.960 0.300 4.095 0.920 ;
        RECT  3.885 0.185 3.960 1.035 ;
        RECT  3.880 0.185 3.885 0.380 ;
        RECT  3.880 0.755 3.885 1.035 ;
        RECT  3.580 0.300 3.880 0.380 ;
        RECT  3.580 0.755 3.880 0.910 ;
        RECT  3.505 0.185 3.580 0.380 ;
        RECT  3.505 0.755 3.580 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.073800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.125 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 -0.115 4.620 0.115 ;
        RECT  4.440 -0.115 4.530 0.460 ;
        RECT  4.165 -0.115 4.440 0.115 ;
        RECT  4.055 -0.115 4.165 0.220 ;
        RECT  3.780 -0.115 4.055 0.115 ;
        RECT  3.680 -0.115 3.780 0.230 ;
        RECT  3.390 -0.115 3.680 0.115 ;
        RECT  3.315 -0.115 3.390 0.260 ;
        RECT  3.050 -0.115 3.315 0.115 ;
        RECT  2.910 -0.115 3.050 0.140 ;
        RECT  2.000 -0.115 2.910 0.115 ;
        RECT  1.880 -0.115 2.000 0.120 ;
        RECT  1.595 -0.115 1.880 0.115 ;
        RECT  1.480 -0.115 1.595 0.145 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.620 1.375 ;
        RECT  4.450 0.720 4.540 1.375 ;
        RECT  4.150 1.145 4.450 1.375 ;
        RECT  4.075 1.005 4.150 1.375 ;
        RECT  3.775 1.145 4.075 1.375 ;
        RECT  3.685 0.985 3.775 1.375 ;
        RECT  3.400 1.145 3.685 1.375 ;
        RECT  3.300 0.850 3.400 1.375 ;
        RECT  3.005 1.145 3.300 1.375 ;
        RECT  2.930 0.860 3.005 1.375 ;
        RECT  2.825 1.145 2.930 1.375 ;
        RECT  2.750 0.925 2.825 1.375 ;
        RECT  2.425 1.145 2.750 1.375 ;
        RECT  2.345 0.865 2.425 1.375 ;
        RECT  1.960 1.145 2.345 1.375 ;
        RECT  1.840 0.985 1.960 1.375 ;
        RECT  1.580 1.145 1.840 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.255 0.755 4.345 1.060 ;
        RECT  4.265 0.185 4.340 0.380 ;
        RECT  4.165 0.300 4.265 0.380 ;
        RECT  4.165 0.755 4.255 0.920 ;
        RECT  3.580 0.300 3.815 0.380 ;
        RECT  3.580 0.755 3.815 0.910 ;
        RECT  3.505 0.185 3.580 0.380 ;
        RECT  3.505 0.755 3.580 1.040 ;
        RECT  3.390 0.545 3.700 0.635 ;
        RECT  3.320 0.350 3.390 0.765 ;
        RECT  2.535 0.350 3.320 0.420 ;
        RECT  3.215 0.695 3.320 0.765 ;
        RECT  2.450 0.210 3.230 0.280 ;
        RECT  3.105 0.695 3.215 1.075 ;
        RECT  2.305 0.545 3.205 0.615 ;
        RECT  2.655 0.695 3.105 0.765 ;
        RECT  2.545 0.695 2.655 1.075 ;
        RECT  2.375 0.210 2.450 0.345 ;
        RECT  2.235 0.215 2.305 0.615 ;
        RECT  1.390 0.215 2.235 0.285 ;
        RECT  1.895 0.355 2.155 0.425 ;
        RECT  2.065 0.845 2.135 1.050 ;
        RECT  1.895 0.845 2.065 0.915 ;
        RECT  1.825 0.355 1.895 0.915 ;
        RECT  1.800 0.520 1.825 0.655 ;
        RECT  1.730 0.355 1.755 0.465 ;
        RECT  1.660 0.355 1.730 1.040 ;
        RECT  0.895 0.880 1.660 0.950 ;
        RECT  1.320 0.215 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD6BWP40

MACRO CKLNQD8BWP40
    CLASS CORE ;
    FOREIGN CKLNQD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN TE
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.840 0.185 4.925 0.455 ;
        RECT  4.840 0.755 4.925 1.060 ;
        RECT  4.540 0.350 4.840 0.455 ;
        RECT  4.545 0.755 4.840 0.920 ;
        RECT  4.515 0.755 4.545 1.060 ;
        RECT  4.515 0.185 4.540 0.455 ;
        RECT  4.465 0.185 4.515 1.060 ;
        RECT  4.455 0.350 4.465 1.060 ;
        RECT  4.165 0.350 4.455 0.920 ;
        RECT  4.160 0.350 4.165 0.455 ;
        RECT  4.160 0.755 4.165 0.920 ;
        RECT  4.080 0.185 4.160 0.455 ;
        RECT  4.080 0.755 4.160 1.035 ;
        RECT  3.780 0.350 4.080 0.455 ;
        RECT  3.780 0.755 4.080 0.910 ;
        RECT  3.705 0.185 3.780 0.455 ;
        RECT  3.705 0.755 3.780 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.475 0.405 0.905 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.096200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.125 0.770 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 -0.115 5.180 0.115 ;
        RECT  5.025 -0.115 5.110 0.460 ;
        RECT  4.745 -0.115 5.025 0.115 ;
        RECT  4.635 -0.115 4.745 0.270 ;
        RECT  4.365 -0.115 4.635 0.115 ;
        RECT  4.255 -0.115 4.365 0.270 ;
        RECT  3.975 -0.115 4.255 0.115 ;
        RECT  3.880 -0.115 3.975 0.245 ;
        RECT  3.590 -0.115 3.880 0.115 ;
        RECT  3.515 -0.115 3.590 0.260 ;
        RECT  3.255 -0.115 3.515 0.115 ;
        RECT  3.095 -0.115 3.255 0.140 ;
        RECT  2.000 -0.115 3.095 0.115 ;
        RECT  1.880 -0.115 2.000 0.120 ;
        RECT  1.595 -0.115 1.880 0.115 ;
        RECT  1.480 -0.115 1.595 0.145 ;
        RECT  1.200 -0.115 1.480 0.115 ;
        RECT  1.130 -0.115 1.200 0.295 ;
        RECT  0.350 -0.115 1.130 0.115 ;
        RECT  0.230 -0.115 0.350 0.235 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.145 5.180 1.375 ;
        RECT  5.035 0.720 5.120 1.375 ;
        RECT  4.745 1.145 5.035 1.375 ;
        RECT  4.645 1.005 4.745 1.375 ;
        RECT  4.350 1.145 4.645 1.375 ;
        RECT  4.275 1.005 4.350 1.375 ;
        RECT  3.975 1.145 4.275 1.375 ;
        RECT  3.885 0.985 3.975 1.375 ;
        RECT  3.600 1.145 3.885 1.375 ;
        RECT  3.500 0.855 3.600 1.375 ;
        RECT  3.205 1.145 3.500 1.375 ;
        RECT  3.130 0.855 3.205 1.375 ;
        RECT  2.825 1.145 3.130 1.375 ;
        RECT  2.750 0.865 2.825 1.375 ;
        RECT  2.435 1.145 2.750 1.375 ;
        RECT  2.355 0.875 2.435 1.375 ;
        RECT  1.960 1.145 2.355 1.375 ;
        RECT  1.840 0.985 1.960 1.375 ;
        RECT  1.580 1.145 1.840 1.375 ;
        RECT  1.460 1.020 1.580 1.375 ;
        RECT  1.170 1.145 1.460 1.375 ;
        RECT  1.050 1.020 1.170 1.375 ;
        RECT  0.130 1.145 1.050 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.840 0.185 4.925 0.455 ;
        RECT  4.840 0.755 4.925 1.060 ;
        RECT  4.585 0.350 4.840 0.455 ;
        RECT  4.585 0.755 4.840 0.920 ;
        RECT  4.080 0.185 4.095 0.455 ;
        RECT  4.080 0.755 4.095 1.035 ;
        RECT  3.780 0.350 4.080 0.455 ;
        RECT  3.780 0.755 4.080 0.910 ;
        RECT  3.705 0.185 3.780 0.455 ;
        RECT  3.705 0.755 3.780 1.040 ;
        RECT  3.625 0.535 3.935 0.625 ;
        RECT  3.555 0.350 3.625 0.765 ;
        RECT  2.445 0.350 3.555 0.420 ;
        RECT  3.400 0.695 3.555 0.765 ;
        RECT  2.540 0.210 3.430 0.280 ;
        RECT  3.315 0.695 3.400 1.075 ;
        RECT  3.025 0.695 3.315 0.765 ;
        RECT  2.305 0.545 3.300 0.615 ;
        RECT  2.940 0.695 3.025 1.075 ;
        RECT  2.650 0.695 2.940 0.765 ;
        RECT  2.540 0.695 2.650 1.075 ;
        RECT  2.375 0.300 2.445 0.420 ;
        RECT  2.235 0.215 2.305 0.615 ;
        RECT  1.390 0.215 2.235 0.285 ;
        RECT  1.895 0.355 2.155 0.425 ;
        RECT  2.065 0.845 2.135 1.050 ;
        RECT  1.895 0.845 2.065 0.915 ;
        RECT  1.825 0.355 1.895 0.915 ;
        RECT  1.800 0.520 1.825 0.655 ;
        RECT  1.730 0.355 1.755 0.465 ;
        RECT  1.660 0.355 1.730 1.040 ;
        RECT  0.895 0.880 1.660 0.950 ;
        RECT  1.320 0.215 1.390 0.810 ;
        RECT  1.055 0.740 1.320 0.810 ;
        RECT  1.170 0.395 1.240 0.630 ;
        RECT  1.060 0.395 1.170 0.465 ;
        RECT  0.980 0.245 1.060 0.465 ;
        RECT  0.975 0.595 1.055 0.810 ;
        RECT  0.720 0.245 0.980 0.315 ;
        RECT  0.895 0.395 0.910 0.515 ;
        RECT  0.825 0.395 0.895 1.055 ;
        RECT  0.570 0.985 0.825 1.055 ;
        RECT  0.650 0.245 0.720 0.905 ;
        RECT  0.500 0.595 0.570 1.055 ;
        RECT  0.465 0.220 0.545 0.375 ;
        RECT  0.130 0.305 0.465 0.375 ;
        RECT  0.050 0.220 0.130 0.375 ;
    END
END CKLNQD8BWP40

MACRO CKMUX2D1BWP40
    CLASS CORE ;
    FOREIGN CKMUX2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.148000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.215 1.505 1.030 ;
        RECT  1.310 0.215 1.425 0.315 ;
        RECT  1.355 0.930 1.425 1.030 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.041000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.021200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.405 0.520 0.430 0.640 ;
        RECT  0.315 0.355 0.405 0.790 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.540 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.540 1.375 ;
        RECT  1.120 1.000 1.220 1.375 ;
        RECT  0.340 1.145 1.120 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.205 0.515 1.285 0.925 ;
        RECT  0.790 0.850 1.205 0.925 ;
        RECT  0.940 0.195 1.040 0.275 ;
        RECT  0.940 0.710 1.040 0.780 ;
        RECT  0.860 0.195 0.940 0.780 ;
        RECT  0.770 0.995 0.940 1.075 ;
        RECT  0.690 0.335 0.790 0.925 ;
        RECT  0.580 0.995 0.770 1.065 ;
        RECT  0.510 0.315 0.580 0.800 ;
        RECT  0.510 0.870 0.580 1.065 ;
        RECT  0.125 0.870 0.510 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END CKMUX2D1BWP40

MACRO CKMUX2D2BWP40
    CLASS CORE ;
    FOREIGN CKMUX2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.385 1.925 0.775 ;
        RECT  1.770 0.385 1.850 0.465 ;
        RECT  1.770 0.695 1.850 0.775 ;
        RECT  1.700 0.215 1.770 0.465 ;
        RECT  1.700 0.695 1.770 1.060 ;
        RECT  1.610 0.215 1.700 0.315 ;
        RECT  1.650 0.900 1.700 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.035000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.026000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.038400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.840 -0.115 1.910 0.275 ;
        RECT  1.540 -0.115 1.840 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.250 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.840 0.965 1.910 1.375 ;
        RECT  1.540 1.145 1.840 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 0.545 1.750 0.615 ;
        RECT  1.500 0.545 1.580 0.925 ;
        RECT  1.085 0.850 1.500 0.925 ;
        RECT  1.225 0.195 1.360 0.275 ;
        RECT  1.225 0.710 1.360 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.155 0.195 1.225 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.010 0.310 1.085 0.925 ;
        RECT  0.830 0.320 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.320 0.830 0.390 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.320 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END CKMUX2D2BWP40

MACRO CKMUX2D4BWP40
    CLASS CORE ;
    FOREIGN CKMUX2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.215 2.570 0.435 ;
        RECT  2.480 0.785 2.550 1.060 ;
        RECT  2.415 0.785 2.480 0.905 ;
        RECT  2.415 0.355 2.470 0.435 ;
        RECT  2.205 0.355 2.415 0.905 ;
        RECT  2.170 0.355 2.205 0.435 ;
        RECT  2.160 0.785 2.205 0.905 ;
        RECT  2.070 0.215 2.170 0.435 ;
        RECT  2.090 0.785 2.160 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.455 0.245 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.027200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.345 1.645 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.510 0.835 0.610 ;
        RECT  0.315 0.510 0.385 0.765 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.680 -0.115 2.750 0.455 ;
        RECT  2.385 -0.115 2.680 0.115 ;
        RECT  2.275 -0.115 2.385 0.265 ;
        RECT  1.970 -0.115 2.275 0.115 ;
        RECT  1.900 -0.115 1.970 0.425 ;
        RECT  1.615 -0.115 1.900 0.115 ;
        RECT  1.505 -0.115 1.615 0.260 ;
        RECT  0.780 -0.115 1.505 0.115 ;
        RECT  0.660 -0.115 0.780 0.295 ;
        RECT  0.345 -0.115 0.660 0.115 ;
        RECT  0.275 -0.115 0.345 0.350 ;
        RECT  0.000 -0.115 0.275 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.680 0.720 2.750 1.375 ;
        RECT  2.385 1.145 2.680 1.375 ;
        RECT  2.275 0.985 2.385 1.375 ;
        RECT  1.990 1.145 2.275 1.375 ;
        RECT  1.865 0.995 1.990 1.375 ;
        RECT  1.610 1.145 1.865 1.375 ;
        RECT  1.510 1.000 1.610 1.375 ;
        RECT  0.780 1.145 1.510 1.375 ;
        RECT  0.660 1.010 0.780 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.215 2.570 0.435 ;
        RECT  2.485 0.785 2.550 1.060 ;
        RECT  2.070 0.215 2.135 0.435 ;
        RECT  2.090 0.785 2.135 1.060 ;
        RECT  2.020 0.515 2.080 0.645 ;
        RECT  1.940 0.515 2.020 0.925 ;
        RECT  1.180 0.850 1.940 0.925 ;
        RECT  1.795 0.670 1.820 0.780 ;
        RECT  1.715 0.245 1.795 0.780 ;
        RECT  1.330 0.710 1.715 0.780 ;
        RECT  1.330 0.195 1.405 0.275 ;
        RECT  1.250 0.195 1.330 0.780 ;
        RECT  1.160 0.995 1.330 1.075 ;
        RECT  1.080 0.335 1.180 0.925 ;
        RECT  0.970 0.995 1.160 1.065 ;
        RECT  0.940 0.365 1.010 0.800 ;
        RECT  0.900 0.870 0.970 1.065 ;
        RECT  0.465 0.365 0.940 0.440 ;
        RECT  0.465 0.710 0.940 0.800 ;
        RECT  0.125 0.870 0.900 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END CKMUX2D4BWP40

MACRO CKMUX2D8BWP40
    CLASS CORE ;
    FOREIGN CKMUX2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.512000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.215 3.970 0.435 ;
        RECT  3.880 0.785 3.950 1.060 ;
        RECT  3.560 0.785 3.880 0.905 ;
        RECT  3.570 0.355 3.870 0.435 ;
        RECT  3.470 0.215 3.570 0.435 ;
        RECT  3.490 0.785 3.560 1.060 ;
        RECT  3.395 0.785 3.490 0.905 ;
        RECT  3.395 0.355 3.470 0.435 ;
        RECT  3.190 0.355 3.395 0.905 ;
        RECT  3.185 0.215 3.190 0.905 ;
        RECT  3.090 0.215 3.185 0.435 ;
        RECT  3.170 0.785 3.185 0.905 ;
        RECT  3.100 0.785 3.170 1.060 ;
        RECT  2.750 0.785 3.100 0.905 ;
        RECT  2.760 0.355 3.090 0.435 ;
        RECT  2.660 0.215 2.760 0.435 ;
        RECT  2.680 0.785 2.750 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.057000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.455 0.245 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.046800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.120 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.041400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.810 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.080 -0.115 4.150 0.450 ;
        RECT  3.785 -0.115 4.080 0.115 ;
        RECT  3.675 -0.115 3.785 0.265 ;
        RECT  3.370 -0.115 3.675 0.115 ;
        RECT  3.300 -0.115 3.370 0.265 ;
        RECT  3.005 -0.115 3.300 0.115 ;
        RECT  2.895 -0.115 3.005 0.265 ;
        RECT  2.530 -0.115 2.895 0.115 ;
        RECT  2.430 -0.115 2.530 0.275 ;
        RECT  2.090 -0.115 2.430 0.115 ;
        RECT  1.990 -0.115 2.090 0.265 ;
        RECT  0.720 -0.115 1.990 0.115 ;
        RECT  0.600 -0.115 0.720 0.280 ;
        RECT  0.320 -0.115 0.600 0.115 ;
        RECT  0.235 -0.115 0.320 0.345 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.080 0.720 4.150 1.375 ;
        RECT  3.785 1.145 4.080 1.375 ;
        RECT  3.675 0.985 3.785 1.375 ;
        RECT  3.390 1.145 3.675 1.375 ;
        RECT  3.265 0.995 3.390 1.375 ;
        RECT  3.005 1.145 3.265 1.375 ;
        RECT  2.895 0.985 3.005 1.375 ;
        RECT  2.530 1.145 2.895 1.375 ;
        RECT  2.430 1.000 2.530 1.375 ;
        RECT  2.090 1.145 2.430 1.375 ;
        RECT  1.990 1.000 2.090 1.375 ;
        RECT  0.720 1.145 1.990 1.375 ;
        RECT  0.600 1.010 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.870 0.215 3.970 0.435 ;
        RECT  3.880 0.785 3.950 1.060 ;
        RECT  3.560 0.785 3.880 0.905 ;
        RECT  3.570 0.355 3.870 0.435 ;
        RECT  3.470 0.215 3.570 0.435 ;
        RECT  3.490 0.785 3.560 1.060 ;
        RECT  3.465 0.785 3.490 0.905 ;
        RECT  3.465 0.355 3.470 0.435 ;
        RECT  3.090 0.215 3.115 0.435 ;
        RECT  3.100 0.785 3.115 1.060 ;
        RECT  2.750 0.785 3.100 0.905 ;
        RECT  2.760 0.355 3.090 0.435 ;
        RECT  2.660 0.215 2.760 0.435 ;
        RECT  2.680 0.785 2.750 1.060 ;
        RECT  2.570 0.515 3.075 0.645 ;
        RECT  2.490 0.515 2.570 0.925 ;
        RECT  1.445 0.855 2.490 0.925 ;
        RECT  2.275 0.705 2.320 0.780 ;
        RECT  2.190 0.345 2.275 0.780 ;
        RECT  1.575 0.345 2.190 0.415 ;
        RECT  1.530 0.710 2.190 0.780 ;
        RECT  1.445 0.195 1.895 0.265 ;
        RECT  0.890 0.995 1.620 1.065 ;
        RECT  1.375 0.195 1.445 0.925 ;
        RECT  0.970 0.195 1.375 0.265 ;
        RECT  0.970 0.855 1.375 0.925 ;
        RECT  1.215 0.350 1.285 0.785 ;
        RECT  0.405 0.350 1.215 0.425 ;
        RECT  0.405 0.710 1.215 0.785 ;
        RECT  0.820 0.870 0.890 1.065 ;
        RECT  0.125 0.870 0.820 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END CKMUX2D8BWP40

MACRO CKND10BWP40
    CLASS CORE ;
    FOREIGN CKND10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.510000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.405 0.695 1.505 1.045 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.155 0.300 1.405 0.465 ;
        RECT  1.155 0.695 1.405 0.885 ;
        RECT  1.095 0.300 1.155 0.885 ;
        RECT  1.015 0.185 1.095 1.045 ;
        RECT  0.945 0.300 1.015 0.885 ;
        RECT  0.715 0.300 0.945 0.465 ;
        RECT  0.715 0.695 0.945 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.272000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.840 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 -0.115 2.100 0.115 ;
        RECT  1.975 -0.115 2.045 0.335 ;
        RECT  1.690 -0.115 1.975 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.290 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.685 2.050 1.375 ;
        RECT  1.690 1.145 1.970 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.405 0.695 1.505 1.045 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.225 0.300 1.405 0.465 ;
        RECT  1.225 0.695 1.405 0.885 ;
        RECT  0.715 0.300 0.875 0.465 ;
        RECT  0.715 0.695 0.875 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END CKND10BWP40

MACRO CKND12BWP40
    CLASS CORE ;
    FOREIGN CKND12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.612000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.435 0.695 1.505 1.045 ;
        RECT  1.435 0.185 1.475 0.465 ;
        RECT  1.405 0.185 1.435 1.045 ;
        RECT  1.095 0.300 1.405 0.885 ;
        RECT  1.085 0.185 1.095 1.035 ;
        RECT  1.025 0.185 1.085 0.465 ;
        RECT  1.025 0.695 1.085 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.326400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.855 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.425 -0.115 2.520 0.115 ;
        RECT  2.355 -0.115 2.425 0.325 ;
        RECT  2.070 -0.115 2.355 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.310 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 1.145 2.520 1.375 ;
        RECT  2.355 0.670 2.435 1.375 ;
        RECT  2.070 1.145 2.355 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.505 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  0.715 0.300 1.015 0.465 ;
        RECT  0.715 0.695 1.015 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END CKND12BWP40

MACRO CKND14BWP40
    CLASS CORE ;
    FOREIGN CKND14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.737800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.595 0.300 1.785 0.465 ;
        RECT  1.595 0.695 1.785 0.885 ;
        RECT  1.505 0.300 1.595 0.885 ;
        RECT  1.475 0.300 1.505 1.045 ;
        RECT  1.405 0.185 1.475 1.045 ;
        RECT  1.225 0.300 1.405 0.885 ;
        RECT  1.095 0.300 1.225 0.465 ;
        RECT  1.095 0.695 1.225 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.380800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.045 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 2.940 0.115 ;
        RECT  2.750 -0.115 2.840 0.350 ;
        RECT  2.450 -0.115 2.750 0.115 ;
        RECT  2.330 -0.115 2.450 0.230 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.315 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.845 1.145 2.940 1.375 ;
        RECT  2.755 0.685 2.845 1.375 ;
        RECT  2.450 1.145 2.755 1.375 ;
        RECT  2.330 0.955 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.645 0.300 1.785 0.465 ;
        RECT  1.645 0.695 1.785 0.885 ;
        RECT  1.095 0.300 1.155 0.465 ;
        RECT  1.095 0.695 1.155 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END CKND14BWP40

MACRO CKND16BWP40
    CLASS CORE ;
    FOREIGN CKND16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.816000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.715 0.300 1.765 0.465 ;
        RECT  1.715 0.695 1.765 0.885 ;
        RECT  1.505 0.300 1.715 0.885 ;
        RECT  1.455 0.300 1.505 1.045 ;
        RECT  1.385 0.185 1.455 1.045 ;
        RECT  1.365 0.300 1.385 0.885 ;
        RECT  1.075 0.300 1.365 0.465 ;
        RECT  1.075 0.695 1.365 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.435200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.260 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.335 ;
        RECT  2.810 -0.115 3.095 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.685 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.785 0.185 1.835 0.465 ;
        RECT  1.785 0.695 1.835 1.035 ;
        RECT  1.075 0.300 1.295 0.465 ;
        RECT  1.075 0.695 1.295 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END CKND16BWP40

MACRO CKND18BWP40
    CLASS CORE ;
    FOREIGN CKND18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.918000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.995 0.300 2.145 0.465 ;
        RECT  1.995 0.695 2.145 0.885 ;
        RECT  1.835 0.300 1.995 0.885 ;
        RECT  1.765 0.185 1.835 1.045 ;
        RECT  1.715 0.300 1.765 1.045 ;
        RECT  1.645 0.300 1.715 0.885 ;
        RECT  1.455 0.300 1.645 0.465 ;
        RECT  1.505 0.695 1.645 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.489600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.565 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 -0.115 3.640 0.115 ;
        RECT  3.515 -0.115 3.585 0.330 ;
        RECT  3.190 -0.115 3.515 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.685 3.590 1.375 ;
        RECT  3.190 1.145 3.510 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.645 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.645 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  2.065 0.300 2.145 0.465 ;
        RECT  2.060 0.695 2.145 0.885 ;
        RECT  1.455 0.300 1.575 0.465 ;
        RECT  1.505 0.695 1.575 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END CKND18BWP40

MACRO CKND1BWP40
    CLASS CORE ;
    FOREIGN CKND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.091000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.185 0.385 1.045 ;
        RECT  0.280 0.185 0.315 0.425 ;
        RECT  0.290 0.710 0.315 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.026000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.080 -0.115 0.150 0.295 ;
        RECT  0.000 -0.115 0.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.145 0.420 1.375 ;
        RECT  0.080 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.080 1.375 ;
        END
    END VDD
END CKND1BWP40

MACRO CKND20BWP40
    CLASS CORE ;
    FOREIGN CKND20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.047200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.275 0.300 2.525 0.465 ;
        RECT  2.275 0.695 2.525 0.885 ;
        RECT  2.215 0.300 2.275 0.885 ;
        RECT  2.135 0.185 2.215 1.045 ;
        RECT  1.925 0.300 2.135 0.885 ;
        RECT  1.835 0.300 1.925 0.465 ;
        RECT  1.835 0.695 1.925 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.505 0.695 1.765 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.544000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.050 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.320 ;
        RECT  3.570 -0.115 3.935 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.685 4.010 1.375 ;
        RECT  3.570 1.145 3.930 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.345 0.300 2.525 0.465 ;
        RECT  2.345 0.695 2.525 0.885 ;
        RECT  1.835 0.300 1.855 0.465 ;
        RECT  1.835 0.695 1.855 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.505 0.695 1.765 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END CKND20BWP40

MACRO CKND24BWP40
    CLASS CORE ;
    FOREIGN CKND24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.224000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.555 0.185 2.595 0.465 ;
        RECT  2.555 0.695 2.595 1.035 ;
        RECT  2.525 0.185 2.555 1.035 ;
        RECT  2.215 0.300 2.525 0.885 ;
        RECT  2.205 0.185 2.215 1.045 ;
        RECT  2.135 0.185 2.205 0.465 ;
        RECT  2.135 0.695 2.205 1.045 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.652800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.815 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.115 4.760 0.115 ;
        RECT  4.600 -0.115 4.700 0.360 ;
        RECT  4.330 -0.115 4.600 0.115 ;
        RECT  4.210 -0.115 4.330 0.230 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.230 ;
        RECT  3.570 -0.115 3.830 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.320 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 1.145 4.760 1.375 ;
        RECT  4.600 0.695 4.700 1.375 ;
        RECT  4.330 1.145 4.600 1.375 ;
        RECT  4.210 0.955 4.330 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 0.955 3.950 1.375 ;
        RECT  3.570 1.145 3.830 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.955 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.625 0.300 2.905 0.465 ;
        RECT  2.625 0.695 2.905 0.885 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END CKND24BWP40

MACRO CKND2BWP40
    CLASS CORE ;
    FOREIGN CKND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.100500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.335 0.385 0.815 ;
        RECT  0.315 0.185 0.320 0.815 ;
        RECT  0.225 0.185 0.315 0.425 ;
        RECT  0.245 0.735 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.053600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.280 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.295 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 0.560 1.375 ;
        RECT  0.430 0.910 0.510 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END CKND2BWP40

MACRO CKND2D1BWP40
    CLASS CORE ;
    FOREIGN CKND2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.106250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.435 0.215 0.455 0.385 ;
        RECT  0.315 0.845 0.455 0.915 ;
        RECT  0.245 0.845 0.315 1.050 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.560 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.145 0.560 1.375 ;
        RECT  0.410 0.985 0.520 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END CKND2D1BWP40

MACRO CKND2D2BWP40
    CLASS CORE ;
    FOREIGN CKND2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.181500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.835 0.720 1.035 ;
        RECT  0.390 0.835 0.640 0.915 ;
        RECT  0.355 0.345 0.390 0.915 ;
        RECT  0.315 0.345 0.355 1.045 ;
        RECT  0.240 0.345 0.315 0.415 ;
        RECT  0.260 0.705 0.315 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.495 0.815 0.765 ;
        RECT  0.595 0.495 0.730 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.980 0.115 ;
        RECT  0.630 -0.115 0.730 0.275 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.835 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.440 0.990 0.540 1.375 ;
        RECT  0.145 1.145 0.440 1.375 ;
        RECT  0.075 0.705 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 0.255 0.910 0.415 ;
        RECT  0.550 0.345 0.830 0.415 ;
        RECT  0.480 0.205 0.550 0.415 ;
        RECT  0.035 0.205 0.480 0.275 ;
    END
END CKND2D2BWP40

MACRO CKND2D4BWP40
    CLASS CORE ;
    FOREIGN CKND2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.375000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.735 1.575 1.045 ;
        RECT  1.430 0.345 1.435 1.045 ;
        RECT  1.365 0.345 1.430 0.945 ;
        RECT  1.250 0.345 1.365 0.415 ;
        RECT  1.160 0.845 1.365 0.945 ;
        RECT  1.080 0.845 1.160 1.075 ;
        RECT  0.720 0.845 1.080 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.585 0.495 1.645 0.640 ;
        RECT  1.515 0.195 1.585 0.640 ;
        RECT  1.155 0.195 1.515 0.265 ;
        RECT  1.085 0.195 1.155 0.415 ;
        RECT  0.950 0.345 1.085 0.415 ;
        RECT  0.850 0.345 0.950 0.630 ;
        RECT  0.715 0.345 0.850 0.415 ;
        RECT  0.645 0.195 0.715 0.415 ;
        RECT  0.290 0.195 0.645 0.265 ;
        RECT  0.210 0.195 0.290 0.625 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.270 0.625 ;
        RECT  1.080 0.495 1.155 0.775 ;
        RECT  0.675 0.705 1.080 0.775 ;
        RECT  0.585 0.495 0.675 0.775 ;
        RECT  0.560 0.495 0.585 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 -0.115 1.820 0.115 ;
        RECT  1.680 -0.115 1.780 0.415 ;
        RECT  0.960 -0.115 1.680 0.115 ;
        RECT  0.840 -0.115 0.960 0.275 ;
        RECT  0.120 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.120 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.145 1.820 1.375 ;
        RECT  1.680 0.990 1.780 1.375 ;
        RECT  1.360 1.145 1.680 1.375 ;
        RECT  1.260 1.030 1.360 1.375 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.840 0.985 0.960 1.375 ;
        RECT  0.550 1.145 0.840 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.345 1.295 0.415 ;
        RECT  1.160 0.845 1.295 0.945 ;
        RECT  1.080 0.845 1.160 1.075 ;
        RECT  0.720 0.845 1.080 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
    END
END CKND2D4BWP40

MACRO CKND2D8BWP40
    CLASS CORE ;
    FOREIGN CKND2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.603600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
        RECT  1.995 0.845 2.770 0.915 ;
        RECT  1.995 0.345 2.050 0.425 ;
        RECT  1.900 0.345 1.995 0.915 ;
        RECT  1.840 0.495 1.900 0.915 ;
        RECT  1.785 0.495 1.840 1.045 ;
        RECT  1.760 0.735 1.785 1.045 ;
        RECT  1.460 0.735 1.760 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  0.440 0.845 1.270 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.208000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.000 0.495 3.185 0.625 ;
        RECT  2.930 0.205 3.000 0.625 ;
        RECT  2.590 0.205 2.930 0.275 ;
        RECT  2.510 0.205 2.590 0.415 ;
        RECT  2.445 0.345 2.510 0.415 ;
        RECT  2.345 0.345 2.445 0.635 ;
        RECT  2.230 0.345 2.345 0.415 ;
        RECT  2.150 0.205 2.230 0.415 ;
        RECT  1.790 0.205 2.150 0.275 ;
        RECT  1.715 0.205 1.790 0.410 ;
        RECT  1.645 0.340 1.715 0.410 ;
        RECT  1.560 0.340 1.645 0.640 ;
        RECT  1.505 0.340 1.560 0.410 ;
        RECT  1.435 0.205 1.505 0.410 ;
        RECT  1.070 0.205 1.435 0.275 ;
        RECT  0.990 0.205 1.070 0.415 ;
        RECT  0.845 0.345 0.990 0.415 ;
        RECT  0.735 0.345 0.845 0.635 ;
        RECT  0.710 0.345 0.735 0.415 ;
        RECT  0.630 0.205 0.710 0.415 ;
        RECT  0.290 0.205 0.630 0.275 ;
        RECT  0.220 0.205 0.290 0.640 ;
        RECT  0.160 0.495 0.220 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.208000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.665 0.705 1.015 0.775 ;
        RECT  0.525 0.495 0.665 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 -0.115 3.220 0.115 ;
        RECT  3.080 -0.115 3.180 0.415 ;
        RECT  2.420 -0.115 3.080 0.115 ;
        RECT  2.320 -0.115 2.420 0.275 ;
        RECT  1.645 -0.115 2.320 0.115 ;
        RECT  1.575 -0.115 1.645 0.260 ;
        RECT  0.900 -0.115 1.575 0.115 ;
        RECT  0.800 -0.115 0.900 0.275 ;
        RECT  0.140 -0.115 0.800 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.755 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 0.985 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.985 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.985 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.025 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.985 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.790 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
        RECT  2.065 0.845 2.770 0.915 ;
        RECT  1.460 0.735 1.715 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  0.440 0.845 1.270 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.495 2.595 0.775 ;
        RECT  2.215 0.705 2.525 0.775 ;
        RECT  2.145 0.495 2.215 0.775 ;
        RECT  2.070 0.495 2.145 0.640 ;
    END
END CKND2D8BWP40

MACRO CKND3BWP40
    CLASS CORE ;
    FOREIGN CKND3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.214400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.655 0.185 0.735 0.445 ;
        RECT  0.665 0.735 0.735 1.045 ;
        RECT  0.525 0.735 0.665 0.815 ;
        RECT  0.525 0.355 0.655 0.445 ;
        RECT  0.455 0.355 0.525 0.815 ;
        RECT  0.320 0.355 0.455 0.445 ;
        RECT  0.315 0.735 0.455 0.815 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.735 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.080400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.840 0.115 ;
        RECT  0.430 -0.115 0.510 0.285 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 0.840 1.375 ;
        RECT  0.430 0.885 0.510 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END CKND3BWP40

MACRO CKND4BWP40
    CLASS CORE ;
    FOREIGN CKND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.201000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.660 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.595 0.705 0.665 0.820 ;
        RECT  0.595 0.310 0.660 0.445 ;
        RECT  0.385 0.310 0.595 0.820 ;
        RECT  0.320 0.310 0.385 0.445 ;
        RECT  0.315 0.705 0.385 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.107200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.335 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.695 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END CKND4BWP40

MACRO CKND5BWP40
    CLASS CORE ;
    FOREIGN CKND5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.304850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.735 0.705 1.105 0.820 ;
        RECT  0.740 0.310 1.100 0.445 ;
        RECT  0.735 0.185 0.740 0.445 ;
        RECT  0.665 0.185 0.735 1.030 ;
        RECT  0.660 0.185 0.665 0.820 ;
        RECT  0.525 0.310 0.660 0.820 ;
        RECT  0.320 0.310 0.525 0.445 ;
        RECT  0.315 0.705 0.525 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.134000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.445 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.980 -0.115 1.260 0.115 ;
        RECT  0.860 -0.115 0.980 0.240 ;
        RECT  0.560 -0.115 0.860 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.145 1.260 1.375 ;
        RECT  0.850 0.890 0.970 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.805 0.705 1.105 0.820 ;
        RECT  0.805 0.310 1.100 0.445 ;
        RECT  0.320 0.310 0.455 0.445 ;
        RECT  0.315 0.705 0.455 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END CKND5BWP40

MACRO CKND6BWP40
    CLASS CORE ;
    FOREIGN CKND6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.301500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.875 0.705 1.045 0.820 ;
        RECT  0.875 0.310 1.040 0.445 ;
        RECT  0.740 0.310 0.875 0.820 ;
        RECT  0.735 0.185 0.740 0.820 ;
        RECT  0.665 0.185 0.735 1.030 ;
        RECT  0.660 0.185 0.665 0.445 ;
        RECT  0.315 0.705 0.665 0.820 ;
        RECT  0.320 0.310 0.660 0.445 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.160800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.515 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.115 1.400 0.115 ;
        RECT  1.210 -0.115 1.330 0.240 ;
        RECT  0.950 -0.115 1.210 0.115 ;
        RECT  0.830 -0.115 0.950 0.240 ;
        RECT  0.560 -0.115 0.830 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.320 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.400 1.375 ;
        RECT  1.210 0.750 1.330 1.375 ;
        RECT  0.960 1.145 1.210 1.375 ;
        RECT  0.830 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.830 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.945 0.705 1.045 0.820 ;
        RECT  0.945 0.310 1.040 0.445 ;
        RECT  0.320 0.310 0.595 0.445 ;
        RECT  0.315 0.705 0.595 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END CKND6BWP40

MACRO CKND8BWP40
    CLASS CORE ;
    FOREIGN CKND8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.431800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.015 0.185 1.095 0.445 ;
        RECT  1.020 0.705 1.090 1.030 ;
        RECT  1.015 0.705 1.020 0.820 ;
        RECT  0.700 0.310 1.015 0.820 ;
        RECT  0.695 0.185 0.700 0.820 ;
        RECT  0.665 0.185 0.695 1.030 ;
        RECT  0.620 0.185 0.665 0.445 ;
        RECT  0.625 0.705 0.665 1.030 ;
        RECT  0.315 0.705 0.625 0.820 ;
        RECT  0.320 0.310 0.620 0.445 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.217600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 -0.115 1.820 0.115 ;
        RECT  1.665 -0.115 1.750 0.345 ;
        RECT  1.305 -0.115 1.665 0.115 ;
        RECT  1.185 -0.115 1.305 0.240 ;
        RECT  0.910 -0.115 1.185 0.115 ;
        RECT  0.790 -0.115 0.910 0.240 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.240 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.145 1.820 1.375 ;
        RECT  1.670 0.725 1.780 1.375 ;
        RECT  1.310 1.145 1.670 1.375 ;
        RECT  1.190 0.890 1.310 1.375 ;
        RECT  0.915 1.145 1.190 1.375 ;
        RECT  0.795 0.890 0.915 1.375 ;
        RECT  0.530 1.145 0.795 1.375 ;
        RECT  0.410 0.890 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.085 0.185 1.095 0.445 ;
        RECT  1.085 0.705 1.090 1.030 ;
        RECT  0.320 0.310 0.595 0.445 ;
        RECT  0.315 0.705 0.595 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END CKND8BWP40

MACRO CKNR2D1BWP40
    CLASS CORE ;
    FOREIGN CKNR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.183350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.715 1.365 1.075 ;
        RECT  0.955 0.715 1.270 0.815 ;
        RECT  0.865 0.325 0.955 0.815 ;
        RECT  0.765 0.325 0.865 0.395 ;
        RECT  0.635 0.210 0.765 0.395 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.065600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.595 0.625 ;
        RECT  0.175 0.355 0.245 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.065600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.365 0.625 ;
        RECT  1.025 0.495 1.295 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 -0.115 1.400 0.115 ;
        RECT  0.870 -0.115 0.950 0.255 ;
        RECT  0.540 -0.115 0.870 0.115 ;
        RECT  0.440 -0.115 0.540 0.415 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 1.400 1.375 ;
        RECT  0.430 0.890 0.550 1.375 ;
        RECT  0.145 1.145 0.430 1.375 ;
        RECT  0.075 0.720 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.755 0.995 1.160 1.065 ;
        RECT  0.645 0.705 0.755 1.065 ;
        RECT  0.355 0.705 0.645 0.785 ;
        RECT  0.240 0.705 0.355 1.065 ;
    END
END CKNR2D1BWP40

MACRO CKNR2D2BWP40
    CLASS CORE ;
    FOREIGN CKNR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.269550 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.215 2.065 1.065 ;
        RECT  1.365 0.215 1.995 0.345 ;
        RECT  1.970 0.635 1.995 1.065 ;
        RECT  1.285 0.215 1.365 0.915 ;
        RECT  0.440 0.215 1.285 0.285 ;
        RECT  1.200 0.845 1.285 0.915 ;
        RECT  0.440 0.845 0.550 0.915 ;
        RECT  0.360 0.215 0.440 0.915 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.109200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.510 0.495 1.785 0.640 ;
        RECT  1.435 0.495 1.510 1.065 ;
        RECT  1.105 0.995 1.435 1.065 ;
        RECT  1.015 0.750 1.105 1.065 ;
        RECT  0.945 0.750 1.015 0.820 ;
        RECT  0.840 0.495 0.945 0.820 ;
        RECT  0.715 0.750 0.840 0.820 ;
        RECT  0.645 0.750 0.715 1.065 ;
        RECT  0.290 0.995 0.645 1.065 ;
        RECT  0.210 0.495 0.290 1.065 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.112400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.495 1.175 0.640 ;
        RECT  1.015 0.355 1.105 0.640 ;
        RECT  0.675 0.355 1.015 0.425 ;
        RECT  0.585 0.355 0.675 0.640 ;
        RECT  0.560 0.495 0.585 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 2.100 0.115 ;
        RECT  1.200 -0.115 1.320 0.145 ;
        RECT  0.930 -0.115 1.200 0.115 ;
        RECT  0.810 -0.115 0.930 0.145 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.140 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.675 1.145 2.100 1.375 ;
        RECT  1.605 0.735 1.675 1.375 ;
        RECT  0.930 1.145 1.605 1.375 ;
        RECT  0.810 0.890 0.930 1.375 ;
        RECT  0.130 1.145 0.810 1.375 ;
        RECT  0.050 0.705 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END CKNR2D2BWP40

MACRO CKNR2D4BWP40
    CLASS CORE ;
    FOREIGN CKNR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.585000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 0.210 4.515 0.370 ;
        RECT  4.340 0.210 4.420 0.915 ;
        RECT  3.480 0.210 4.340 0.280 ;
        RECT  4.230 0.845 4.340 0.915 ;
        RECT  3.480 0.845 3.570 0.915 ;
        RECT  3.410 0.210 3.480 0.915 ;
        RECT  2.850 0.210 3.410 0.280 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  1.995 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.995 0.835 2.065 0.915 ;
        RECT  1.910 0.210 1.995 0.915 ;
        RECT  1.785 0.210 1.910 0.625 ;
        RECT  1.350 0.210 1.785 0.280 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.264000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 0.495 4.655 0.640 ;
        RECT  4.490 0.495 4.570 1.065 ;
        RECT  4.135 0.995 4.490 1.065 ;
        RECT  4.065 0.710 4.135 1.065 ;
        RECT  3.940 0.710 4.065 0.780 ;
        RECT  3.815 0.495 3.940 0.780 ;
        RECT  3.745 0.710 3.815 0.780 ;
        RECT  3.665 0.710 3.745 1.065 ;
        RECT  3.330 0.995 3.665 1.065 ;
        RECT  3.255 0.495 3.330 1.065 ;
        RECT  3.000 0.495 3.255 0.625 ;
        RECT  2.930 0.495 3.000 1.055 ;
        RECT  2.590 0.985 2.930 1.055 ;
        RECT  2.510 0.745 2.590 1.055 ;
        RECT  2.445 0.745 2.510 0.815 ;
        RECT  2.345 0.525 2.445 0.815 ;
        RECT  2.230 0.745 2.345 0.815 ;
        RECT  2.135 0.745 2.230 1.065 ;
        RECT  1.790 0.995 2.135 1.065 ;
        RECT  1.715 0.710 1.790 1.065 ;
        RECT  1.655 0.710 1.715 0.780 ;
        RECT  1.575 0.495 1.655 0.780 ;
        RECT  1.505 0.710 1.575 0.780 ;
        RECT  1.435 0.710 1.505 1.055 ;
        RECT  1.085 0.985 1.435 1.055 ;
        RECT  0.990 0.745 1.085 1.055 ;
        RECT  0.845 0.745 0.990 0.815 ;
        RECT  0.735 0.495 0.845 0.815 ;
        RECT  0.710 0.745 0.735 0.815 ;
        RECT  0.630 0.745 0.710 1.055 ;
        RECT  0.290 0.985 0.630 1.055 ;
        RECT  0.220 0.495 0.290 1.055 ;
        RECT  0.125 0.495 0.220 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.264000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.350 1.085 0.625 ;
        RECT  0.665 0.350 1.015 0.420 ;
        RECT  0.525 0.350 0.665 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.720 -0.115 4.760 0.115 ;
        RECT  4.620 -0.115 4.720 0.415 ;
        RECT  4.350 -0.115 4.620 0.115 ;
        RECT  4.230 -0.115 4.350 0.140 ;
        RECT  3.960 -0.115 4.230 0.115 ;
        RECT  3.840 -0.115 3.960 0.140 ;
        RECT  0.910 -0.115 3.840 0.115 ;
        RECT  0.790 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.640 0.720 4.710 1.375 ;
        RECT  3.960 1.145 4.640 1.375 ;
        RECT  3.840 0.860 3.960 1.375 ;
        RECT  3.180 1.145 3.840 1.375 ;
        RECT  3.080 0.745 3.180 1.375 ;
        RECT  2.420 1.145 3.080 1.375 ;
        RECT  2.320 0.885 2.420 1.375 ;
        RECT  1.645 1.145 2.320 1.375 ;
        RECT  1.575 0.860 1.645 1.375 ;
        RECT  0.900 1.145 1.575 1.375 ;
        RECT  0.800 0.885 0.900 1.375 ;
        RECT  0.140 1.145 0.800 1.375 ;
        RECT  0.040 0.725 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.420 0.210 4.515 0.370 ;
        RECT  4.340 0.210 4.420 0.915 ;
        RECT  3.480 0.210 4.340 0.280 ;
        RECT  4.230 0.845 4.340 0.915 ;
        RECT  3.480 0.845 3.570 0.915 ;
        RECT  3.410 0.210 3.480 0.915 ;
        RECT  2.850 0.210 3.410 0.280 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  2.065 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.350 0.210 1.715 0.280 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        RECT  4.195 0.520 4.220 0.640 ;
        RECT  4.105 0.350 4.195 0.640 ;
        RECT  3.725 0.350 4.105 0.420 ;
        RECT  3.650 0.350 3.725 0.630 ;
        RECT  3.550 0.510 3.650 0.630 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.350 2.595 0.640 ;
        RECT  2.215 0.350 2.525 0.420 ;
        RECT  2.145 0.350 2.215 0.665 ;
        RECT  2.070 0.495 2.145 0.665 ;
    END
END CKNR2D4BWP40

MACRO CKNR2D8BWP40
    CLASS CORE ;
    FOREIGN CKNR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.176000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.010 0.210 9.145 0.395 ;
        RECT  8.940 0.210 9.010 0.915 ;
        RECT  8.080 0.210 8.940 0.285 ;
        RECT  8.850 0.845 8.940 0.915 ;
        RECT  8.080 0.845 8.190 0.915 ;
        RECT  8.000 0.210 8.080 0.915 ;
        RECT  7.470 0.210 8.000 0.370 ;
        RECT  7.390 0.210 7.470 0.915 ;
        RECT  6.560 0.210 7.390 0.280 ;
        RECT  7.310 0.845 7.390 0.915 ;
        RECT  6.560 0.845 6.650 0.915 ;
        RECT  6.490 0.210 6.560 0.915 ;
        RECT  5.930 0.210 6.490 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.075 0.210 5.850 0.280 ;
        RECT  5.770 0.835 5.850 0.915 ;
        RECT  5.075 0.835 5.145 0.915 ;
        RECT  4.990 0.210 5.075 0.915 ;
        RECT  4.865 0.210 4.990 0.625 ;
        RECT  4.430 0.210 4.865 0.350 ;
        RECT  4.350 0.210 4.430 0.915 ;
        RECT  3.520 0.210 4.350 0.280 ;
        RECT  4.250 0.835 4.350 0.915 ;
        RECT  3.520 0.835 3.610 0.915 ;
        RECT  3.440 0.210 3.520 0.915 ;
        RECT  2.895 0.210 3.440 0.370 ;
        RECT  2.825 0.210 2.895 0.915 ;
        RECT  1.960 0.210 2.825 0.285 ;
        RECT  2.730 0.845 2.825 0.915 ;
        RECT  1.960 0.845 2.070 0.915 ;
        RECT  1.880 0.210 1.960 0.915 ;
        RECT  1.355 0.210 1.880 0.375 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.170 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.528000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.170 0.495 9.320 0.625 ;
        RECT  9.100 0.495 9.170 1.065 ;
        RECT  8.755 0.995 9.100 1.065 ;
        RECT  8.685 0.720 8.755 1.065 ;
        RECT  8.550 0.720 8.685 0.790 ;
        RECT  8.435 0.495 8.550 0.790 ;
        RECT  8.365 0.720 8.435 0.790 ;
        RECT  8.285 0.720 8.365 1.065 ;
        RECT  7.930 0.995 8.285 1.065 ;
        RECT  7.850 0.495 7.930 1.065 ;
        RECT  7.630 0.495 7.850 0.625 ;
        RECT  7.550 0.495 7.630 1.065 ;
        RECT  7.215 0.995 7.550 1.065 ;
        RECT  7.145 0.745 7.215 1.065 ;
        RECT  7.020 0.745 7.145 0.815 ;
        RECT  6.895 0.495 7.020 0.815 ;
        RECT  6.825 0.745 6.895 0.815 ;
        RECT  6.745 0.745 6.825 1.065 ;
        RECT  6.410 0.995 6.745 1.065 ;
        RECT  6.335 0.495 6.410 1.065 ;
        RECT  6.080 0.495 6.335 0.625 ;
        RECT  6.010 0.495 6.080 1.055 ;
        RECT  5.670 0.985 6.010 1.055 ;
        RECT  5.590 0.745 5.670 1.055 ;
        RECT  5.525 0.745 5.590 0.815 ;
        RECT  5.425 0.525 5.525 0.815 ;
        RECT  5.310 0.745 5.425 0.815 ;
        RECT  5.215 0.745 5.310 1.065 ;
        RECT  4.870 0.995 5.215 1.065 ;
        RECT  4.795 0.710 4.870 1.065 ;
        RECT  4.735 0.710 4.795 0.780 ;
        RECT  4.655 0.495 4.735 0.780 ;
        RECT  4.585 0.710 4.655 0.780 ;
        RECT  4.515 0.710 4.585 1.055 ;
        RECT  4.165 0.985 4.515 1.055 ;
        RECT  4.070 0.745 4.165 1.055 ;
        RECT  3.925 0.745 4.070 0.815 ;
        RECT  3.815 0.495 3.925 0.815 ;
        RECT  3.790 0.745 3.815 0.815 ;
        RECT  3.710 0.745 3.790 1.055 ;
        RECT  3.370 0.985 3.710 1.055 ;
        RECT  3.300 0.495 3.370 1.055 ;
        RECT  3.055 0.495 3.300 0.665 ;
        RECT  2.975 0.495 3.055 1.065 ;
        RECT  2.635 0.995 2.975 1.065 ;
        RECT  2.555 0.720 2.635 1.065 ;
        RECT  2.485 0.720 2.555 0.790 ;
        RECT  2.275 0.495 2.485 0.790 ;
        RECT  2.235 0.720 2.275 0.790 ;
        RECT  2.165 0.720 2.235 1.065 ;
        RECT  1.810 0.995 2.165 1.065 ;
        RECT  1.730 0.495 1.810 1.065 ;
        RECT  1.515 0.495 1.730 0.625 ;
        RECT  1.430 0.495 1.515 1.065 ;
        RECT  1.085 0.995 1.430 1.065 ;
        RECT  1.015 0.720 1.085 1.065 ;
        RECT  0.905 0.720 1.015 0.790 ;
        RECT  0.805 0.495 0.905 0.790 ;
        RECT  0.695 0.720 0.805 0.790 ;
        RECT  0.625 0.720 0.695 1.065 ;
        RECT  0.270 0.995 0.625 1.065 ;
        RECT  0.190 0.495 0.270 1.065 ;
        RECT  0.070 0.495 0.190 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.528000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.280 0.625 ;
        RECT  4.095 0.350 4.165 0.625 ;
        RECT  3.745 0.350 4.095 0.420 ;
        RECT  3.605 0.350 3.745 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.340 -0.115 9.380 0.115 ;
        RECT  9.240 -0.115 9.340 0.410 ;
        RECT  8.970 -0.115 9.240 0.115 ;
        RECT  8.850 -0.115 8.970 0.140 ;
        RECT  8.585 -0.115 8.850 0.115 ;
        RECT  8.445 -0.115 8.585 0.140 ;
        RECT  7.430 -0.115 8.445 0.115 ;
        RECT  7.310 -0.115 7.430 0.140 ;
        RECT  7.040 -0.115 7.310 0.115 ;
        RECT  6.920 -0.115 7.040 0.140 ;
        RECT  6.650 -0.115 6.920 0.115 ;
        RECT  6.530 -0.115 6.650 0.140 ;
        RECT  2.850 -0.115 6.530 0.115 ;
        RECT  2.730 -0.115 2.850 0.140 ;
        RECT  2.460 -0.115 2.730 0.115 ;
        RECT  2.330 -0.115 2.460 0.140 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.140 ;
        RECT  0.910 -0.115 1.950 0.115 ;
        RECT  0.785 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.785 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.325 1.145 9.380 1.375 ;
        RECT  9.255 0.720 9.325 1.375 ;
        RECT  8.580 1.145 9.255 1.375 ;
        RECT  8.460 0.860 8.580 1.375 ;
        RECT  7.780 1.145 8.460 1.375 ;
        RECT  7.710 0.715 7.780 1.375 ;
        RECT  7.040 1.145 7.710 1.375 ;
        RECT  6.920 0.885 7.040 1.375 ;
        RECT  6.260 1.145 6.920 1.375 ;
        RECT  6.160 0.740 6.260 1.375 ;
        RECT  5.500 1.145 6.160 1.375 ;
        RECT  5.400 0.885 5.500 1.375 ;
        RECT  4.725 1.145 5.400 1.375 ;
        RECT  4.655 0.860 4.725 1.375 ;
        RECT  3.980 1.145 4.655 1.375 ;
        RECT  3.880 0.885 3.980 1.375 ;
        RECT  3.210 1.145 3.880 1.375 ;
        RECT  3.140 0.735 3.210 1.375 ;
        RECT  2.460 1.145 3.140 1.375 ;
        RECT  2.340 0.870 2.460 1.375 ;
        RECT  1.660 1.145 2.340 1.375 ;
        RECT  1.590 0.705 1.660 1.375 ;
        RECT  0.910 1.145 1.590 1.375 ;
        RECT  0.790 0.860 0.910 1.375 ;
        RECT  0.120 1.145 0.790 1.375 ;
        RECT  0.050 0.720 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.010 0.210 9.145 0.395 ;
        RECT  8.940 0.210 9.010 0.915 ;
        RECT  8.080 0.210 8.940 0.285 ;
        RECT  8.850 0.845 8.940 0.915 ;
        RECT  8.080 0.845 8.190 0.915 ;
        RECT  8.000 0.210 8.080 0.915 ;
        RECT  7.470 0.210 8.000 0.370 ;
        RECT  7.390 0.210 7.470 0.915 ;
        RECT  6.560 0.210 7.390 0.280 ;
        RECT  7.310 0.845 7.390 0.915 ;
        RECT  6.560 0.845 6.650 0.915 ;
        RECT  6.490 0.210 6.560 0.915 ;
        RECT  5.930 0.210 6.490 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.145 0.210 5.850 0.280 ;
        RECT  5.770 0.835 5.850 0.915 ;
        RECT  4.430 0.210 4.795 0.350 ;
        RECT  4.350 0.210 4.430 0.915 ;
        RECT  3.520 0.210 4.350 0.280 ;
        RECT  4.250 0.835 4.350 0.915 ;
        RECT  3.520 0.835 3.610 0.915 ;
        RECT  3.440 0.210 3.520 0.915 ;
        RECT  2.895 0.210 3.440 0.370 ;
        RECT  2.825 0.210 2.895 0.915 ;
        RECT  1.960 0.210 2.825 0.285 ;
        RECT  2.730 0.845 2.825 0.915 ;
        RECT  1.960 0.845 2.070 0.915 ;
        RECT  1.880 0.210 1.960 0.915 ;
        RECT  1.355 0.210 1.880 0.375 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.170 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        RECT  8.755 0.495 8.825 0.640 ;
        RECT  8.680 0.355 8.755 0.640 ;
        RECT  8.315 0.355 8.680 0.425 ;
        RECT  8.225 0.355 8.315 0.640 ;
        RECT  8.200 0.495 8.225 0.640 ;
        RECT  7.275 0.520 7.300 0.665 ;
        RECT  7.185 0.350 7.275 0.665 ;
        RECT  6.805 0.350 7.185 0.420 ;
        RECT  6.730 0.350 6.805 0.630 ;
        RECT  6.630 0.510 6.730 0.630 ;
        RECT  5.675 0.495 5.775 0.640 ;
        RECT  5.605 0.350 5.675 0.640 ;
        RECT  5.295 0.350 5.605 0.420 ;
        RECT  5.225 0.350 5.295 0.665 ;
        RECT  5.150 0.495 5.225 0.665 ;
        RECT  2.640 0.495 2.705 0.640 ;
        RECT  2.565 0.355 2.640 0.640 ;
        RECT  2.190 0.355 2.565 0.425 ;
        RECT  2.105 0.355 2.190 0.640 ;
        RECT  2.080 0.495 2.105 0.640 ;
        RECT  1.085 0.495 1.155 0.640 ;
        RECT  1.010 0.355 1.085 0.640 ;
        RECT  0.655 0.355 1.010 0.425 ;
        RECT  0.565 0.355 0.655 0.640 ;
        RECT  0.540 0.495 0.565 0.640 ;
    END
END CKNR2D8BWP40

MACRO CKOR2D1BWP40
    CLASS CORE ;
    FOREIGN CKOR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.144000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.195 1.225 1.075 ;
        RECT  1.110 0.195 1.155 0.445 ;
        RECT  1.125 0.685 1.155 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.495 0.770 0.785 ;
        RECT  0.245 0.715 0.695 0.785 ;
        RECT  0.170 0.495 0.245 0.785 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.625 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.115 1.260 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.510 -0.115 0.800 0.115 ;
        RECT  0.430 -0.115 0.510 0.255 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 1.260 1.375 ;
        RECT  0.810 1.030 0.910 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.050 0.940 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 1.025 0.640 ;
        RECT  0.850 0.345 0.920 0.925 ;
        RECT  0.705 0.345 0.850 0.415 ;
        RECT  0.415 0.855 0.850 0.925 ;
        RECT  0.220 0.995 0.715 1.065 ;
        RECT  0.620 0.230 0.705 0.415 ;
    END
END CKOR2D1BWP40

MACRO CKOR2D2BWP40
    CLASS CORE ;
    FOREIGN CKOR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.235 0.905 ;
        RECT  1.095 0.355 1.155 0.435 ;
        RECT  1.095 0.785 1.155 0.905 ;
        RECT  1.025 0.215 1.095 0.435 ;
        RECT  1.015 0.785 1.095 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.040000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.495 0.770 0.785 ;
        RECT  0.245 0.715 0.695 0.785 ;
        RECT  0.170 0.495 0.245 0.785 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.043600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.625 0.640 ;
        RECT  0.315 0.355 0.385 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.115 1.400 0.115 ;
        RECT  1.250 -0.115 1.330 0.280 ;
        RECT  0.920 -0.115 1.250 0.115 ;
        RECT  0.800 -0.115 0.920 0.275 ;
        RECT  0.510 -0.115 0.800 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.400 1.375 ;
        RECT  1.250 0.980 1.330 1.375 ;
        RECT  0.910 1.145 1.250 1.375 ;
        RECT  0.810 1.030 0.910 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.050 0.865 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.520 1.000 0.640 ;
        RECT  0.850 0.345 0.920 0.925 ;
        RECT  0.705 0.345 0.850 0.415 ;
        RECT  0.415 0.855 0.850 0.925 ;
        RECT  0.220 0.995 0.715 1.065 ;
        RECT  0.620 0.240 0.705 0.415 ;
    END
END CKOR2D2BWP40

MACRO CKOR2D4BWP40
    CLASS CORE ;
    FOREIGN CKOR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.284000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 0.445 ;
        RECT  1.855 0.700 1.925 1.045 ;
        RECT  1.830 0.185 1.855 1.045 ;
        RECT  1.645 0.325 1.830 0.820 ;
        RECT  1.500 0.325 1.645 0.445 ;
        RECT  1.500 0.700 1.645 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.069600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.490 1.160 0.765 ;
        RECT  0.535 0.695 1.015 0.765 ;
        RECT  0.445 0.495 0.535 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.069600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.540 0.915 0.625 ;
        RECT  0.730 0.355 0.815 0.625 ;
        RECT  0.300 0.355 0.730 0.425 ;
        RECT  0.220 0.355 0.300 0.650 ;
        RECT  0.125 0.495 0.220 0.650 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.175 -0.115 2.240 0.115 ;
        RECT  2.055 -0.115 2.175 0.415 ;
        RECT  1.720 -0.115 2.055 0.115 ;
        RECT  1.600 -0.115 1.720 0.255 ;
        RECT  1.330 -0.115 1.600 0.115 ;
        RECT  1.190 -0.115 1.330 0.235 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.145 ;
        RECT  0.540 -0.115 0.810 0.115 ;
        RECT  0.420 -0.115 0.540 0.255 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.175 1.145 2.240 1.375 ;
        RECT  2.055 0.745 2.175 1.375 ;
        RECT  1.720 1.145 2.055 1.375 ;
        RECT  1.600 0.890 1.720 1.375 ;
        RECT  1.300 1.145 1.600 1.375 ;
        RECT  1.220 0.995 1.300 1.375 ;
        RECT  0.540 1.145 1.220 1.375 ;
        RECT  0.420 1.000 0.540 1.375 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.500 0.325 1.575 0.445 ;
        RECT  1.500 0.700 1.575 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        RECT  1.320 0.545 1.565 0.615 ;
        RECT  1.250 0.325 1.320 0.915 ;
        RECT  1.040 0.325 1.250 0.395 ;
        RECT  0.905 0.845 1.250 0.915 ;
        RECT  0.970 0.215 1.040 0.395 ;
        RECT  0.620 0.215 0.970 0.285 ;
        RECT  0.835 0.845 0.905 1.075 ;
        RECT  0.145 0.845 0.835 0.915 ;
        RECT  0.035 0.845 0.145 1.075 ;
    END
END CKOR2D4BWP40

MACRO CKOR2D8BWP40
    CLASS CORE ;
    FOREIGN CKOR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.185 3.820 0.445 ;
        RECT  3.740 0.700 3.820 0.990 ;
        RECT  3.420 0.325 3.740 0.445 ;
        RECT  3.420 0.700 3.740 0.820 ;
        RECT  3.340 0.185 3.420 0.445 ;
        RECT  3.340 0.700 3.420 0.990 ;
        RECT  3.255 0.325 3.340 0.445 ;
        RECT  3.255 0.700 3.340 0.820 ;
        RECT  3.045 0.325 3.255 0.820 ;
        RECT  3.020 0.325 3.045 0.445 ;
        RECT  3.020 0.700 3.045 0.820 ;
        RECT  2.925 0.185 3.020 0.445 ;
        RECT  2.925 0.700 3.020 1.045 ;
        RECT  2.620 0.325 2.925 0.445 ;
        RECT  2.620 0.700 2.925 0.820 ;
        RECT  2.540 0.185 2.620 0.445 ;
        RECT  2.540 0.700 2.620 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.147600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.495 2.295 0.625 ;
        RECT  1.435 0.355 1.530 0.625 ;
        RECT  0.245 0.355 1.435 0.425 ;
        RECT  0.135 0.355 0.245 0.645 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.147600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 1.325 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.445 ;
        RECT  3.640 -0.115 3.930 0.115 ;
        RECT  3.520 -0.115 3.640 0.255 ;
        RECT  3.240 -0.115 3.520 0.115 ;
        RECT  3.120 -0.115 3.240 0.255 ;
        RECT  2.840 -0.115 3.120 0.115 ;
        RECT  2.720 -0.115 2.840 0.255 ;
        RECT  2.430 -0.115 2.720 0.115 ;
        RECT  2.350 -0.115 2.430 0.275 ;
        RECT  2.025 -0.115 2.350 0.115 ;
        RECT  1.955 -0.115 2.025 0.255 ;
        RECT  1.290 -0.115 1.955 0.115 ;
        RECT  1.170 -0.115 1.290 0.145 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.145 ;
        RECT  0.000 -0.115 0.790 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.700 4.010 1.375 ;
        RECT  3.640 1.145 3.930 1.375 ;
        RECT  3.520 0.890 3.640 1.375 ;
        RECT  3.240 1.145 3.520 1.375 ;
        RECT  3.120 0.890 3.240 1.375 ;
        RECT  2.840 1.145 3.120 1.375 ;
        RECT  2.720 0.890 2.840 1.375 ;
        RECT  2.430 1.145 2.720 1.375 ;
        RECT  2.350 0.880 2.430 1.375 ;
        RECT  2.050 1.145 2.350 1.375 ;
        RECT  1.970 0.985 2.050 1.375 ;
        RECT  1.655 1.145 1.970 1.375 ;
        RECT  1.565 0.985 1.655 1.375 ;
        RECT  0.125 1.145 1.565 1.375 ;
        RECT  0.055 0.720 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.740 0.185 3.820 0.445 ;
        RECT  3.740 0.700 3.820 0.990 ;
        RECT  3.420 0.325 3.740 0.445 ;
        RECT  3.420 0.700 3.740 0.820 ;
        RECT  3.340 0.185 3.420 0.445 ;
        RECT  3.340 0.700 3.420 0.990 ;
        RECT  3.325 0.325 3.340 0.445 ;
        RECT  3.325 0.700 3.340 0.820 ;
        RECT  2.925 0.185 2.975 0.445 ;
        RECT  2.925 0.700 2.975 1.045 ;
        RECT  2.620 0.325 2.925 0.445 ;
        RECT  2.620 0.700 2.925 0.820 ;
        RECT  2.540 0.185 2.620 0.445 ;
        RECT  2.540 0.700 2.620 0.990 ;
        RECT  2.445 0.545 2.895 0.615 ;
        RECT  2.375 0.345 2.445 0.765 ;
        RECT  2.235 0.345 2.375 0.415 ;
        RECT  0.410 0.695 2.375 0.765 ;
        RECT  2.165 0.845 2.255 1.075 ;
        RECT  2.165 0.185 2.235 0.415 ;
        RECT  1.835 0.345 2.165 0.415 ;
        RECT  1.835 0.845 2.165 0.915 ;
        RECT  1.765 0.215 1.835 0.415 ;
        RECT  1.765 0.845 1.835 1.075 ;
        RECT  0.600 0.215 1.765 0.285 ;
        RECT  1.455 0.845 1.765 0.915 ;
        RECT  1.385 0.845 1.455 1.075 ;
        RECT  1.075 0.845 1.385 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.335 0.845 0.625 0.915 ;
        RECT  0.220 0.845 0.335 1.075 ;
    END
END CKOR2D8BWP40

MACRO CKXOR2D1BWP40
    CLASS CORE ;
    FOREIGN CKXOR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.050 ;
        RECT  1.415 0.185 1.435 0.435 ;
        RECT  1.410 0.870 1.435 1.050 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.355 1.225 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.047600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.780 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 -0.115 1.540 0.115 ;
        RECT  1.185 -0.115 1.265 0.275 ;
        RECT  0.270 -0.115 1.185 0.115 ;
        RECT  0.270 0.345 0.340 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.150 1.135 1.300 1.375 ;
        RECT  0.340 1.145 1.150 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.520 1.365 0.810 ;
        RECT  1.235 0.740 1.295 0.810 ;
        RECT  1.165 0.740 1.235 1.065 ;
        RECT  0.805 0.995 1.165 1.065 ;
        RECT  0.950 0.195 1.020 0.925 ;
        RECT  0.340 0.195 0.950 0.265 ;
        RECT  0.725 0.350 0.805 1.065 ;
        RECT  0.545 0.860 0.635 1.070 ;
        RECT  0.465 0.355 0.565 0.790 ;
        RECT  0.125 0.860 0.545 0.930 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.280 0.120 0.420 ;
        RECT  0.035 0.280 0.105 1.040 ;
    END
END CKXOR2D1BWP40

MACRO CKXOR2D2BWP40
    CLASS CORE ;
    FOREIGN CKXOR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.355 2.205 0.905 ;
        RECT  1.975 0.355 2.125 0.430 ;
        RECT  1.975 0.780 2.125 0.905 ;
        RECT  1.905 0.205 1.975 0.430 ;
        RECT  1.905 0.780 1.975 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.355 0.385 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.034600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.685 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.180 -0.115 2.240 0.115 ;
        RECT  2.080 -0.115 2.180 0.275 ;
        RECT  1.810 -0.115 2.080 0.115 ;
        RECT  1.715 -0.115 1.810 0.415 ;
        RECT  0.620 -0.115 1.715 0.115 ;
        RECT  0.500 -0.115 0.620 0.140 ;
        RECT  0.000 -0.115 0.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.180 1.145 2.240 1.375 ;
        RECT  2.080 0.985 2.180 1.375 ;
        RECT  1.810 1.145 2.080 1.375 ;
        RECT  1.690 1.130 1.810 1.375 ;
        RECT  0.615 1.145 1.690 1.375 ;
        RECT  0.505 0.865 0.615 1.375 ;
        RECT  0.175 1.145 0.505 1.375 ;
        RECT  0.065 0.830 0.175 1.375 ;
        RECT  0.000 1.145 0.065 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.755 0.540 1.825 1.060 ;
        RECT  0.960 0.990 1.755 1.060 ;
        RECT  1.440 0.350 1.630 0.420 ;
        RECT  1.440 0.840 1.620 0.910 ;
        RECT  1.350 0.350 1.440 0.910 ;
        RECT  1.105 0.210 1.185 0.920 ;
        RECT  0.665 0.210 1.105 0.280 ;
        RECT  0.960 0.400 1.015 0.470 ;
        RECT  0.890 0.400 0.960 1.060 ;
        RECT  0.735 0.360 0.805 0.970 ;
        RECT  0.595 0.210 0.665 0.775 ;
        RECT  0.310 0.210 0.595 0.280 ;
        RECT  0.420 0.705 0.595 0.775 ;
        RECT  0.330 0.705 0.420 1.075 ;
        RECT  1.825 0.540 2.025 0.610 ;
    END
END CKXOR2D2BWP40

MACRO CKXOR2D4BWP40
    CLASS CORE ;
    FOREIGN CKXOR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 0.205 2.835 1.065 ;
        RECT  2.755 0.355 2.765 1.065 ;
        RECT  2.625 0.355 2.755 0.915 ;
        RECT  2.455 0.355 2.625 0.475 ;
        RECT  2.455 0.780 2.625 0.915 ;
        RECT  2.385 0.205 2.455 0.475 ;
        RECT  2.385 0.780 2.455 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.074000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.485 0.530 0.635 ;
        RECT  0.035 0.355 0.105 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.034600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.105 0.665 2.160 0.765 ;
        RECT  1.995 0.495 2.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 -0.115 3.080 0.115 ;
        RECT  2.940 -0.115 3.040 0.445 ;
        RECT  2.660 -0.115 2.940 0.115 ;
        RECT  2.560 -0.115 2.660 0.285 ;
        RECT  2.280 -0.115 2.560 0.115 ;
        RECT  2.160 -0.115 2.280 0.265 ;
        RECT  1.100 -0.115 2.160 0.115 ;
        RECT  0.980 -0.115 1.100 0.140 ;
        RECT  0.680 -0.115 0.980 0.115 ;
        RECT  0.560 -0.115 0.680 0.140 ;
        RECT  0.180 -0.115 0.560 0.115 ;
        RECT  0.070 -0.115 0.180 0.275 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.145 3.080 1.375 ;
        RECT  2.940 0.705 3.040 1.375 ;
        RECT  2.670 1.145 2.940 1.375 ;
        RECT  2.550 0.995 2.670 1.375 ;
        RECT  2.280 1.145 2.550 1.375 ;
        RECT  2.160 1.130 2.280 1.375 ;
        RECT  1.100 1.145 2.160 1.375 ;
        RECT  0.980 1.005 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 0.890 0.720 1.375 ;
        RECT  0.330 1.145 0.600 1.375 ;
        RECT  0.230 0.890 0.330 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.455 0.355 2.555 0.475 ;
        RECT  2.455 0.780 2.555 0.915 ;
        RECT  2.385 0.205 2.455 0.475 ;
        RECT  2.385 0.780 2.455 1.065 ;
        RECT  2.305 0.545 2.445 0.615 ;
        RECT  2.235 0.545 2.305 1.060 ;
        RECT  1.425 0.990 2.235 1.060 ;
        RECT  1.870 0.350 2.100 0.420 ;
        RECT  1.870 0.850 2.100 0.920 ;
        RECT  1.800 0.350 1.870 0.920 ;
        RECT  1.600 0.210 1.680 0.905 ;
        RECT  0.690 0.210 1.600 0.280 ;
        RECT  1.425 0.400 1.520 0.470 ;
        RECT  1.355 0.400 1.425 1.060 ;
        RECT  1.025 0.360 1.280 0.470 ;
        RECT  1.175 0.810 1.265 1.065 ;
        RECT  1.025 0.810 1.175 0.880 ;
        RECT  0.940 0.360 1.025 0.880 ;
        RECT  0.790 0.360 0.940 0.440 ;
        RECT  0.905 0.810 0.940 0.880 ;
        RECT  0.805 0.810 0.905 1.015 ;
        RECT  0.690 0.510 0.870 0.640 ;
        RECT  0.610 0.210 0.690 0.820 ;
        RECT  0.340 0.210 0.610 0.370 ;
        RECT  0.520 0.750 0.610 0.820 ;
        RECT  0.430 0.750 0.520 1.075 ;
        RECT  0.055 0.750 0.130 1.075 ;
        RECT  0.130 0.750 0.430 0.820 ;
    END
END CKXOR2D4BWP40

MACRO CKXOR2D8BWP40
    CLASS CORE ;
    FOREIGN CKXOR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.468000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.205 4.795 0.485 ;
        RECT  4.725 0.780 4.795 1.065 ;
        RECT  4.415 0.355 4.725 0.485 ;
        RECT  4.425 0.780 4.725 0.905 ;
        RECT  4.345 0.780 4.425 1.065 ;
        RECT  4.345 0.205 4.415 0.485 ;
        RECT  4.235 0.355 4.345 0.485 ;
        RECT  4.235 0.780 4.345 0.905 ;
        RECT  4.030 0.355 4.235 0.905 ;
        RECT  4.025 0.205 4.030 1.065 ;
        RECT  3.960 0.205 4.025 0.480 ;
        RECT  3.955 0.780 4.025 1.065 ;
        RECT  3.650 0.355 3.960 0.480 ;
        RECT  3.650 0.780 3.955 0.905 ;
        RECT  3.580 0.195 3.650 0.480 ;
        RECT  3.580 0.780 3.650 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.855 0.625 ;
        RECT  0.175 0.355 0.245 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.056200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.220 0.495 3.335 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.000 -0.115 5.040 0.115 ;
        RECT  4.900 -0.115 5.000 0.485 ;
        RECT  4.620 -0.115 4.900 0.115 ;
        RECT  4.520 -0.115 4.620 0.275 ;
        RECT  4.240 -0.115 4.520 0.115 ;
        RECT  4.140 -0.115 4.240 0.275 ;
        RECT  3.855 -0.115 4.140 0.115 ;
        RECT  3.755 -0.115 3.855 0.275 ;
        RECT  3.475 -0.115 3.755 0.115 ;
        RECT  3.355 -0.115 3.475 0.250 ;
        RECT  1.485 -0.115 3.355 0.115 ;
        RECT  1.360 -0.115 1.485 0.245 ;
        RECT  1.100 -0.115 1.360 0.115 ;
        RECT  0.980 -0.115 1.100 0.215 ;
        RECT  0.725 -0.115 0.980 0.115 ;
        RECT  0.595 -0.115 0.725 0.240 ;
        RECT  0.000 -0.115 0.595 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.000 1.145 5.040 1.375 ;
        RECT  4.900 0.705 5.000 1.375 ;
        RECT  4.620 1.145 4.900 1.375 ;
        RECT  4.520 0.985 4.620 1.375 ;
        RECT  4.240 1.145 4.520 1.375 ;
        RECT  4.140 0.985 4.240 1.375 ;
        RECT  3.855 1.145 4.140 1.375 ;
        RECT  3.755 0.985 3.855 1.375 ;
        RECT  3.475 1.145 3.755 1.375 ;
        RECT  3.355 1.130 3.475 1.375 ;
        RECT  1.840 1.145 3.355 1.375 ;
        RECT  1.765 0.850 1.840 1.375 ;
        RECT  1.460 1.145 1.765 1.375 ;
        RECT  1.380 0.850 1.460 1.375 ;
        RECT  1.095 1.145 1.380 1.375 ;
        RECT  0.985 0.880 1.095 1.375 ;
        RECT  0.705 1.145 0.985 1.375 ;
        RECT  0.620 0.880 0.705 1.375 ;
        RECT  0.325 1.145 0.620 1.375 ;
        RECT  0.240 0.880 0.325 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.205 4.795 0.485 ;
        RECT  4.725 0.780 4.795 1.065 ;
        RECT  4.415 0.355 4.725 0.485 ;
        RECT  4.425 0.780 4.725 0.905 ;
        RECT  4.345 0.780 4.425 1.065 ;
        RECT  4.345 0.205 4.415 0.485 ;
        RECT  4.305 0.355 4.345 0.485 ;
        RECT  4.305 0.780 4.345 0.905 ;
        RECT  3.650 0.355 3.955 0.480 ;
        RECT  3.650 0.780 3.955 0.905 ;
        RECT  3.580 0.195 3.650 0.480 ;
        RECT  3.580 0.780 3.650 1.065 ;
        RECT  3.500 0.550 3.915 0.625 ;
        RECT  3.430 0.550 3.500 1.060 ;
        RECT  2.975 0.990 3.430 1.060 ;
        RECT  3.125 0.350 3.295 0.420 ;
        RECT  3.125 0.850 3.295 0.920 ;
        RECT  3.055 0.350 3.125 0.920 ;
        RECT  2.975 0.195 3.105 0.265 ;
        RECT  2.905 0.195 2.975 1.060 ;
        RECT  2.115 0.195 2.905 0.265 ;
        RECT  2.120 0.990 2.905 1.060 ;
        RECT  2.745 0.340 2.825 0.920 ;
        RECT  1.540 0.535 2.745 0.605 ;
        RECT  1.650 0.360 2.425 0.430 ;
        RECT  2.330 0.700 2.405 0.900 ;
        RECT  2.030 0.700 2.330 0.770 ;
        RECT  1.960 0.700 2.030 1.065 ;
        RECT  1.655 0.700 1.960 0.770 ;
        RECT  1.570 0.700 1.655 1.075 ;
        RECT  1.570 0.265 1.650 0.430 ;
        RECT  1.420 0.360 1.570 0.430 ;
        RECT  1.420 0.700 1.570 0.770 ;
        RECT  1.335 0.360 1.420 0.770 ;
        RECT  1.285 0.360 1.335 0.430 ;
        RECT  1.285 0.700 1.335 0.770 ;
        RECT  1.175 0.195 1.285 0.430 ;
        RECT  1.175 0.700 1.285 1.065 ;
        RECT  1.045 0.530 1.255 0.620 ;
        RECT  0.965 0.310 1.045 0.800 ;
        RECT  0.410 0.310 0.965 0.380 ;
        RECT  0.900 0.705 0.965 0.800 ;
        RECT  0.810 0.705 0.900 1.075 ;
        RECT  0.515 0.705 0.810 0.800 ;
        RECT  0.425 0.705 0.515 1.035 ;
        RECT  0.135 0.705 0.425 0.800 ;
        RECT  0.050 0.705 0.135 1.035 ;
    END
END CKXOR2D8BWP40

MACRO DCAP16BWP40
    CLASS CORE ;
    FOREIGN DCAP16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.970 -0.115 2.240 0.115 ;
        RECT  1.890 -0.115 1.970 0.335 ;
        RECT  1.760 -0.115 1.890 0.115 ;
        RECT  1.680 -0.115 1.760 0.335 ;
        RECT  1.550 -0.115 1.680 0.115 ;
        RECT  1.470 -0.115 1.550 0.335 ;
        RECT  1.340 -0.115 1.470 0.115 ;
        RECT  1.260 -0.115 1.340 0.335 ;
        RECT  1.130 -0.115 1.260 0.115 ;
        RECT  1.050 -0.115 1.130 0.335 ;
        RECT  0.920 -0.115 1.050 0.115 ;
        RECT  0.840 -0.115 0.920 0.335 ;
        RECT  0.710 -0.115 0.840 0.115 ;
        RECT  0.630 -0.115 0.710 0.335 ;
        RECT  0.510 -0.115 0.630 0.115 ;
        RECT  0.430 -0.115 0.510 0.335 ;
        RECT  0.320 -0.115 0.430 0.115 ;
        RECT  0.240 -0.115 0.320 0.335 ;
        RECT  0.130 -0.115 0.240 0.115 ;
        RECT  0.050 -0.115 0.130 0.335 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.970 1.145 2.240 1.375 ;
        RECT  1.890 0.945 1.970 1.375 ;
        RECT  1.760 1.145 1.890 1.375 ;
        RECT  1.680 0.945 1.760 1.375 ;
        RECT  1.550 1.145 1.680 1.375 ;
        RECT  1.470 0.795 1.550 1.375 ;
        RECT  1.340 1.145 1.470 1.375 ;
        RECT  1.260 0.795 1.340 1.375 ;
        RECT  1.130 1.145 1.260 1.375 ;
        RECT  1.050 0.795 1.130 1.375 ;
        RECT  0.920 1.145 1.050 1.375 ;
        RECT  0.840 0.795 0.920 1.375 ;
        RECT  0.710 1.145 0.840 1.375 ;
        RECT  0.630 0.795 0.710 1.375 ;
        RECT  0.510 1.145 0.630 1.375 ;
        RECT  0.430 0.795 0.510 1.375 ;
        RECT  0.320 1.145 0.430 1.375 ;
        RECT  0.240 0.795 0.320 1.375 ;
        RECT  0.130 1.145 0.240 1.375 ;
        RECT  0.050 0.795 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.110 0.210 2.190 0.710 ;
        RECT  2.110 0.790 2.190 1.060 ;
        RECT  1.850 0.630 2.110 0.710 ;
        RECT  1.780 0.790 2.110 0.870 ;
        RECT  1.700 0.430 1.780 0.870 ;
        RECT  0.205 0.430 1.700 0.510 ;
    END
END DCAP16BWP40

MACRO DCAP32BWP40
    CLASS CORE ;
    FOREIGN DCAP32BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.210 -0.115 4.480 0.115 ;
        RECT  4.130 -0.115 4.210 0.335 ;
        RECT  4.000 -0.115 4.130 0.115 ;
        RECT  3.920 -0.115 4.000 0.335 ;
        RECT  3.790 -0.115 3.920 0.115 ;
        RECT  3.710 -0.115 3.790 0.335 ;
        RECT  3.580 -0.115 3.710 0.115 ;
        RECT  3.500 -0.115 3.580 0.335 ;
        RECT  3.370 -0.115 3.500 0.115 ;
        RECT  3.290 -0.115 3.370 0.335 ;
        RECT  3.160 -0.115 3.290 0.115 ;
        RECT  3.080 -0.115 3.160 0.335 ;
        RECT  2.950 -0.115 3.080 0.115 ;
        RECT  2.870 -0.115 2.950 0.335 ;
        RECT  2.750 -0.115 2.870 0.115 ;
        RECT  2.670 -0.115 2.750 0.335 ;
        RECT  2.560 -0.115 2.670 0.115 ;
        RECT  2.480 -0.115 2.560 0.335 ;
        RECT  2.370 -0.115 2.480 0.115 ;
        RECT  2.290 -0.115 2.370 0.335 ;
        RECT  2.175 -0.115 2.290 0.115 ;
        RECT  2.095 -0.115 2.175 0.335 ;
        RECT  1.970 -0.115 2.095 0.115 ;
        RECT  1.890 -0.115 1.970 0.335 ;
        RECT  1.760 -0.115 1.890 0.115 ;
        RECT  1.680 -0.115 1.760 0.335 ;
        RECT  1.550 -0.115 1.680 0.115 ;
        RECT  1.470 -0.115 1.550 0.335 ;
        RECT  1.340 -0.115 1.470 0.115 ;
        RECT  1.260 -0.115 1.340 0.335 ;
        RECT  1.130 -0.115 1.260 0.115 ;
        RECT  1.050 -0.115 1.130 0.335 ;
        RECT  0.920 -0.115 1.050 0.115 ;
        RECT  0.840 -0.115 0.920 0.335 ;
        RECT  0.710 -0.115 0.840 0.115 ;
        RECT  0.630 -0.115 0.710 0.335 ;
        RECT  0.510 -0.115 0.630 0.115 ;
        RECT  0.430 -0.115 0.510 0.335 ;
        RECT  0.320 -0.115 0.430 0.115 ;
        RECT  0.240 -0.115 0.320 0.335 ;
        RECT  0.130 -0.115 0.240 0.115 ;
        RECT  0.050 -0.115 0.130 0.335 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.210 1.145 4.480 1.375 ;
        RECT  4.130 0.945 4.210 1.375 ;
        RECT  4.000 1.145 4.130 1.375 ;
        RECT  3.920 0.945 4.000 1.375 ;
        RECT  3.790 1.145 3.920 1.375 ;
        RECT  3.710 0.795 3.790 1.375 ;
        RECT  3.580 1.145 3.710 1.375 ;
        RECT  3.500 0.795 3.580 1.375 ;
        RECT  3.370 1.145 3.500 1.375 ;
        RECT  3.290 0.795 3.370 1.375 ;
        RECT  3.160 1.145 3.290 1.375 ;
        RECT  3.080 0.795 3.160 1.375 ;
        RECT  2.950 1.145 3.080 1.375 ;
        RECT  2.870 0.795 2.950 1.375 ;
        RECT  2.750 1.145 2.870 1.375 ;
        RECT  2.670 0.795 2.750 1.375 ;
        RECT  2.560 1.145 2.670 1.375 ;
        RECT  2.480 0.795 2.560 1.375 ;
        RECT  2.370 1.145 2.480 1.375 ;
        RECT  2.290 0.795 2.370 1.375 ;
        RECT  2.175 1.145 2.290 1.375 ;
        RECT  2.095 0.795 2.175 1.375 ;
        RECT  1.970 1.145 2.095 1.375 ;
        RECT  1.890 0.795 1.970 1.375 ;
        RECT  1.760 1.145 1.890 1.375 ;
        RECT  1.680 0.795 1.760 1.375 ;
        RECT  1.550 1.145 1.680 1.375 ;
        RECT  1.470 0.795 1.550 1.375 ;
        RECT  1.340 1.145 1.470 1.375 ;
        RECT  1.260 0.795 1.340 1.375 ;
        RECT  1.130 1.145 1.260 1.375 ;
        RECT  1.050 0.795 1.130 1.375 ;
        RECT  0.920 1.145 1.050 1.375 ;
        RECT  0.840 0.795 0.920 1.375 ;
        RECT  0.710 1.145 0.840 1.375 ;
        RECT  0.630 0.795 0.710 1.375 ;
        RECT  0.510 1.145 0.630 1.375 ;
        RECT  0.430 0.795 0.510 1.375 ;
        RECT  0.320 1.145 0.430 1.375 ;
        RECT  0.240 0.795 0.320 1.375 ;
        RECT  0.130 1.145 0.240 1.375 ;
        RECT  0.050 0.795 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.350 0.210 4.430 0.710 ;
        RECT  4.350 0.790 4.430 1.060 ;
        RECT  4.090 0.630 4.350 0.710 ;
        RECT  4.020 0.790 4.350 0.870 ;
        RECT  3.940 0.430 4.020 0.870 ;
        RECT  0.205 0.430 3.940 0.510 ;
    END
END DCAP32BWP40

MACRO DCAP4BWP40
    CLASS CORE ;
    FOREIGN DCAP4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 -0.115 0.560 0.115 ;
        RECT  0.240 -0.115 0.320 0.350 ;
        RECT  0.130 -0.115 0.240 0.115 ;
        RECT  0.050 -0.115 0.130 0.350 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.145 0.560 1.375 ;
        RECT  0.240 0.945 0.320 1.375 ;
        RECT  0.130 1.145 0.240 1.375 ;
        RECT  0.050 0.945 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.430 0.210 0.510 0.700 ;
        RECT  0.430 0.785 0.510 1.075 ;
        RECT  0.320 0.620 0.430 0.700 ;
        RECT  0.225 0.785 0.430 0.865 ;
        RECT  0.155 0.440 0.225 0.865 ;
    END
END DCAP4BWP40

MACRO DCAP64BWP40
    CLASS CORE ;
    FOREIGN DCAP64BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.690 -0.115 8.960 0.115 ;
        RECT  8.610 -0.115 8.690 0.335 ;
        RECT  8.480 -0.115 8.610 0.115 ;
        RECT  8.400 -0.115 8.480 0.335 ;
        RECT  8.270 -0.115 8.400 0.115 ;
        RECT  8.190 -0.115 8.270 0.335 ;
        RECT  8.060 -0.115 8.190 0.115 ;
        RECT  7.980 -0.115 8.060 0.335 ;
        RECT  7.850 -0.115 7.980 0.115 ;
        RECT  7.770 -0.115 7.850 0.335 ;
        RECT  7.640 -0.115 7.770 0.115 ;
        RECT  7.560 -0.115 7.640 0.335 ;
        RECT  7.430 -0.115 7.560 0.115 ;
        RECT  7.350 -0.115 7.430 0.335 ;
        RECT  7.230 -0.115 7.350 0.115 ;
        RECT  7.150 -0.115 7.230 0.335 ;
        RECT  7.040 -0.115 7.150 0.115 ;
        RECT  6.960 -0.115 7.040 0.335 ;
        RECT  6.850 -0.115 6.960 0.115 ;
        RECT  6.770 -0.115 6.850 0.335 ;
        RECT  6.655 -0.115 6.770 0.115 ;
        RECT  6.575 -0.115 6.655 0.335 ;
        RECT  6.450 -0.115 6.575 0.115 ;
        RECT  6.370 -0.115 6.450 0.335 ;
        RECT  6.240 -0.115 6.370 0.115 ;
        RECT  6.160 -0.115 6.240 0.335 ;
        RECT  6.030 -0.115 6.160 0.115 ;
        RECT  5.950 -0.115 6.030 0.335 ;
        RECT  5.820 -0.115 5.950 0.115 ;
        RECT  5.740 -0.115 5.820 0.335 ;
        RECT  5.610 -0.115 5.740 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.190 -0.115 5.320 0.115 ;
        RECT  5.110 -0.115 5.190 0.335 ;
        RECT  4.990 -0.115 5.110 0.115 ;
        RECT  4.910 -0.115 4.990 0.335 ;
        RECT  4.800 -0.115 4.910 0.115 ;
        RECT  4.720 -0.115 4.800 0.335 ;
        RECT  4.610 -0.115 4.720 0.115 ;
        RECT  4.530 -0.115 4.610 0.335 ;
        RECT  4.420 -0.115 4.530 0.115 ;
        RECT  4.340 -0.115 4.420 0.335 ;
        RECT  4.210 -0.115 4.340 0.115 ;
        RECT  4.130 -0.115 4.210 0.335 ;
        RECT  4.000 -0.115 4.130 0.115 ;
        RECT  3.920 -0.115 4.000 0.335 ;
        RECT  3.790 -0.115 3.920 0.115 ;
        RECT  3.710 -0.115 3.790 0.335 ;
        RECT  3.580 -0.115 3.710 0.115 ;
        RECT  3.500 -0.115 3.580 0.335 ;
        RECT  3.370 -0.115 3.500 0.115 ;
        RECT  3.290 -0.115 3.370 0.335 ;
        RECT  3.160 -0.115 3.290 0.115 ;
        RECT  3.080 -0.115 3.160 0.335 ;
        RECT  2.950 -0.115 3.080 0.115 ;
        RECT  2.870 -0.115 2.950 0.335 ;
        RECT  2.750 -0.115 2.870 0.115 ;
        RECT  2.670 -0.115 2.750 0.335 ;
        RECT  2.560 -0.115 2.670 0.115 ;
        RECT  2.480 -0.115 2.560 0.335 ;
        RECT  2.370 -0.115 2.480 0.115 ;
        RECT  2.290 -0.115 2.370 0.335 ;
        RECT  2.175 -0.115 2.290 0.115 ;
        RECT  2.095 -0.115 2.175 0.335 ;
        RECT  1.970 -0.115 2.095 0.115 ;
        RECT  1.890 -0.115 1.970 0.335 ;
        RECT  1.760 -0.115 1.890 0.115 ;
        RECT  1.680 -0.115 1.760 0.335 ;
        RECT  1.550 -0.115 1.680 0.115 ;
        RECT  1.470 -0.115 1.550 0.335 ;
        RECT  1.340 -0.115 1.470 0.115 ;
        RECT  1.260 -0.115 1.340 0.335 ;
        RECT  1.130 -0.115 1.260 0.115 ;
        RECT  1.050 -0.115 1.130 0.335 ;
        RECT  0.920 -0.115 1.050 0.115 ;
        RECT  0.840 -0.115 0.920 0.335 ;
        RECT  0.710 -0.115 0.840 0.115 ;
        RECT  0.630 -0.115 0.710 0.335 ;
        RECT  0.510 -0.115 0.630 0.115 ;
        RECT  0.430 -0.115 0.510 0.335 ;
        RECT  0.320 -0.115 0.430 0.115 ;
        RECT  0.240 -0.115 0.320 0.335 ;
        RECT  0.130 -0.115 0.240 0.115 ;
        RECT  0.050 -0.115 0.130 0.335 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.690 1.145 8.960 1.375 ;
        RECT  8.610 0.945 8.690 1.375 ;
        RECT  8.480 1.145 8.610 1.375 ;
        RECT  8.400 0.945 8.480 1.375 ;
        RECT  8.270 1.145 8.400 1.375 ;
        RECT  8.190 0.795 8.270 1.375 ;
        RECT  8.060 1.145 8.190 1.375 ;
        RECT  7.980 0.795 8.060 1.375 ;
        RECT  7.850 1.145 7.980 1.375 ;
        RECT  7.770 0.795 7.850 1.375 ;
        RECT  7.640 1.145 7.770 1.375 ;
        RECT  7.560 0.795 7.640 1.375 ;
        RECT  7.430 1.145 7.560 1.375 ;
        RECT  7.350 0.795 7.430 1.375 ;
        RECT  7.230 1.145 7.350 1.375 ;
        RECT  7.150 0.795 7.230 1.375 ;
        RECT  7.040 1.145 7.150 1.375 ;
        RECT  6.960 0.795 7.040 1.375 ;
        RECT  6.850 1.145 6.960 1.375 ;
        RECT  6.770 0.795 6.850 1.375 ;
        RECT  6.655 1.145 6.770 1.375 ;
        RECT  6.575 0.795 6.655 1.375 ;
        RECT  6.450 1.145 6.575 1.375 ;
        RECT  6.370 0.795 6.450 1.375 ;
        RECT  6.240 1.145 6.370 1.375 ;
        RECT  6.160 0.795 6.240 1.375 ;
        RECT  6.030 1.145 6.160 1.375 ;
        RECT  5.950 0.795 6.030 1.375 ;
        RECT  5.820 1.145 5.950 1.375 ;
        RECT  5.740 0.795 5.820 1.375 ;
        RECT  5.610 1.145 5.740 1.375 ;
        RECT  5.530 0.795 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.795 5.400 1.375 ;
        RECT  5.190 1.145 5.320 1.375 ;
        RECT  5.110 0.795 5.190 1.375 ;
        RECT  4.990 1.145 5.110 1.375 ;
        RECT  4.910 0.795 4.990 1.375 ;
        RECT  4.800 1.145 4.910 1.375 ;
        RECT  4.720 0.795 4.800 1.375 ;
        RECT  4.610 1.145 4.720 1.375 ;
        RECT  4.530 0.795 4.610 1.375 ;
        RECT  4.415 1.145 4.530 1.375 ;
        RECT  4.335 0.795 4.415 1.375 ;
        RECT  4.210 1.145 4.335 1.375 ;
        RECT  4.130 0.795 4.210 1.375 ;
        RECT  4.000 1.145 4.130 1.375 ;
        RECT  3.920 0.795 4.000 1.375 ;
        RECT  3.790 1.145 3.920 1.375 ;
        RECT  3.710 0.795 3.790 1.375 ;
        RECT  3.580 1.145 3.710 1.375 ;
        RECT  3.500 0.795 3.580 1.375 ;
        RECT  3.370 1.145 3.500 1.375 ;
        RECT  3.290 0.795 3.370 1.375 ;
        RECT  3.160 1.145 3.290 1.375 ;
        RECT  3.080 0.795 3.160 1.375 ;
        RECT  2.950 1.145 3.080 1.375 ;
        RECT  2.870 0.795 2.950 1.375 ;
        RECT  2.750 1.145 2.870 1.375 ;
        RECT  2.670 0.795 2.750 1.375 ;
        RECT  2.560 1.145 2.670 1.375 ;
        RECT  2.480 0.795 2.560 1.375 ;
        RECT  2.370 1.145 2.480 1.375 ;
        RECT  2.290 0.795 2.370 1.375 ;
        RECT  2.175 1.145 2.290 1.375 ;
        RECT  2.095 0.795 2.175 1.375 ;
        RECT  1.970 1.145 2.095 1.375 ;
        RECT  1.890 0.795 1.970 1.375 ;
        RECT  1.760 1.145 1.890 1.375 ;
        RECT  1.680 0.795 1.760 1.375 ;
        RECT  1.550 1.145 1.680 1.375 ;
        RECT  1.470 0.795 1.550 1.375 ;
        RECT  1.340 1.145 1.470 1.375 ;
        RECT  1.260 0.795 1.340 1.375 ;
        RECT  1.130 1.145 1.260 1.375 ;
        RECT  1.050 0.795 1.130 1.375 ;
        RECT  0.920 1.145 1.050 1.375 ;
        RECT  0.840 0.795 0.920 1.375 ;
        RECT  0.710 1.145 0.840 1.375 ;
        RECT  0.630 0.795 0.710 1.375 ;
        RECT  0.510 1.145 0.630 1.375 ;
        RECT  0.430 0.795 0.510 1.375 ;
        RECT  0.320 1.145 0.430 1.375 ;
        RECT  0.240 0.795 0.320 1.375 ;
        RECT  0.130 1.145 0.240 1.375 ;
        RECT  0.050 0.795 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.830 0.210 8.910 0.710 ;
        RECT  8.830 0.790 8.910 1.060 ;
        RECT  8.570 0.630 8.830 0.710 ;
        RECT  8.500 0.790 8.830 0.870 ;
        RECT  8.420 0.430 8.500 0.870 ;
        RECT  0.205 0.430 8.420 0.510 ;
    END
END DCAP64BWP40

MACRO DCAP8BWP40
    CLASS CORE ;
    FOREIGN DCAP8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.835 -0.115 1.120 0.115 ;
        RECT  0.755 -0.115 0.835 0.330 ;
        RECT  0.600 -0.115 0.755 0.115 ;
        RECT  0.520 -0.115 0.600 0.330 ;
        RECT  0.365 -0.115 0.520 0.115 ;
        RECT  0.285 -0.115 0.365 0.330 ;
        RECT  0.150 -0.115 0.285 0.115 ;
        RECT  0.070 -0.115 0.150 0.330 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.145 1.120 1.375 ;
        RECT  0.750 0.955 0.830 1.375 ;
        RECT  0.595 1.145 0.750 1.375 ;
        RECT  0.515 0.955 0.595 1.375 ;
        RECT  0.370 1.145 0.515 1.375 ;
        RECT  0.290 0.805 0.370 1.375 ;
        RECT  0.150 1.145 0.290 1.375 ;
        RECT  0.070 0.805 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.975 0.210 1.055 0.710 ;
        RECT  0.975 0.790 1.055 1.050 ;
        RECT  0.740 0.630 0.975 0.710 ;
        RECT  0.670 0.790 0.975 0.870 ;
        RECT  0.590 0.430 0.670 0.870 ;
        RECT  0.280 0.430 0.590 0.510 ;
    END
END DCAP8BWP40

MACRO DCCKBD10BWP40
    CLASS CORE ;
    FOREIGN DCCKBD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.600000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  1.995 0.305 2.195 0.465 ;
        RECT  1.885 0.305 1.995 0.950 ;
        RECT  1.815 0.185 1.885 0.950 ;
        RECT  1.785 0.305 1.815 0.950 ;
        RECT  1.505 0.305 1.785 0.465 ;
        RECT  1.030 0.720 1.785 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.610 -0.115 5.880 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.170 -0.115 5.320 0.115 ;
        RECT  5.090 -0.115 5.170 0.335 ;
        RECT  4.935 -0.115 5.090 0.115 ;
        RECT  4.855 -0.115 4.935 0.335 ;
        RECT  4.700 -0.115 4.855 0.115 ;
        RECT  4.620 -0.115 4.700 0.335 ;
        RECT  4.490 -0.115 4.620 0.115 ;
        RECT  4.410 -0.115 4.490 0.335 ;
        RECT  4.280 -0.115 4.410 0.115 ;
        RECT  4.200 -0.115 4.280 0.335 ;
        RECT  4.070 -0.115 4.200 0.115 ;
        RECT  3.990 -0.115 4.070 0.335 ;
        RECT  3.860 -0.115 3.990 0.115 ;
        RECT  3.780 -0.115 3.860 0.335 ;
        RECT  3.650 -0.115 3.780 0.115 ;
        RECT  3.570 -0.115 3.650 0.335 ;
        RECT  3.450 -0.115 3.570 0.115 ;
        RECT  3.370 -0.115 3.450 0.335 ;
        RECT  3.260 -0.115 3.370 0.115 ;
        RECT  3.180 -0.115 3.260 0.335 ;
        RECT  3.070 -0.115 3.180 0.115 ;
        RECT  2.990 -0.115 3.070 0.335 ;
        RECT  2.840 -0.115 2.990 0.115 ;
        RECT  2.760 -0.115 2.840 0.465 ;
        RECT  2.480 -0.115 2.760 0.115 ;
        RECT  2.360 -0.115 2.480 0.235 ;
        RECT  2.100 -0.115 2.360 0.115 ;
        RECT  1.980 -0.115 2.100 0.235 ;
        RECT  1.720 -0.115 1.980 0.115 ;
        RECT  1.600 -0.115 1.720 0.235 ;
        RECT  1.340 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.340 0.235 ;
        RECT  0.940 -0.115 1.220 0.115 ;
        RECT  0.860 -0.115 0.940 0.465 ;
        RECT  0.565 -0.115 0.860 0.115 ;
        RECT  0.475 -0.115 0.565 0.260 ;
        RECT  0.190 -0.115 0.475 0.115 ;
        RECT  0.090 -0.115 0.190 0.410 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.610 1.145 5.880 1.375 ;
        RECT  5.530 0.945 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.945 5.400 1.375 ;
        RECT  5.170 1.145 5.320 1.375 ;
        RECT  5.090 0.795 5.170 1.375 ;
        RECT  4.935 1.145 5.090 1.375 ;
        RECT  4.855 0.795 4.935 1.375 ;
        RECT  4.700 1.145 4.855 1.375 ;
        RECT  4.620 0.795 4.700 1.375 ;
        RECT  4.490 1.145 4.620 1.375 ;
        RECT  4.410 0.795 4.490 1.375 ;
        RECT  4.280 1.145 4.410 1.375 ;
        RECT  4.200 0.795 4.280 1.375 ;
        RECT  4.070 1.145 4.200 1.375 ;
        RECT  3.990 0.795 4.070 1.375 ;
        RECT  3.860 1.145 3.990 1.375 ;
        RECT  3.780 0.795 3.860 1.375 ;
        RECT  3.650 1.145 3.780 1.375 ;
        RECT  3.570 0.795 3.650 1.375 ;
        RECT  3.450 1.145 3.570 1.375 ;
        RECT  3.370 0.795 3.450 1.375 ;
        RECT  3.260 1.145 3.370 1.375 ;
        RECT  3.180 0.795 3.260 1.375 ;
        RECT  3.070 1.145 3.180 1.375 ;
        RECT  2.990 0.795 3.070 1.375 ;
        RECT  2.840 1.145 2.990 1.375 ;
        RECT  2.760 0.700 2.840 1.375 ;
        RECT  2.480 1.145 2.760 1.375 ;
        RECT  2.360 1.020 2.480 1.375 ;
        RECT  2.100 1.145 2.360 1.375 ;
        RECT  1.980 1.020 2.100 1.375 ;
        RECT  1.720 1.145 1.980 1.375 ;
        RECT  1.600 1.020 1.720 1.375 ;
        RECT  1.340 1.145 1.600 1.375 ;
        RECT  1.220 1.020 1.340 1.375 ;
        RECT  0.940 1.145 1.220 1.375 ;
        RECT  0.860 0.720 0.940 1.375 ;
        RECT  0.560 1.145 0.860 1.375 ;
        RECT  0.480 0.995 0.560 1.375 ;
        RECT  0.190 1.145 0.480 1.375 ;
        RECT  0.090 0.845 0.190 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.065 0.720 2.670 0.950 ;
        RECT  2.575 0.185 2.645 0.465 ;
        RECT  2.265 0.305 2.575 0.465 ;
        RECT  2.195 0.185 2.265 0.465 ;
        RECT  2.065 0.305 2.195 0.465 ;
        RECT  1.505 0.305 1.715 0.465 ;
        RECT  1.030 0.720 1.715 0.950 ;
        RECT  1.435 0.185 1.505 0.465 ;
        RECT  1.125 0.305 1.435 0.465 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  5.750 0.210 5.830 0.710 ;
        RECT  5.750 0.790 5.830 1.060 ;
        RECT  5.490 0.630 5.750 0.710 ;
        RECT  5.420 0.790 5.750 0.870 ;
        RECT  5.340 0.430 5.420 0.870 ;
        RECT  3.145 0.430 5.340 0.510 ;
        RECT  0.770 0.545 1.705 0.615 ;
        RECT  0.660 0.195 0.770 1.050 ;
        RECT  0.390 0.335 0.660 0.415 ;
        RECT  0.365 0.770 0.660 0.850 ;
        RECT  0.270 0.205 0.390 0.415 ;
        RECT  0.295 0.770 0.365 1.050 ;
    END
END DCCKBD10BWP40

MACRO DCCKBD12BWP40
    CLASS CORE ;
    FOREIGN DCCKBD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.275 0.305 2.525 0.465 ;
        RECT  2.215 0.305 2.275 0.950 ;
        RECT  2.135 0.185 2.215 0.950 ;
        RECT  1.925 0.305 2.135 0.950 ;
        RECT  1.835 0.305 1.925 0.465 ;
        RECT  0.980 0.720 1.925 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.123200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.170 -0.115 6.440 0.115 ;
        RECT  6.090 -0.115 6.170 0.335 ;
        RECT  5.960 -0.115 6.090 0.115 ;
        RECT  5.880 -0.115 5.960 0.335 ;
        RECT  5.760 -0.115 5.880 0.115 ;
        RECT  5.680 -0.115 5.760 0.335 ;
        RECT  5.570 -0.115 5.680 0.115 ;
        RECT  5.490 -0.115 5.570 0.335 ;
        RECT  5.375 -0.115 5.490 0.115 ;
        RECT  5.295 -0.115 5.375 0.335 ;
        RECT  5.180 -0.115 5.295 0.115 ;
        RECT  5.100 -0.115 5.180 0.335 ;
        RECT  4.980 -0.115 5.100 0.115 ;
        RECT  4.900 -0.115 4.980 0.335 ;
        RECT  4.770 -0.115 4.900 0.115 ;
        RECT  4.690 -0.115 4.770 0.335 ;
        RECT  4.560 -0.115 4.690 0.115 ;
        RECT  4.480 -0.115 4.560 0.335 ;
        RECT  4.350 -0.115 4.480 0.115 ;
        RECT  4.270 -0.115 4.350 0.335 ;
        RECT  4.140 -0.115 4.270 0.115 ;
        RECT  4.060 -0.115 4.140 0.335 ;
        RECT  3.930 -0.115 4.060 0.115 ;
        RECT  3.850 -0.115 3.930 0.335 ;
        RECT  3.730 -0.115 3.850 0.115 ;
        RECT  3.650 -0.115 3.730 0.335 ;
        RECT  3.540 -0.115 3.650 0.115 ;
        RECT  3.460 -0.115 3.540 0.335 ;
        RECT  3.350 -0.115 3.460 0.115 ;
        RECT  3.270 -0.115 3.350 0.335 ;
        RECT  3.170 -0.115 3.270 0.115 ;
        RECT  3.090 -0.115 3.170 0.465 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.235 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.235 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.890 -0.115 1.170 0.115 ;
        RECT  0.810 -0.115 0.890 0.465 ;
        RECT  0.515 -0.115 0.810 0.115 ;
        RECT  0.425 -0.115 0.515 0.260 ;
        RECT  0.140 -0.115 0.425 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.145 6.440 1.375 ;
        RECT  6.090 0.945 6.170 1.375 ;
        RECT  5.960 1.145 6.090 1.375 ;
        RECT  5.880 0.945 5.960 1.375 ;
        RECT  5.760 1.145 5.880 1.375 ;
        RECT  5.680 0.795 5.760 1.375 ;
        RECT  5.570 1.145 5.680 1.375 ;
        RECT  5.490 0.795 5.570 1.375 ;
        RECT  5.375 1.145 5.490 1.375 ;
        RECT  5.295 0.795 5.375 1.375 ;
        RECT  5.180 1.145 5.295 1.375 ;
        RECT  5.100 0.795 5.180 1.375 ;
        RECT  4.980 1.145 5.100 1.375 ;
        RECT  4.900 0.795 4.980 1.375 ;
        RECT  4.770 1.145 4.900 1.375 ;
        RECT  4.690 0.795 4.770 1.375 ;
        RECT  4.560 1.145 4.690 1.375 ;
        RECT  4.480 0.795 4.560 1.375 ;
        RECT  4.350 1.145 4.480 1.375 ;
        RECT  4.270 0.795 4.350 1.375 ;
        RECT  4.140 1.145 4.270 1.375 ;
        RECT  4.060 0.795 4.140 1.375 ;
        RECT  3.930 1.145 4.060 1.375 ;
        RECT  3.850 0.795 3.930 1.375 ;
        RECT  3.730 1.145 3.850 1.375 ;
        RECT  3.650 0.795 3.730 1.375 ;
        RECT  3.540 1.145 3.650 1.375 ;
        RECT  3.460 0.795 3.540 1.375 ;
        RECT  3.350 1.145 3.460 1.375 ;
        RECT  3.270 0.795 3.350 1.375 ;
        RECT  3.170 1.145 3.270 1.375 ;
        RECT  3.090 0.700 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 1.020 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 1.020 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 1.020 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.020 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 1.020 1.290 1.375 ;
        RECT  0.890 1.145 1.170 1.375 ;
        RECT  0.810 0.720 0.890 1.375 ;
        RECT  0.530 1.145 0.810 1.375 ;
        RECT  0.410 0.910 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.720 3.000 0.950 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.595 0.305 2.905 0.465 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.345 0.305 2.525 0.465 ;
        RECT  1.835 0.305 1.855 0.465 ;
        RECT  0.980 0.720 1.855 0.950 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.455 0.305 1.765 0.465 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.305 1.385 0.465 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  6.310 0.210 6.390 0.710 ;
        RECT  6.310 0.790 6.390 1.060 ;
        RECT  6.050 0.630 6.310 0.710 ;
        RECT  5.980 0.790 6.310 0.870 ;
        RECT  5.900 0.430 5.980 0.870 ;
        RECT  3.425 0.430 5.900 0.510 ;
        RECT  0.720 0.545 1.765 0.615 ;
        RECT  0.610 0.195 0.720 1.050 ;
        RECT  0.340 0.335 0.610 0.415 ;
        RECT  0.315 0.750 0.610 0.830 ;
        RECT  0.220 0.205 0.340 0.415 ;
        RECT  0.245 0.750 0.315 1.050 ;
    END
END DCCKBD12BWP40

MACRO DCCKBD14BWP40
    CLASS CORE ;
    FOREIGN DCCKBD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.872000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.835 0.305 3.125 0.465 ;
        RECT  2.815 0.305 2.835 0.945 ;
        RECT  2.745 0.185 2.815 0.945 ;
        RECT  2.485 0.305 2.745 0.945 ;
        RECT  2.435 0.305 2.485 0.465 ;
        RECT  1.200 0.715 2.485 0.945 ;
        RECT  2.365 0.185 2.435 0.465 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.156000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.665 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.570 -0.115 7.840 0.115 ;
        RECT  7.490 -0.115 7.570 0.335 ;
        RECT  7.360 -0.115 7.490 0.115 ;
        RECT  7.280 -0.115 7.360 0.335 ;
        RECT  7.150 -0.115 7.280 0.115 ;
        RECT  7.070 -0.115 7.150 0.335 ;
        RECT  6.940 -0.115 7.070 0.115 ;
        RECT  6.860 -0.115 6.940 0.335 ;
        RECT  6.705 -0.115 6.860 0.115 ;
        RECT  6.625 -0.115 6.705 0.335 ;
        RECT  6.480 -0.115 6.625 0.115 ;
        RECT  6.400 -0.115 6.480 0.335 ;
        RECT  6.290 -0.115 6.400 0.115 ;
        RECT  6.210 -0.115 6.290 0.335 ;
        RECT  6.095 -0.115 6.210 0.115 ;
        RECT  6.015 -0.115 6.095 0.335 ;
        RECT  5.890 -0.115 6.015 0.115 ;
        RECT  5.810 -0.115 5.890 0.335 ;
        RECT  5.680 -0.115 5.810 0.115 ;
        RECT  5.600 -0.115 5.680 0.335 ;
        RECT  5.470 -0.115 5.600 0.115 ;
        RECT  5.390 -0.115 5.470 0.335 ;
        RECT  5.260 -0.115 5.390 0.115 ;
        RECT  5.180 -0.115 5.260 0.335 ;
        RECT  5.050 -0.115 5.180 0.115 ;
        RECT  4.970 -0.115 5.050 0.335 ;
        RECT  4.840 -0.115 4.970 0.115 ;
        RECT  4.760 -0.115 4.840 0.335 ;
        RECT  4.630 -0.115 4.760 0.115 ;
        RECT  4.550 -0.115 4.630 0.335 ;
        RECT  4.430 -0.115 4.550 0.115 ;
        RECT  4.350 -0.115 4.430 0.335 ;
        RECT  4.240 -0.115 4.350 0.115 ;
        RECT  4.160 -0.115 4.240 0.335 ;
        RECT  4.050 -0.115 4.160 0.115 ;
        RECT  3.970 -0.115 4.050 0.335 ;
        RECT  3.835 -0.115 3.970 0.115 ;
        RECT  3.730 -0.115 3.835 0.465 ;
        RECT  3.410 -0.115 3.730 0.115 ;
        RECT  3.290 -0.115 3.410 0.235 ;
        RECT  3.030 -0.115 3.290 0.115 ;
        RECT  2.910 -0.115 3.030 0.235 ;
        RECT  2.650 -0.115 2.910 0.115 ;
        RECT  2.530 -0.115 2.650 0.235 ;
        RECT  2.270 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.270 0.235 ;
        RECT  1.890 -0.115 2.150 0.115 ;
        RECT  1.770 -0.115 1.890 0.235 ;
        RECT  1.510 -0.115 1.770 0.115 ;
        RECT  1.390 -0.115 1.510 0.235 ;
        RECT  1.100 -0.115 1.390 0.115 ;
        RECT  1.020 -0.115 1.100 0.465 ;
        RECT  0.720 -0.115 1.020 0.115 ;
        RECT  0.600 -0.115 0.720 0.265 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.570 1.145 7.840 1.375 ;
        RECT  7.490 0.945 7.570 1.375 ;
        RECT  7.360 1.145 7.490 1.375 ;
        RECT  7.280 0.945 7.360 1.375 ;
        RECT  7.150 1.145 7.280 1.375 ;
        RECT  7.070 0.795 7.150 1.375 ;
        RECT  6.940 1.145 7.070 1.375 ;
        RECT  6.860 0.795 6.940 1.375 ;
        RECT  6.705 1.145 6.860 1.375 ;
        RECT  6.625 0.795 6.705 1.375 ;
        RECT  6.480 1.145 6.625 1.375 ;
        RECT  6.400 0.795 6.480 1.375 ;
        RECT  6.290 1.145 6.400 1.375 ;
        RECT  6.210 0.795 6.290 1.375 ;
        RECT  6.095 1.145 6.210 1.375 ;
        RECT  6.015 0.795 6.095 1.375 ;
        RECT  5.890 1.145 6.015 1.375 ;
        RECT  5.810 0.795 5.890 1.375 ;
        RECT  5.680 1.145 5.810 1.375 ;
        RECT  5.600 0.795 5.680 1.375 ;
        RECT  5.470 1.145 5.600 1.375 ;
        RECT  5.390 0.795 5.470 1.375 ;
        RECT  5.260 1.145 5.390 1.375 ;
        RECT  5.180 0.795 5.260 1.375 ;
        RECT  5.050 1.145 5.180 1.375 ;
        RECT  4.970 0.795 5.050 1.375 ;
        RECT  4.840 1.145 4.970 1.375 ;
        RECT  4.760 0.795 4.840 1.375 ;
        RECT  4.630 1.145 4.760 1.375 ;
        RECT  4.550 0.795 4.630 1.375 ;
        RECT  4.430 1.145 4.550 1.375 ;
        RECT  4.350 0.795 4.430 1.375 ;
        RECT  4.240 1.145 4.350 1.375 ;
        RECT  4.160 0.795 4.240 1.375 ;
        RECT  4.050 1.145 4.160 1.375 ;
        RECT  3.970 0.795 4.050 1.375 ;
        RECT  3.835 1.145 3.970 1.375 ;
        RECT  3.730 0.690 3.835 1.375 ;
        RECT  3.410 1.145 3.730 1.375 ;
        RECT  3.290 1.015 3.410 1.375 ;
        RECT  3.030 1.145 3.290 1.375 ;
        RECT  2.910 1.015 3.030 1.375 ;
        RECT  2.650 1.145 2.910 1.375 ;
        RECT  2.530 1.015 2.650 1.375 ;
        RECT  2.270 1.145 2.530 1.375 ;
        RECT  2.150 1.015 2.270 1.375 ;
        RECT  1.890 1.145 2.150 1.375 ;
        RECT  1.770 1.015 1.890 1.375 ;
        RECT  1.510 1.145 1.770 1.375 ;
        RECT  1.390 1.015 1.510 1.375 ;
        RECT  1.120 1.145 1.390 1.375 ;
        RECT  1.000 0.710 1.120 1.375 ;
        RECT  0.700 1.145 1.000 1.375 ;
        RECT  0.620 1.000 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 1.000 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.675 0.305 1.985 0.465 ;
        RECT  1.605 0.185 1.675 0.465 ;
        RECT  1.295 0.305 1.605 0.465 ;
        RECT  1.225 0.185 1.295 0.465 ;
        RECT  7.710 0.210 7.790 0.710 ;
        RECT  7.710 0.790 7.790 1.060 ;
        RECT  7.450 0.630 7.710 0.710 ;
        RECT  7.380 0.790 7.710 0.870 ;
        RECT  7.300 0.430 7.380 0.870 ;
        RECT  4.125 0.430 7.300 0.510 ;
        RECT  0.920 0.545 2.405 0.615 ;
        RECT  0.790 0.195 0.920 1.065 ;
        RECT  0.510 0.335 0.790 0.415 ;
        RECT  0.525 0.845 0.790 0.915 ;
        RECT  0.415 0.845 0.525 1.075 ;
        RECT  0.430 0.185 0.510 0.415 ;
        RECT  0.130 0.335 0.430 0.415 ;
        RECT  0.125 0.845 0.415 0.915 ;
        RECT  0.055 0.255 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.075 ;
        RECT  2.905 0.715 3.640 0.945 ;
        RECT  3.505 0.185 3.575 0.465 ;
        RECT  3.195 0.305 3.505 0.465 ;
        RECT  3.125 0.185 3.195 0.465 ;
        RECT  2.905 0.305 3.125 0.465 ;
        RECT  2.365 0.185 2.415 0.465 ;
        RECT  1.200 0.715 2.415 0.945 ;
        RECT  2.055 0.305 2.365 0.465 ;
        RECT  1.985 0.185 2.055 0.465 ;
    END
END DCCKBD14BWP40

MACRO DCCKBD16BWP40
    CLASS CORE ;
    FOREIGN DCCKBD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.115 0.305 3.405 0.465 ;
        RECT  3.095 0.305 3.115 0.945 ;
        RECT  3.025 0.185 3.095 0.945 ;
        RECT  2.765 0.305 3.025 0.945 ;
        RECT  2.715 0.305 2.765 0.465 ;
        RECT  1.480 0.715 2.765 0.945 ;
        RECT  2.645 0.185 2.715 0.465 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.184800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.945 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.690 -0.115 8.960 0.115 ;
        RECT  8.610 -0.115 8.690 0.335 ;
        RECT  8.480 -0.115 8.610 0.115 ;
        RECT  8.400 -0.115 8.480 0.335 ;
        RECT  8.270 -0.115 8.400 0.115 ;
        RECT  8.190 -0.115 8.270 0.335 ;
        RECT  8.060 -0.115 8.190 0.115 ;
        RECT  7.980 -0.115 8.060 0.335 ;
        RECT  7.850 -0.115 7.980 0.115 ;
        RECT  7.770 -0.115 7.850 0.335 ;
        RECT  7.640 -0.115 7.770 0.115 ;
        RECT  7.560 -0.115 7.640 0.335 ;
        RECT  7.430 -0.115 7.560 0.115 ;
        RECT  7.350 -0.115 7.430 0.335 ;
        RECT  7.230 -0.115 7.350 0.115 ;
        RECT  7.150 -0.115 7.230 0.335 ;
        RECT  7.040 -0.115 7.150 0.115 ;
        RECT  6.960 -0.115 7.040 0.335 ;
        RECT  6.850 -0.115 6.960 0.115 ;
        RECT  6.770 -0.115 6.850 0.335 ;
        RECT  6.655 -0.115 6.770 0.115 ;
        RECT  6.575 -0.115 6.655 0.335 ;
        RECT  6.450 -0.115 6.575 0.115 ;
        RECT  6.370 -0.115 6.450 0.335 ;
        RECT  6.240 -0.115 6.370 0.115 ;
        RECT  6.160 -0.115 6.240 0.335 ;
        RECT  6.030 -0.115 6.160 0.115 ;
        RECT  5.950 -0.115 6.030 0.335 ;
        RECT  5.820 -0.115 5.950 0.115 ;
        RECT  5.740 -0.115 5.820 0.335 ;
        RECT  5.610 -0.115 5.740 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.190 -0.115 5.320 0.115 ;
        RECT  5.110 -0.115 5.190 0.335 ;
        RECT  4.990 -0.115 5.110 0.115 ;
        RECT  4.910 -0.115 4.990 0.335 ;
        RECT  4.800 -0.115 4.910 0.115 ;
        RECT  4.720 -0.115 4.800 0.335 ;
        RECT  4.610 -0.115 4.720 0.115 ;
        RECT  4.530 -0.115 4.610 0.335 ;
        RECT  4.430 -0.115 4.530 0.115 ;
        RECT  4.350 -0.115 4.430 0.465 ;
        RECT  4.070 -0.115 4.350 0.115 ;
        RECT  3.950 -0.115 4.070 0.235 ;
        RECT  3.690 -0.115 3.950 0.115 ;
        RECT  3.570 -0.115 3.690 0.235 ;
        RECT  3.310 -0.115 3.570 0.115 ;
        RECT  3.190 -0.115 3.310 0.235 ;
        RECT  2.930 -0.115 3.190 0.115 ;
        RECT  2.810 -0.115 2.930 0.235 ;
        RECT  2.550 -0.115 2.810 0.115 ;
        RECT  2.430 -0.115 2.550 0.235 ;
        RECT  2.170 -0.115 2.430 0.115 ;
        RECT  2.050 -0.115 2.170 0.235 ;
        RECT  1.790 -0.115 2.050 0.115 ;
        RECT  1.670 -0.115 1.790 0.235 ;
        RECT  1.380 -0.115 1.670 0.115 ;
        RECT  1.300 -0.115 1.380 0.465 ;
        RECT  1.000 -0.115 1.300 0.115 ;
        RECT  0.880 -0.115 1.000 0.265 ;
        RECT  0.620 -0.115 0.880 0.115 ;
        RECT  0.500 -0.115 0.620 0.265 ;
        RECT  0.180 -0.115 0.500 0.115 ;
        RECT  0.060 -0.115 0.180 0.415 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.690 1.145 8.960 1.375 ;
        RECT  8.610 0.945 8.690 1.375 ;
        RECT  8.480 1.145 8.610 1.375 ;
        RECT  8.400 0.945 8.480 1.375 ;
        RECT  8.270 1.145 8.400 1.375 ;
        RECT  8.190 0.795 8.270 1.375 ;
        RECT  8.060 1.145 8.190 1.375 ;
        RECT  7.980 0.795 8.060 1.375 ;
        RECT  7.850 1.145 7.980 1.375 ;
        RECT  7.770 0.795 7.850 1.375 ;
        RECT  7.640 1.145 7.770 1.375 ;
        RECT  7.560 0.795 7.640 1.375 ;
        RECT  7.430 1.145 7.560 1.375 ;
        RECT  7.350 0.795 7.430 1.375 ;
        RECT  7.230 1.145 7.350 1.375 ;
        RECT  7.150 0.795 7.230 1.375 ;
        RECT  7.040 1.145 7.150 1.375 ;
        RECT  6.960 0.795 7.040 1.375 ;
        RECT  6.850 1.145 6.960 1.375 ;
        RECT  6.770 0.795 6.850 1.375 ;
        RECT  6.655 1.145 6.770 1.375 ;
        RECT  6.575 0.795 6.655 1.375 ;
        RECT  6.450 1.145 6.575 1.375 ;
        RECT  6.370 0.795 6.450 1.375 ;
        RECT  6.240 1.145 6.370 1.375 ;
        RECT  6.160 0.795 6.240 1.375 ;
        RECT  6.030 1.145 6.160 1.375 ;
        RECT  5.950 0.795 6.030 1.375 ;
        RECT  5.820 1.145 5.950 1.375 ;
        RECT  5.740 0.795 5.820 1.375 ;
        RECT  5.610 1.145 5.740 1.375 ;
        RECT  5.530 0.795 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.795 5.400 1.375 ;
        RECT  5.190 1.145 5.320 1.375 ;
        RECT  5.110 0.795 5.190 1.375 ;
        RECT  4.990 1.145 5.110 1.375 ;
        RECT  4.910 0.795 4.990 1.375 ;
        RECT  4.800 1.145 4.910 1.375 ;
        RECT  4.720 0.795 4.800 1.375 ;
        RECT  4.610 1.145 4.720 1.375 ;
        RECT  4.530 0.795 4.610 1.375 ;
        RECT  4.430 1.145 4.530 1.375 ;
        RECT  4.350 0.690 4.430 1.375 ;
        RECT  4.070 1.145 4.350 1.375 ;
        RECT  3.950 1.015 4.070 1.375 ;
        RECT  3.690 1.145 3.950 1.375 ;
        RECT  3.570 1.015 3.690 1.375 ;
        RECT  3.310 1.145 3.570 1.375 ;
        RECT  3.190 1.015 3.310 1.375 ;
        RECT  2.930 1.145 3.190 1.375 ;
        RECT  2.810 1.015 2.930 1.375 ;
        RECT  2.550 1.145 2.810 1.375 ;
        RECT  2.430 1.015 2.550 1.375 ;
        RECT  2.170 1.145 2.430 1.375 ;
        RECT  2.050 1.015 2.170 1.375 ;
        RECT  1.790 1.145 2.050 1.375 ;
        RECT  1.670 1.015 1.790 1.375 ;
        RECT  1.400 1.145 1.670 1.375 ;
        RECT  1.280 0.710 1.400 1.375 ;
        RECT  0.980 1.145 1.280 1.375 ;
        RECT  0.900 0.860 0.980 1.375 ;
        RECT  0.600 1.145 0.900 1.375 ;
        RECT  0.520 0.860 0.600 1.375 ;
        RECT  0.170 1.145 0.520 1.375 ;
        RECT  0.090 0.845 0.170 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.260 0.945 ;
        RECT  4.165 0.185 4.235 0.465 ;
        RECT  3.855 0.305 4.165 0.465 ;
        RECT  3.785 0.185 3.855 0.465 ;
        RECT  3.475 0.305 3.785 0.465 ;
        RECT  3.405 0.185 3.475 0.465 ;
        RECT  3.185 0.305 3.405 0.465 ;
        RECT  2.645 0.185 2.695 0.465 ;
        RECT  1.480 0.715 2.695 0.945 ;
        RECT  4.685 0.430 8.420 0.510 ;
        RECT  1.200 0.545 2.685 0.615 ;
        RECT  1.070 0.195 1.200 1.065 ;
        RECT  0.790 0.335 1.070 0.415 ;
        RECT  0.785 0.705 1.070 0.785 ;
        RECT  0.710 0.185 0.790 0.415 ;
        RECT  0.715 0.705 0.785 1.035 ;
        RECT  0.405 0.705 0.715 0.785 ;
        RECT  0.410 0.335 0.710 0.415 ;
        RECT  0.310 0.185 0.410 0.415 ;
        RECT  0.335 0.705 0.405 1.035 ;
        RECT  2.335 0.305 2.645 0.465 ;
        RECT  2.265 0.185 2.335 0.465 ;
        RECT  1.955 0.305 2.265 0.465 ;
        RECT  1.885 0.185 1.955 0.465 ;
        RECT  1.575 0.305 1.885 0.465 ;
        RECT  1.505 0.185 1.575 0.465 ;
        RECT  8.830 0.210 8.910 0.710 ;
        RECT  8.830 0.790 8.910 1.060 ;
        RECT  8.570 0.630 8.830 0.710 ;
        RECT  8.500 0.790 8.830 0.870 ;
        RECT  8.420 0.430 8.500 0.870 ;
    END
END DCCKBD16BWP40

MACRO DCCKBD18BWP40
    CLASS CORE ;
    FOREIGN DCCKBD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.080000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.105 0.305 3.305 0.465 ;
        RECT  2.995 0.305 3.105 0.945 ;
        RECT  2.925 0.185 2.995 0.945 ;
        RECT  2.765 0.305 2.925 0.945 ;
        RECT  2.615 0.305 2.765 0.465 ;
        RECT  1.380 0.715 2.765 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  1.405 0.185 1.475 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.184800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.855 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.250 -0.115 9.520 0.115 ;
        RECT  9.170 -0.115 9.250 0.335 ;
        RECT  9.040 -0.115 9.170 0.115 ;
        RECT  8.960 -0.115 9.040 0.335 ;
        RECT  8.830 -0.115 8.960 0.115 ;
        RECT  8.750 -0.115 8.830 0.335 ;
        RECT  8.620 -0.115 8.750 0.115 ;
        RECT  8.540 -0.115 8.620 0.335 ;
        RECT  8.375 -0.115 8.540 0.115 ;
        RECT  8.295 -0.115 8.375 0.335 ;
        RECT  8.130 -0.115 8.295 0.115 ;
        RECT  8.050 -0.115 8.130 0.335 ;
        RECT  7.920 -0.115 8.050 0.115 ;
        RECT  7.840 -0.115 7.920 0.335 ;
        RECT  7.710 -0.115 7.840 0.115 ;
        RECT  7.630 -0.115 7.710 0.335 ;
        RECT  7.510 -0.115 7.630 0.115 ;
        RECT  7.430 -0.115 7.510 0.335 ;
        RECT  7.320 -0.115 7.430 0.115 ;
        RECT  7.240 -0.115 7.320 0.335 ;
        RECT  7.130 -0.115 7.240 0.115 ;
        RECT  7.050 -0.115 7.130 0.335 ;
        RECT  6.935 -0.115 7.050 0.115 ;
        RECT  6.855 -0.115 6.935 0.335 ;
        RECT  6.730 -0.115 6.855 0.115 ;
        RECT  6.650 -0.115 6.730 0.335 ;
        RECT  6.520 -0.115 6.650 0.115 ;
        RECT  6.440 -0.115 6.520 0.335 ;
        RECT  6.310 -0.115 6.440 0.115 ;
        RECT  6.230 -0.115 6.310 0.335 ;
        RECT  6.100 -0.115 6.230 0.115 ;
        RECT  6.020 -0.115 6.100 0.335 ;
        RECT  5.890 -0.115 6.020 0.115 ;
        RECT  5.810 -0.115 5.890 0.335 ;
        RECT  5.680 -0.115 5.810 0.115 ;
        RECT  5.600 -0.115 5.680 0.335 ;
        RECT  5.470 -0.115 5.600 0.115 ;
        RECT  5.390 -0.115 5.470 0.335 ;
        RECT  5.270 -0.115 5.390 0.115 ;
        RECT  5.190 -0.115 5.270 0.335 ;
        RECT  5.080 -0.115 5.190 0.115 ;
        RECT  5.000 -0.115 5.080 0.335 ;
        RECT  4.890 -0.115 5.000 0.115 ;
        RECT  4.810 -0.115 4.890 0.335 ;
        RECT  4.710 -0.115 4.810 0.115 ;
        RECT  4.630 -0.115 4.710 0.465 ;
        RECT  4.350 -0.115 4.630 0.115 ;
        RECT  4.230 -0.115 4.350 0.235 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.235 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.235 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.235 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.235 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.235 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.235 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.235 ;
        RECT  1.280 -0.115 1.570 0.115 ;
        RECT  1.200 -0.115 1.280 0.465 ;
        RECT  0.910 -0.115 1.200 0.115 ;
        RECT  0.790 -0.115 0.910 0.265 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.265 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.250 1.145 9.520 1.375 ;
        RECT  9.170 0.945 9.250 1.375 ;
        RECT  9.040 1.145 9.170 1.375 ;
        RECT  8.960 0.945 9.040 1.375 ;
        RECT  8.830 1.145 8.960 1.375 ;
        RECT  8.750 0.795 8.830 1.375 ;
        RECT  8.620 1.145 8.750 1.375 ;
        RECT  8.540 0.795 8.620 1.375 ;
        RECT  8.375 1.145 8.540 1.375 ;
        RECT  8.295 0.795 8.375 1.375 ;
        RECT  8.130 1.145 8.295 1.375 ;
        RECT  8.050 0.795 8.130 1.375 ;
        RECT  7.920 1.145 8.050 1.375 ;
        RECT  7.840 0.795 7.920 1.375 ;
        RECT  7.710 1.145 7.840 1.375 ;
        RECT  7.630 0.795 7.710 1.375 ;
        RECT  7.510 1.145 7.630 1.375 ;
        RECT  7.430 0.795 7.510 1.375 ;
        RECT  7.320 1.145 7.430 1.375 ;
        RECT  7.240 0.795 7.320 1.375 ;
        RECT  7.130 1.145 7.240 1.375 ;
        RECT  7.050 0.795 7.130 1.375 ;
        RECT  6.935 1.145 7.050 1.375 ;
        RECT  6.855 0.795 6.935 1.375 ;
        RECT  6.730 1.145 6.855 1.375 ;
        RECT  6.650 0.795 6.730 1.375 ;
        RECT  6.520 1.145 6.650 1.375 ;
        RECT  6.440 0.795 6.520 1.375 ;
        RECT  6.310 1.145 6.440 1.375 ;
        RECT  6.230 0.795 6.310 1.375 ;
        RECT  6.100 1.145 6.230 1.375 ;
        RECT  6.020 0.795 6.100 1.375 ;
        RECT  5.890 1.145 6.020 1.375 ;
        RECT  5.810 0.795 5.890 1.375 ;
        RECT  5.680 1.145 5.810 1.375 ;
        RECT  5.600 0.795 5.680 1.375 ;
        RECT  5.470 1.145 5.600 1.375 ;
        RECT  5.390 0.795 5.470 1.375 ;
        RECT  5.270 1.145 5.390 1.375 ;
        RECT  5.190 0.795 5.270 1.375 ;
        RECT  5.080 1.145 5.190 1.375 ;
        RECT  5.000 0.795 5.080 1.375 ;
        RECT  4.890 1.145 5.000 1.375 ;
        RECT  4.810 0.795 4.890 1.375 ;
        RECT  4.710 1.145 4.810 1.375 ;
        RECT  4.630 0.690 4.710 1.375 ;
        RECT  4.350 1.145 4.630 1.375 ;
        RECT  4.230 1.015 4.350 1.375 ;
        RECT  3.970 1.145 4.230 1.375 ;
        RECT  3.850 1.015 3.970 1.375 ;
        RECT  3.590 1.145 3.850 1.375 ;
        RECT  3.470 1.015 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.090 1.015 3.210 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 1.015 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.330 1.015 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 1.015 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.570 1.015 1.690 1.375 ;
        RECT  1.300 1.145 1.570 1.375 ;
        RECT  1.180 0.710 1.300 1.375 ;
        RECT  0.890 1.145 1.180 1.375 ;
        RECT  0.810 0.860 0.890 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.860 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.715 4.540 0.945 ;
        RECT  4.435 0.185 4.515 0.465 ;
        RECT  4.135 0.305 4.435 0.465 ;
        RECT  4.065 0.185 4.135 0.465 ;
        RECT  3.755 0.305 4.065 0.465 ;
        RECT  3.685 0.185 3.755 0.465 ;
        RECT  3.375 0.305 3.685 0.465 ;
        RECT  3.305 0.185 3.375 0.465 ;
        RECT  3.185 0.305 3.305 0.465 ;
        RECT  2.615 0.305 2.695 0.465 ;
        RECT  1.380 0.715 2.695 0.945 ;
        RECT  2.545 0.185 2.615 0.465 ;
        RECT  2.235 0.305 2.545 0.465 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  1.855 0.305 2.165 0.465 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.475 0.305 1.785 0.465 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.625 0.705 0.695 1.035 ;
        RECT  0.315 0.705 0.625 0.785 ;
        RECT  0.320 0.335 0.620 0.415 ;
        RECT  0.220 0.185 0.320 0.415 ;
        RECT  0.245 0.705 0.315 1.035 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  9.390 0.210 9.470 0.710 ;
        RECT  9.390 0.790 9.470 1.060 ;
        RECT  9.130 0.630 9.390 0.710 ;
        RECT  9.060 0.790 9.390 0.870 ;
        RECT  8.980 0.430 9.060 0.870 ;
        RECT  4.965 0.430 8.980 0.510 ;
        RECT  1.110 0.545 2.585 0.615 ;
        RECT  0.980 0.195 1.110 1.065 ;
        RECT  0.700 0.335 0.980 0.415 ;
        RECT  0.695 0.705 0.980 0.785 ;
    END
END DCCKBD18BWP40

MACRO DCCKBD20BWP40
    CLASS CORE ;
    FOREIGN DCCKBD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.200000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.555 0.305 3.865 0.465 ;
        RECT  3.535 0.185 3.555 0.465 ;
        RECT  3.485 0.185 3.535 0.960 ;
        RECT  3.185 0.305 3.485 0.960 ;
        RECT  3.175 0.305 3.185 0.465 ;
        RECT  1.560 0.730 3.185 0.960 ;
        RECT  3.105 0.185 3.175 0.465 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.224000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.065 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.370 -0.115 10.640 0.115 ;
        RECT  10.290 -0.115 10.370 0.335 ;
        RECT  10.160 -0.115 10.290 0.115 ;
        RECT  10.080 -0.115 10.160 0.335 ;
        RECT  9.950 -0.115 10.080 0.115 ;
        RECT  9.870 -0.115 9.950 0.335 ;
        RECT  9.740 -0.115 9.870 0.115 ;
        RECT  9.660 -0.115 9.740 0.335 ;
        RECT  9.530 -0.115 9.660 0.115 ;
        RECT  9.450 -0.115 9.530 0.335 ;
        RECT  9.320 -0.115 9.450 0.115 ;
        RECT  9.240 -0.115 9.320 0.335 ;
        RECT  9.110 -0.115 9.240 0.115 ;
        RECT  9.030 -0.115 9.110 0.335 ;
        RECT  8.900 -0.115 9.030 0.115 ;
        RECT  8.820 -0.115 8.900 0.335 ;
        RECT  8.690 -0.115 8.820 0.115 ;
        RECT  8.610 -0.115 8.690 0.335 ;
        RECT  8.480 -0.115 8.610 0.115 ;
        RECT  8.400 -0.115 8.480 0.335 ;
        RECT  8.270 -0.115 8.400 0.115 ;
        RECT  8.190 -0.115 8.270 0.335 ;
        RECT  8.070 -0.115 8.190 0.115 ;
        RECT  7.990 -0.115 8.070 0.335 ;
        RECT  7.880 -0.115 7.990 0.115 ;
        RECT  7.800 -0.115 7.880 0.335 ;
        RECT  7.690 -0.115 7.800 0.115 ;
        RECT  7.610 -0.115 7.690 0.335 ;
        RECT  7.495 -0.115 7.610 0.115 ;
        RECT  7.415 -0.115 7.495 0.335 ;
        RECT  7.290 -0.115 7.415 0.115 ;
        RECT  7.210 -0.115 7.290 0.335 ;
        RECT  7.080 -0.115 7.210 0.115 ;
        RECT  7.000 -0.115 7.080 0.335 ;
        RECT  6.870 -0.115 7.000 0.115 ;
        RECT  6.790 -0.115 6.870 0.335 ;
        RECT  6.660 -0.115 6.790 0.115 ;
        RECT  6.580 -0.115 6.660 0.335 ;
        RECT  6.450 -0.115 6.580 0.115 ;
        RECT  6.370 -0.115 6.450 0.335 ;
        RECT  6.240 -0.115 6.370 0.115 ;
        RECT  6.160 -0.115 6.240 0.335 ;
        RECT  6.030 -0.115 6.160 0.115 ;
        RECT  5.950 -0.115 6.030 0.335 ;
        RECT  5.830 -0.115 5.950 0.115 ;
        RECT  5.750 -0.115 5.830 0.335 ;
        RECT  5.640 -0.115 5.750 0.115 ;
        RECT  5.560 -0.115 5.640 0.335 ;
        RECT  5.450 -0.115 5.560 0.115 ;
        RECT  5.370 -0.115 5.450 0.335 ;
        RECT  5.270 -0.115 5.370 0.115 ;
        RECT  5.190 -0.115 5.270 0.465 ;
        RECT  4.910 -0.115 5.190 0.115 ;
        RECT  4.790 -0.115 4.910 0.235 ;
        RECT  4.530 -0.115 4.790 0.115 ;
        RECT  4.410 -0.115 4.530 0.235 ;
        RECT  4.150 -0.115 4.410 0.115 ;
        RECT  4.030 -0.115 4.150 0.235 ;
        RECT  3.770 -0.115 4.030 0.115 ;
        RECT  3.650 -0.115 3.770 0.235 ;
        RECT  3.390 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.390 0.235 ;
        RECT  3.010 -0.115 3.270 0.115 ;
        RECT  2.890 -0.115 3.010 0.235 ;
        RECT  2.630 -0.115 2.890 0.115 ;
        RECT  2.510 -0.115 2.630 0.235 ;
        RECT  2.250 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.250 0.235 ;
        RECT  1.870 -0.115 2.130 0.115 ;
        RECT  1.750 -0.115 1.870 0.235 ;
        RECT  1.465 -0.115 1.750 0.115 ;
        RECT  1.395 -0.115 1.465 0.465 ;
        RECT  1.085 -0.115 1.395 0.115 ;
        RECT  1.015 -0.115 1.085 0.255 ;
        RECT  0.695 -0.115 1.015 0.115 ;
        RECT  0.625 -0.115 0.695 0.255 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.245 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.370 1.145 10.640 1.375 ;
        RECT  10.290 0.945 10.370 1.375 ;
        RECT  10.160 1.145 10.290 1.375 ;
        RECT  10.080 0.945 10.160 1.375 ;
        RECT  9.950 1.145 10.080 1.375 ;
        RECT  9.870 0.795 9.950 1.375 ;
        RECT  9.740 1.145 9.870 1.375 ;
        RECT  9.660 0.795 9.740 1.375 ;
        RECT  9.530 1.145 9.660 1.375 ;
        RECT  9.450 0.795 9.530 1.375 ;
        RECT  9.320 1.145 9.450 1.375 ;
        RECT  9.240 0.795 9.320 1.375 ;
        RECT  9.110 1.145 9.240 1.375 ;
        RECT  9.030 0.795 9.110 1.375 ;
        RECT  8.900 1.145 9.030 1.375 ;
        RECT  8.820 0.795 8.900 1.375 ;
        RECT  8.690 1.145 8.820 1.375 ;
        RECT  8.610 0.795 8.690 1.375 ;
        RECT  8.480 1.145 8.610 1.375 ;
        RECT  8.400 0.795 8.480 1.375 ;
        RECT  8.270 1.145 8.400 1.375 ;
        RECT  8.190 0.795 8.270 1.375 ;
        RECT  8.070 1.145 8.190 1.375 ;
        RECT  7.990 0.795 8.070 1.375 ;
        RECT  7.880 1.145 7.990 1.375 ;
        RECT  7.800 0.795 7.880 1.375 ;
        RECT  7.690 1.145 7.800 1.375 ;
        RECT  7.610 0.795 7.690 1.375 ;
        RECT  7.495 1.145 7.610 1.375 ;
        RECT  7.415 0.795 7.495 1.375 ;
        RECT  7.290 1.145 7.415 1.375 ;
        RECT  7.210 0.795 7.290 1.375 ;
        RECT  7.080 1.145 7.210 1.375 ;
        RECT  7.000 0.795 7.080 1.375 ;
        RECT  6.870 1.145 7.000 1.375 ;
        RECT  6.790 0.795 6.870 1.375 ;
        RECT  6.660 1.145 6.790 1.375 ;
        RECT  6.580 0.795 6.660 1.375 ;
        RECT  6.450 1.145 6.580 1.375 ;
        RECT  6.370 0.795 6.450 1.375 ;
        RECT  6.240 1.145 6.370 1.375 ;
        RECT  6.160 0.795 6.240 1.375 ;
        RECT  6.030 1.145 6.160 1.375 ;
        RECT  5.950 0.795 6.030 1.375 ;
        RECT  5.830 1.145 5.950 1.375 ;
        RECT  5.750 0.795 5.830 1.375 ;
        RECT  5.640 1.145 5.750 1.375 ;
        RECT  5.560 0.795 5.640 1.375 ;
        RECT  5.450 1.145 5.560 1.375 ;
        RECT  5.370 0.795 5.450 1.375 ;
        RECT  5.270 1.145 5.370 1.375 ;
        RECT  5.190 0.700 5.270 1.375 ;
        RECT  4.910 1.145 5.190 1.375 ;
        RECT  4.790 1.030 4.910 1.375 ;
        RECT  4.530 1.145 4.790 1.375 ;
        RECT  4.410 1.030 4.530 1.375 ;
        RECT  4.150 1.145 4.410 1.375 ;
        RECT  4.030 1.030 4.150 1.375 ;
        RECT  3.770 1.145 4.030 1.375 ;
        RECT  3.650 1.030 3.770 1.375 ;
        RECT  3.390 1.145 3.650 1.375 ;
        RECT  3.270 1.030 3.390 1.375 ;
        RECT  3.010 1.145 3.270 1.375 ;
        RECT  2.890 1.030 3.010 1.375 ;
        RECT  2.630 1.145 2.890 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.250 1.145 2.510 1.375 ;
        RECT  2.130 1.030 2.250 1.375 ;
        RECT  1.870 1.145 2.130 1.375 ;
        RECT  1.750 1.030 1.870 1.375 ;
        RECT  1.465 1.145 1.750 1.375 ;
        RECT  1.395 0.720 1.465 1.375 ;
        RECT  1.085 1.145 1.395 1.375 ;
        RECT  1.015 1.005 1.085 1.375 ;
        RECT  0.710 1.145 1.015 1.375 ;
        RECT  0.610 1.015 0.710 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.230 1.015 0.330 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.730 5.100 0.960 ;
        RECT  5.005 0.185 5.075 0.465 ;
        RECT  4.695 0.305 5.005 0.465 ;
        RECT  4.625 0.185 4.695 0.465 ;
        RECT  4.315 0.305 4.625 0.465 ;
        RECT  4.245 0.185 4.315 0.465 ;
        RECT  3.935 0.305 4.245 0.465 ;
        RECT  3.865 0.185 3.935 0.465 ;
        RECT  3.605 0.305 3.865 0.465 ;
        RECT  3.105 0.185 3.115 0.465 ;
        RECT  1.560 0.730 3.115 0.960 ;
        RECT  2.795 0.305 3.105 0.465 ;
        RECT  2.725 0.185 2.795 0.465 ;
        RECT  2.415 0.305 2.725 0.465 ;
        RECT  2.345 0.185 2.415 0.465 ;
        RECT  2.035 0.305 2.345 0.465 ;
        RECT  1.965 0.185 2.035 0.465 ;
        RECT  1.655 0.305 1.965 0.465 ;
        RECT  1.585 0.185 1.655 0.465 ;
        RECT  10.510 0.210 10.590 0.710 ;
        RECT  10.510 0.790 10.590 1.060 ;
        RECT  10.250 0.630 10.510 0.710 ;
        RECT  10.180 0.790 10.510 0.870 ;
        RECT  10.100 0.430 10.180 0.870 ;
        RECT  5.525 0.430 10.100 0.510 ;
        RECT  1.315 0.545 3.105 0.615 ;
        RECT  1.155 0.185 1.315 1.065 ;
        RECT  0.895 0.335 1.155 0.415 ;
        RECT  0.920 0.845 1.155 0.925 ;
        RECT  0.800 0.845 0.920 1.065 ;
        RECT  0.825 0.185 0.895 0.415 ;
        RECT  0.505 0.335 0.825 0.415 ;
        RECT  0.530 0.845 0.800 0.925 ;
        RECT  0.410 0.845 0.530 1.075 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.130 0.335 0.435 0.415 ;
        RECT  0.125 0.845 0.410 0.920 ;
        RECT  0.055 0.275 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.075 ;
    END
END DCCKBD20BWP40

MACRO DCCKBD24BWP40
    CLASS CORE ;
    FOREIGN DCCKBD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 1.440000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.155 0.305 4.465 0.465 ;
        RECT  4.095 0.185 4.155 0.465 ;
        RECT  4.085 0.185 4.095 0.945 ;
        RECT  3.775 0.305 4.085 0.945 ;
        RECT  3.745 0.185 3.775 0.945 ;
        RECT  3.705 0.185 3.745 0.465 ;
        RECT  1.780 0.715 3.745 0.945 ;
        RECT  3.395 0.305 3.705 0.465 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.246400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 1.155 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.330 -0.115 12.600 0.115 ;
        RECT  12.250 -0.115 12.330 0.335 ;
        RECT  12.120 -0.115 12.250 0.115 ;
        RECT  12.040 -0.115 12.120 0.335 ;
        RECT  11.890 -0.115 12.040 0.115 ;
        RECT  11.810 -0.115 11.890 0.335 ;
        RECT  11.640 -0.115 11.810 0.115 ;
        RECT  11.560 -0.115 11.640 0.335 ;
        RECT  11.385 -0.115 11.560 0.115 ;
        RECT  11.305 -0.115 11.385 0.335 ;
        RECT  11.140 -0.115 11.305 0.115 ;
        RECT  11.060 -0.115 11.140 0.335 ;
        RECT  10.930 -0.115 11.060 0.115 ;
        RECT  10.850 -0.115 10.930 0.335 ;
        RECT  10.720 -0.115 10.850 0.115 ;
        RECT  10.640 -0.115 10.720 0.335 ;
        RECT  10.510 -0.115 10.640 0.115 ;
        RECT  10.430 -0.115 10.510 0.335 ;
        RECT  10.300 -0.115 10.430 0.115 ;
        RECT  10.220 -0.115 10.300 0.335 ;
        RECT  10.090 -0.115 10.220 0.115 ;
        RECT  10.010 -0.115 10.090 0.335 ;
        RECT  9.880 -0.115 10.010 0.115 ;
        RECT  9.800 -0.115 9.880 0.335 ;
        RECT  9.670 -0.115 9.800 0.115 ;
        RECT  9.590 -0.115 9.670 0.335 ;
        RECT  9.460 -0.115 9.590 0.115 ;
        RECT  9.380 -0.115 9.460 0.335 ;
        RECT  9.250 -0.115 9.380 0.115 ;
        RECT  9.170 -0.115 9.250 0.335 ;
        RECT  9.050 -0.115 9.170 0.115 ;
        RECT  8.970 -0.115 9.050 0.335 ;
        RECT  8.860 -0.115 8.970 0.115 ;
        RECT  8.780 -0.115 8.860 0.335 ;
        RECT  8.670 -0.115 8.780 0.115 ;
        RECT  8.590 -0.115 8.670 0.335 ;
        RECT  8.475 -0.115 8.590 0.115 ;
        RECT  8.395 -0.115 8.475 0.335 ;
        RECT  8.270 -0.115 8.395 0.115 ;
        RECT  8.190 -0.115 8.270 0.335 ;
        RECT  8.060 -0.115 8.190 0.115 ;
        RECT  7.980 -0.115 8.060 0.335 ;
        RECT  7.850 -0.115 7.980 0.115 ;
        RECT  7.770 -0.115 7.850 0.335 ;
        RECT  7.640 -0.115 7.770 0.115 ;
        RECT  7.560 -0.115 7.640 0.335 ;
        RECT  7.430 -0.115 7.560 0.115 ;
        RECT  7.350 -0.115 7.430 0.335 ;
        RECT  7.220 -0.115 7.350 0.115 ;
        RECT  7.140 -0.115 7.220 0.335 ;
        RECT  7.010 -0.115 7.140 0.115 ;
        RECT  6.930 -0.115 7.010 0.335 ;
        RECT  6.810 -0.115 6.930 0.115 ;
        RECT  6.730 -0.115 6.810 0.335 ;
        RECT  6.620 -0.115 6.730 0.115 ;
        RECT  6.540 -0.115 6.620 0.335 ;
        RECT  6.430 -0.115 6.540 0.115 ;
        RECT  6.350 -0.115 6.430 0.335 ;
        RECT  6.250 -0.115 6.350 0.115 ;
        RECT  6.170 -0.115 6.250 0.475 ;
        RECT  5.890 -0.115 6.170 0.115 ;
        RECT  5.770 -0.115 5.890 0.235 ;
        RECT  5.510 -0.115 5.770 0.115 ;
        RECT  5.390 -0.115 5.510 0.235 ;
        RECT  5.130 -0.115 5.390 0.115 ;
        RECT  5.010 -0.115 5.130 0.235 ;
        RECT  4.750 -0.115 5.010 0.115 ;
        RECT  4.630 -0.115 4.750 0.235 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.235 ;
        RECT  3.990 -0.115 4.250 0.115 ;
        RECT  3.870 -0.115 3.990 0.235 ;
        RECT  3.610 -0.115 3.870 0.115 ;
        RECT  3.490 -0.115 3.610 0.235 ;
        RECT  3.230 -0.115 3.490 0.115 ;
        RECT  3.110 -0.115 3.230 0.235 ;
        RECT  2.850 -0.115 3.110 0.115 ;
        RECT  2.730 -0.115 2.850 0.235 ;
        RECT  2.470 -0.115 2.730 0.115 ;
        RECT  2.350 -0.115 2.470 0.235 ;
        RECT  2.090 -0.115 2.350 0.115 ;
        RECT  1.970 -0.115 2.090 0.235 ;
        RECT  1.685 -0.115 1.970 0.115 ;
        RECT  1.615 -0.115 1.685 0.465 ;
        RECT  1.295 -0.115 1.615 0.115 ;
        RECT  1.225 -0.115 1.295 0.245 ;
        RECT  0.895 -0.115 1.225 0.115 ;
        RECT  0.825 -0.115 0.895 0.245 ;
        RECT  0.505 -0.115 0.825 0.115 ;
        RECT  0.435 -0.115 0.505 0.245 ;
        RECT  0.125 -0.115 0.435 0.115 ;
        RECT  0.055 -0.115 0.125 0.415 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.330 1.145 12.600 1.375 ;
        RECT  12.250 0.945 12.330 1.375 ;
        RECT  12.120 1.145 12.250 1.375 ;
        RECT  12.040 0.945 12.120 1.375 ;
        RECT  11.890 1.145 12.040 1.375 ;
        RECT  11.810 0.795 11.890 1.375 ;
        RECT  11.640 1.145 11.810 1.375 ;
        RECT  11.560 0.795 11.640 1.375 ;
        RECT  11.385 1.145 11.560 1.375 ;
        RECT  11.305 0.795 11.385 1.375 ;
        RECT  11.140 1.145 11.305 1.375 ;
        RECT  11.060 0.795 11.140 1.375 ;
        RECT  10.930 1.145 11.060 1.375 ;
        RECT  10.850 0.795 10.930 1.375 ;
        RECT  10.720 1.145 10.850 1.375 ;
        RECT  10.640 0.795 10.720 1.375 ;
        RECT  10.510 1.145 10.640 1.375 ;
        RECT  10.430 0.795 10.510 1.375 ;
        RECT  10.300 1.145 10.430 1.375 ;
        RECT  10.220 0.795 10.300 1.375 ;
        RECT  10.090 1.145 10.220 1.375 ;
        RECT  10.010 0.795 10.090 1.375 ;
        RECT  9.880 1.145 10.010 1.375 ;
        RECT  9.800 0.795 9.880 1.375 ;
        RECT  9.670 1.145 9.800 1.375 ;
        RECT  9.590 0.795 9.670 1.375 ;
        RECT  9.460 1.145 9.590 1.375 ;
        RECT  9.380 0.795 9.460 1.375 ;
        RECT  9.250 1.145 9.380 1.375 ;
        RECT  9.170 0.795 9.250 1.375 ;
        RECT  9.050 1.145 9.170 1.375 ;
        RECT  8.970 0.795 9.050 1.375 ;
        RECT  8.860 1.145 8.970 1.375 ;
        RECT  8.780 0.795 8.860 1.375 ;
        RECT  8.670 1.145 8.780 1.375 ;
        RECT  8.590 0.795 8.670 1.375 ;
        RECT  8.475 1.145 8.590 1.375 ;
        RECT  8.395 0.795 8.475 1.375 ;
        RECT  8.270 1.145 8.395 1.375 ;
        RECT  8.190 0.795 8.270 1.375 ;
        RECT  8.060 1.145 8.190 1.375 ;
        RECT  7.980 0.795 8.060 1.375 ;
        RECT  7.850 1.145 7.980 1.375 ;
        RECT  7.770 0.795 7.850 1.375 ;
        RECT  7.640 1.145 7.770 1.375 ;
        RECT  7.560 0.795 7.640 1.375 ;
        RECT  7.430 1.145 7.560 1.375 ;
        RECT  7.350 0.795 7.430 1.375 ;
        RECT  7.220 1.145 7.350 1.375 ;
        RECT  7.140 0.795 7.220 1.375 ;
        RECT  7.010 1.145 7.140 1.375 ;
        RECT  6.930 0.795 7.010 1.375 ;
        RECT  6.810 1.145 6.930 1.375 ;
        RECT  6.730 0.795 6.810 1.375 ;
        RECT  6.620 1.145 6.730 1.375 ;
        RECT  6.540 0.795 6.620 1.375 ;
        RECT  6.430 1.145 6.540 1.375 ;
        RECT  6.350 0.795 6.430 1.375 ;
        RECT  6.250 1.145 6.350 1.375 ;
        RECT  6.170 0.720 6.250 1.375 ;
        RECT  5.890 1.145 6.170 1.375 ;
        RECT  5.770 1.015 5.890 1.375 ;
        RECT  5.510 1.145 5.770 1.375 ;
        RECT  5.390 1.015 5.510 1.375 ;
        RECT  5.130 1.145 5.390 1.375 ;
        RECT  5.010 1.015 5.130 1.375 ;
        RECT  4.750 1.145 5.010 1.375 ;
        RECT  4.630 1.015 4.750 1.375 ;
        RECT  4.370 1.145 4.630 1.375 ;
        RECT  4.250 1.015 4.370 1.375 ;
        RECT  3.990 1.145 4.250 1.375 ;
        RECT  3.870 1.015 3.990 1.375 ;
        RECT  3.610 1.145 3.870 1.375 ;
        RECT  3.490 1.015 3.610 1.375 ;
        RECT  3.230 1.145 3.490 1.375 ;
        RECT  3.110 1.015 3.230 1.375 ;
        RECT  2.850 1.145 3.110 1.375 ;
        RECT  2.730 1.015 2.850 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 1.015 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 1.015 2.090 1.375 ;
        RECT  1.685 1.145 1.970 1.375 ;
        RECT  1.615 0.740 1.685 1.375 ;
        RECT  1.295 1.145 1.615 1.375 ;
        RECT  1.225 0.880 1.295 1.375 ;
        RECT  0.900 1.145 1.225 1.375 ;
        RECT  0.820 0.880 0.900 1.375 ;
        RECT  0.510 1.145 0.820 1.375 ;
        RECT  0.430 0.880 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.165 0.715 6.080 0.945 ;
        RECT  5.985 0.185 6.055 0.465 ;
        RECT  5.675 0.305 5.985 0.465 ;
        RECT  5.605 0.185 5.675 0.465 ;
        RECT  5.295 0.305 5.605 0.465 ;
        RECT  5.225 0.185 5.295 0.465 ;
        RECT  4.915 0.305 5.225 0.465 ;
        RECT  4.845 0.185 4.915 0.465 ;
        RECT  4.535 0.305 4.845 0.465 ;
        RECT  4.465 0.185 4.535 0.465 ;
        RECT  4.165 0.305 4.465 0.465 ;
        RECT  3.395 0.305 3.675 0.465 ;
        RECT  1.780 0.715 3.675 0.945 ;
        RECT  3.325 0.185 3.395 0.465 ;
        RECT  3.015 0.305 3.325 0.465 ;
        RECT  2.945 0.185 3.015 0.465 ;
        RECT  2.635 0.305 2.945 0.465 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.305 2.565 0.465 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.875 0.305 2.185 0.465 ;
        RECT  1.805 0.185 1.875 0.465 ;
        RECT  12.470 0.210 12.550 0.710 ;
        RECT  12.470 0.790 12.550 1.060 ;
        RECT  12.210 0.630 12.470 0.710 ;
        RECT  12.140 0.790 12.470 0.870 ;
        RECT  12.060 0.430 12.140 0.870 ;
        RECT  6.505 0.430 12.060 0.510 ;
        RECT  1.535 0.545 3.645 0.615 ;
        RECT  1.365 0.195 1.535 1.070 ;
        RECT  1.100 0.325 1.365 0.415 ;
        RECT  1.120 0.705 1.365 0.795 ;
        RECT  1.000 0.705 1.120 1.070 ;
        RECT  1.020 0.185 1.100 0.415 ;
        RECT  0.700 0.325 1.020 0.415 ;
        RECT  0.720 0.705 1.000 0.795 ;
        RECT  0.600 0.705 0.720 1.070 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.320 0.325 0.620 0.415 ;
        RECT  0.340 0.705 0.600 0.795 ;
        RECT  0.220 0.705 0.340 1.065 ;
        RECT  0.220 0.185 0.320 0.415 ;
    END
END DCCKBD24BWP40

MACRO DCCKBD4BWP40
    CLASS CORE ;
    FOREIGN DCCKBD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.185 1.125 0.465 ;
        RECT  1.055 0.700 1.125 1.045 ;
        RECT  1.015 0.355 1.055 0.465 ;
        RECT  1.015 0.700 1.055 0.820 ;
        RECT  0.805 0.355 1.015 0.820 ;
        RECT  0.725 0.355 0.805 0.465 ;
        RECT  0.725 0.700 0.805 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.280 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.115 2.800 0.115 ;
        RECT  2.450 -0.115 2.530 0.335 ;
        RECT  2.320 -0.115 2.450 0.115 ;
        RECT  2.240 -0.115 2.320 0.335 ;
        RECT  2.110 -0.115 2.240 0.115 ;
        RECT  2.030 -0.115 2.110 0.335 ;
        RECT  1.910 -0.115 2.030 0.115 ;
        RECT  1.830 -0.115 1.910 0.335 ;
        RECT  1.720 -0.115 1.830 0.115 ;
        RECT  1.640 -0.115 1.720 0.335 ;
        RECT  1.530 -0.115 1.640 0.115 ;
        RECT  1.450 -0.115 1.530 0.335 ;
        RECT  1.350 -0.115 1.450 0.115 ;
        RECT  1.270 -0.115 1.350 0.475 ;
        RECT  0.950 -0.115 1.270 0.115 ;
        RECT  0.830 -0.115 0.950 0.280 ;
        RECT  0.530 -0.115 0.830 0.115 ;
        RECT  0.450 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.450 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.145 2.800 1.375 ;
        RECT  2.450 0.945 2.530 1.375 ;
        RECT  2.320 1.145 2.450 1.375 ;
        RECT  2.240 0.945 2.320 1.375 ;
        RECT  2.110 1.145 2.240 1.375 ;
        RECT  2.030 0.795 2.110 1.375 ;
        RECT  1.910 1.145 2.030 1.375 ;
        RECT  1.830 0.795 1.910 1.375 ;
        RECT  1.720 1.145 1.830 1.375 ;
        RECT  1.640 0.795 1.720 1.375 ;
        RECT  1.530 1.145 1.640 1.375 ;
        RECT  1.450 0.795 1.530 1.375 ;
        RECT  1.350 1.145 1.450 1.375 ;
        RECT  1.270 0.700 1.350 1.375 ;
        RECT  0.950 1.145 1.270 1.375 ;
        RECT  0.830 0.890 0.950 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.440 0.975 0.540 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.185 1.125 0.465 ;
        RECT  1.085 0.700 1.125 1.045 ;
        RECT  0.725 0.355 0.735 0.465 ;
        RECT  0.725 0.700 0.735 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  2.670 0.210 2.750 0.710 ;
        RECT  2.670 0.790 2.750 1.060 ;
        RECT  2.410 0.630 2.670 0.710 ;
        RECT  2.340 0.790 2.670 0.870 ;
        RECT  2.260 0.430 2.340 0.870 ;
        RECT  1.605 0.430 2.260 0.510 ;
        RECT  0.585 0.545 0.720 0.615 ;
        RECT  0.510 0.345 0.585 0.905 ;
        RECT  0.325 0.345 0.510 0.415 ;
        RECT  0.325 0.835 0.510 0.905 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.835 0.325 0.995 ;
    END
END DCCKBD4BWP40

MACRO DCCKBD5BWP40
    CLASS CORE ;
    FOREIGN DCCKBD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.340000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.155 0.355 1.415 0.465 ;
        RECT  1.155 0.700 1.415 0.820 ;
        RECT  1.105 0.355 1.155 0.820 ;
        RECT  1.085 0.355 1.105 1.045 ;
        RECT  1.015 0.185 1.085 1.045 ;
        RECT  0.945 0.355 1.015 0.820 ;
        RECT  0.695 0.355 0.945 0.465 ;
        RECT  0.695 0.700 0.945 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.063200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.385 0.635 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.810 -0.115 3.080 0.115 ;
        RECT  2.730 -0.115 2.810 0.335 ;
        RECT  2.600 -0.115 2.730 0.115 ;
        RECT  2.520 -0.115 2.600 0.335 ;
        RECT  2.390 -0.115 2.520 0.115 ;
        RECT  2.310 -0.115 2.390 0.335 ;
        RECT  2.155 -0.115 2.310 0.115 ;
        RECT  2.075 -0.115 2.155 0.335 ;
        RECT  1.860 -0.115 2.075 0.115 ;
        RECT  1.780 -0.115 1.860 0.335 ;
        RECT  1.670 -0.115 1.780 0.115 ;
        RECT  1.590 -0.115 1.670 0.335 ;
        RECT  1.320 -0.115 1.590 0.115 ;
        RECT  1.200 -0.115 1.320 0.280 ;
        RECT  0.920 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.920 0.280 ;
        RECT  0.510 -0.115 0.800 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.145 3.080 1.375 ;
        RECT  2.730 0.945 2.810 1.375 ;
        RECT  2.600 1.145 2.730 1.375 ;
        RECT  2.520 0.945 2.600 1.375 ;
        RECT  2.390 1.145 2.520 1.375 ;
        RECT  2.310 0.795 2.390 1.375 ;
        RECT  2.155 1.145 2.310 1.375 ;
        RECT  2.075 0.795 2.155 1.375 ;
        RECT  1.860 1.145 2.075 1.375 ;
        RECT  1.780 0.795 1.860 1.375 ;
        RECT  1.670 1.145 1.780 1.375 ;
        RECT  1.590 0.795 1.670 1.375 ;
        RECT  1.320 1.145 1.590 1.375 ;
        RECT  1.200 0.890 1.320 1.375 ;
        RECT  0.920 1.145 1.200 1.375 ;
        RECT  0.800 0.890 0.920 1.375 ;
        RECT  0.530 1.145 0.800 1.375 ;
        RECT  0.410 0.890 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.860 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.485 0.465 ;
        RECT  1.415 0.700 1.485 1.045 ;
        RECT  1.225 0.355 1.415 0.465 ;
        RECT  1.225 0.700 1.415 0.820 ;
        RECT  0.695 0.355 0.875 0.465 ;
        RECT  0.695 0.700 0.875 0.820 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.700 0.695 1.045 ;
        RECT  2.950 0.210 3.030 0.710 ;
        RECT  2.950 0.790 3.030 1.060 ;
        RECT  2.690 0.630 2.950 0.710 ;
        RECT  2.620 0.790 2.950 0.870 ;
        RECT  2.540 0.430 2.620 0.870 ;
        RECT  1.745 0.430 2.540 0.510 ;
        RECT  0.535 0.545 0.825 0.615 ;
        RECT  0.465 0.345 0.535 0.820 ;
        RECT  0.315 0.345 0.465 0.415 ;
        RECT  0.315 0.750 0.465 0.820 ;
        RECT  0.245 0.245 0.315 0.415 ;
        RECT  0.245 0.750 0.315 0.995 ;
    END
END DCCKBD5BWP40

MACRO DCCKBD6BWP40
    CLASS CORE ;
    FOREIGN DCCKBD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.384000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.155 0.355 1.455 0.465 ;
        RECT  1.155 0.700 1.455 0.820 ;
        RECT  1.145 0.355 1.155 0.820 ;
        RECT  1.125 0.355 1.145 1.045 ;
        RECT  1.055 0.185 1.125 1.045 ;
        RECT  0.945 0.355 1.055 0.820 ;
        RECT  0.725 0.355 0.945 0.465 ;
        RECT  0.725 0.700 0.945 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.385 0.635 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 -0.115 3.640 0.115 ;
        RECT  3.290 -0.115 3.370 0.335 ;
        RECT  3.160 -0.115 3.290 0.115 ;
        RECT  3.080 -0.115 3.160 0.335 ;
        RECT  2.950 -0.115 3.080 0.115 ;
        RECT  2.870 -0.115 2.950 0.335 ;
        RECT  2.740 -0.115 2.870 0.115 ;
        RECT  2.660 -0.115 2.740 0.335 ;
        RECT  2.530 -0.115 2.660 0.115 ;
        RECT  2.450 -0.115 2.530 0.335 ;
        RECT  2.330 -0.115 2.450 0.115 ;
        RECT  2.250 -0.115 2.330 0.335 ;
        RECT  2.140 -0.115 2.250 0.115 ;
        RECT  2.060 -0.115 2.140 0.335 ;
        RECT  1.950 -0.115 2.060 0.115 ;
        RECT  1.870 -0.115 1.950 0.335 ;
        RECT  1.770 -0.115 1.870 0.115 ;
        RECT  1.690 -0.115 1.770 0.465 ;
        RECT  1.360 -0.115 1.690 0.115 ;
        RECT  1.240 -0.115 1.360 0.280 ;
        RECT  0.960 -0.115 1.240 0.115 ;
        RECT  0.840 -0.115 0.960 0.280 ;
        RECT  0.540 -0.115 0.840 0.115 ;
        RECT  0.460 -0.115 0.540 0.270 ;
        RECT  0.140 -0.115 0.460 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.145 3.640 1.375 ;
        RECT  3.290 0.945 3.370 1.375 ;
        RECT  3.160 1.145 3.290 1.375 ;
        RECT  3.080 0.945 3.160 1.375 ;
        RECT  2.950 1.145 3.080 1.375 ;
        RECT  2.870 0.795 2.950 1.375 ;
        RECT  2.740 1.145 2.870 1.375 ;
        RECT  2.660 0.795 2.740 1.375 ;
        RECT  2.530 1.145 2.660 1.375 ;
        RECT  2.450 0.795 2.530 1.375 ;
        RECT  2.330 1.145 2.450 1.375 ;
        RECT  2.250 0.795 2.330 1.375 ;
        RECT  2.140 1.145 2.250 1.375 ;
        RECT  2.060 0.795 2.140 1.375 ;
        RECT  1.950 1.145 2.060 1.375 ;
        RECT  1.870 0.795 1.950 1.375 ;
        RECT  1.770 1.145 1.870 1.375 ;
        RECT  1.690 0.735 1.770 1.375 ;
        RECT  1.360 1.145 1.690 1.375 ;
        RECT  1.240 0.890 1.360 1.375 ;
        RECT  0.960 1.145 1.240 1.375 ;
        RECT  0.840 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.000 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.455 0.185 1.525 0.465 ;
        RECT  1.455 0.700 1.525 1.045 ;
        RECT  1.225 0.355 1.455 0.465 ;
        RECT  1.225 0.700 1.455 0.820 ;
        RECT  0.725 0.355 0.875 0.465 ;
        RECT  0.725 0.700 0.875 0.820 ;
        RECT  0.655 0.185 0.725 0.465 ;
        RECT  0.655 0.700 0.725 1.045 ;
        RECT  3.510 0.210 3.590 0.710 ;
        RECT  3.510 0.790 3.590 1.060 ;
        RECT  3.250 0.630 3.510 0.710 ;
        RECT  3.180 0.790 3.510 0.870 ;
        RECT  3.100 0.430 3.180 0.870 ;
        RECT  2.025 0.430 3.100 0.510 ;
        RECT  0.565 0.545 0.865 0.615 ;
        RECT  0.485 0.345 0.565 0.915 ;
        RECT  0.325 0.345 0.485 0.415 ;
        RECT  0.325 0.845 0.485 0.915 ;
        RECT  0.255 0.245 0.325 0.415 ;
        RECT  0.255 0.845 0.325 0.995 ;
    END
END DCCKBD6BWP40

MACRO DCCKBD8BWP40
    CLASS CORE ;
    FOREIGN DCCKBD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.512000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.765 0.305 2.055 0.465 ;
        RECT  1.715 0.185 1.765 0.465 ;
        RECT  1.655 0.185 1.715 0.950 ;
        RECT  1.365 0.305 1.655 0.950 ;
        RECT  1.325 0.305 1.365 0.465 ;
        RECT  0.825 0.720 1.365 0.950 ;
        RECT  1.235 0.185 1.325 0.465 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.092400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.495 0.300 0.625 ;
        RECT  0.035 0.495 0.120 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.490 -0.115 4.760 0.115 ;
        RECT  4.410 -0.115 4.490 0.335 ;
        RECT  4.280 -0.115 4.410 0.115 ;
        RECT  4.200 -0.115 4.280 0.335 ;
        RECT  4.045 -0.115 4.200 0.115 ;
        RECT  3.965 -0.115 4.045 0.335 ;
        RECT  3.790 -0.115 3.965 0.115 ;
        RECT  3.710 -0.115 3.790 0.335 ;
        RECT  3.535 -0.115 3.710 0.115 ;
        RECT  3.455 -0.115 3.535 0.335 ;
        RECT  3.300 -0.115 3.455 0.115 ;
        RECT  3.220 -0.115 3.300 0.335 ;
        RECT  3.090 -0.115 3.220 0.115 ;
        RECT  3.010 -0.115 3.090 0.335 ;
        RECT  2.890 -0.115 3.010 0.115 ;
        RECT  2.810 -0.115 2.890 0.335 ;
        RECT  2.700 -0.115 2.810 0.115 ;
        RECT  2.620 -0.115 2.700 0.335 ;
        RECT  2.510 -0.115 2.620 0.115 ;
        RECT  2.430 -0.115 2.510 0.335 ;
        RECT  2.330 -0.115 2.430 0.115 ;
        RECT  2.250 -0.115 2.330 0.465 ;
        RECT  1.960 -0.115 2.250 0.115 ;
        RECT  1.840 -0.115 1.960 0.235 ;
        RECT  1.560 -0.115 1.840 0.115 ;
        RECT  1.440 -0.115 1.560 0.235 ;
        RECT  1.160 -0.115 1.440 0.115 ;
        RECT  1.040 -0.115 1.160 0.235 ;
        RECT  0.730 -0.115 1.040 0.115 ;
        RECT  0.650 -0.115 0.730 0.465 ;
        RECT  0.360 -0.115 0.650 0.115 ;
        RECT  0.240 -0.115 0.360 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.490 1.145 4.760 1.375 ;
        RECT  4.410 0.945 4.490 1.375 ;
        RECT  4.280 1.145 4.410 1.375 ;
        RECT  4.200 0.945 4.280 1.375 ;
        RECT  4.045 1.145 4.200 1.375 ;
        RECT  3.965 0.795 4.045 1.375 ;
        RECT  3.790 1.145 3.965 1.375 ;
        RECT  3.710 0.795 3.790 1.375 ;
        RECT  3.535 1.145 3.710 1.375 ;
        RECT  3.455 0.795 3.535 1.375 ;
        RECT  3.300 1.145 3.455 1.375 ;
        RECT  3.220 0.795 3.300 1.375 ;
        RECT  3.090 1.145 3.220 1.375 ;
        RECT  3.010 0.795 3.090 1.375 ;
        RECT  2.890 1.145 3.010 1.375 ;
        RECT  2.810 0.795 2.890 1.375 ;
        RECT  2.700 1.145 2.810 1.375 ;
        RECT  2.620 0.795 2.700 1.375 ;
        RECT  2.510 1.145 2.620 1.375 ;
        RECT  2.430 0.795 2.510 1.375 ;
        RECT  2.330 1.145 2.430 1.375 ;
        RECT  2.250 0.700 2.330 1.375 ;
        RECT  1.960 1.145 2.250 1.375 ;
        RECT  1.840 1.020 1.960 1.375 ;
        RECT  1.560 1.145 1.840 1.375 ;
        RECT  1.440 1.020 1.560 1.375 ;
        RECT  1.160 1.145 1.440 1.375 ;
        RECT  1.040 1.020 1.160 1.375 ;
        RECT  0.730 1.145 1.040 1.375 ;
        RECT  0.650 0.700 0.730 1.375 ;
        RECT  0.360 1.145 0.650 1.375 ;
        RECT  0.240 1.015 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.720 2.155 0.950 ;
        RECT  2.055 0.185 2.125 0.465 ;
        RECT  1.785 0.305 2.055 0.465 ;
        RECT  1.235 0.185 1.295 0.465 ;
        RECT  0.825 0.720 1.295 0.950 ;
        RECT  0.925 0.305 1.235 0.465 ;
        RECT  0.855 0.185 0.925 0.465 ;
        RECT  4.630 0.210 4.710 0.710 ;
        RECT  4.630 0.790 4.710 1.060 ;
        RECT  4.370 0.630 4.630 0.710 ;
        RECT  4.300 0.790 4.630 0.870 ;
        RECT  4.220 0.430 4.300 0.870 ;
        RECT  2.585 0.430 4.220 0.510 ;
        RECT  0.535 0.545 1.215 0.615 ;
        RECT  0.445 0.185 0.535 1.055 ;
        RECT  0.125 0.335 0.445 0.415 ;
        RECT  0.125 0.850 0.445 0.930 ;
        RECT  0.055 0.245 0.125 0.415 ;
        RECT  0.055 0.850 0.125 1.035 ;
    END
END DCCKBD8BWP40

MACRO DCCKND10BWP40
    CLASS CORE ;
    FOREIGN DCCKND10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.510000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.405 0.695 1.505 1.045 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.155 0.300 1.405 0.465 ;
        RECT  1.155 0.695 1.405 0.885 ;
        RECT  1.095 0.300 1.155 0.885 ;
        RECT  1.015 0.185 1.095 1.045 ;
        RECT  0.945 0.300 1.015 0.885 ;
        RECT  0.715 0.300 0.945 0.465 ;
        RECT  0.715 0.695 0.945 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.272000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.840 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 -0.115 4.200 0.115 ;
        RECT  3.850 -0.115 3.930 0.335 ;
        RECT  3.720 -0.115 3.850 0.115 ;
        RECT  3.640 -0.115 3.720 0.335 ;
        RECT  3.510 -0.115 3.640 0.115 ;
        RECT  3.430 -0.115 3.510 0.335 ;
        RECT  3.255 -0.115 3.430 0.115 ;
        RECT  3.175 -0.115 3.255 0.335 ;
        RECT  3.020 -0.115 3.175 0.115 ;
        RECT  2.940 -0.115 3.020 0.335 ;
        RECT  2.810 -0.115 2.940 0.115 ;
        RECT  2.730 -0.115 2.810 0.335 ;
        RECT  2.610 -0.115 2.730 0.115 ;
        RECT  2.530 -0.115 2.610 0.335 ;
        RECT  2.420 -0.115 2.530 0.115 ;
        RECT  2.340 -0.115 2.420 0.335 ;
        RECT  2.230 -0.115 2.340 0.115 ;
        RECT  2.150 -0.115 2.230 0.335 ;
        RECT  2.045 -0.115 2.150 0.115 ;
        RECT  1.975 -0.115 2.045 0.335 ;
        RECT  1.690 -0.115 1.975 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.290 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.145 4.200 1.375 ;
        RECT  3.850 0.945 3.930 1.375 ;
        RECT  3.720 1.145 3.850 1.375 ;
        RECT  3.640 0.945 3.720 1.375 ;
        RECT  3.510 1.145 3.640 1.375 ;
        RECT  3.430 0.795 3.510 1.375 ;
        RECT  3.255 1.145 3.430 1.375 ;
        RECT  3.175 0.795 3.255 1.375 ;
        RECT  3.020 1.145 3.175 1.375 ;
        RECT  2.940 0.795 3.020 1.375 ;
        RECT  2.810 1.145 2.940 1.375 ;
        RECT  2.730 0.795 2.810 1.375 ;
        RECT  2.610 1.145 2.730 1.375 ;
        RECT  2.530 0.795 2.610 1.375 ;
        RECT  2.420 1.145 2.530 1.375 ;
        RECT  2.340 0.795 2.420 1.375 ;
        RECT  2.230 1.145 2.340 1.375 ;
        RECT  2.150 0.795 2.230 1.375 ;
        RECT  2.050 1.145 2.150 1.375 ;
        RECT  1.970 0.685 2.050 1.375 ;
        RECT  1.690 1.145 1.970 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.405 0.695 1.505 1.045 ;
        RECT  1.405 0.185 1.475 0.465 ;
        RECT  1.225 0.300 1.405 0.465 ;
        RECT  1.225 0.695 1.405 0.885 ;
        RECT  0.715 0.300 0.875 0.465 ;
        RECT  0.715 0.695 0.875 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        RECT  4.070 0.210 4.150 0.710 ;
        RECT  4.070 0.790 4.150 1.060 ;
        RECT  3.810 0.630 4.070 0.710 ;
        RECT  3.740 0.790 4.070 0.870 ;
        RECT  3.660 0.430 3.740 0.870 ;
        RECT  2.305 0.430 3.660 0.510 ;
    END
END DCCKND10BWP40

MACRO DCCKND12BWP40
    CLASS CORE ;
    FOREIGN DCCKND12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.612000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.435 0.695 1.505 1.045 ;
        RECT  1.435 0.185 1.475 0.465 ;
        RECT  1.405 0.185 1.435 1.045 ;
        RECT  1.095 0.300 1.405 0.885 ;
        RECT  1.085 0.185 1.095 1.035 ;
        RECT  1.025 0.185 1.085 0.465 ;
        RECT  1.025 0.695 1.085 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.326400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.855 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.770 -0.115 5.040 0.115 ;
        RECT  4.690 -0.115 4.770 0.335 ;
        RECT  4.560 -0.115 4.690 0.115 ;
        RECT  4.480 -0.115 4.560 0.335 ;
        RECT  4.325 -0.115 4.480 0.115 ;
        RECT  4.245 -0.115 4.325 0.335 ;
        RECT  4.120 -0.115 4.245 0.115 ;
        RECT  4.040 -0.115 4.120 0.335 ;
        RECT  3.890 -0.115 4.040 0.115 ;
        RECT  3.810 -0.115 3.890 0.335 ;
        RECT  3.675 -0.115 3.810 0.115 ;
        RECT  3.595 -0.115 3.675 0.335 ;
        RECT  3.440 -0.115 3.595 0.115 ;
        RECT  3.360 -0.115 3.440 0.335 ;
        RECT  3.230 -0.115 3.360 0.115 ;
        RECT  3.150 -0.115 3.230 0.335 ;
        RECT  3.030 -0.115 3.150 0.115 ;
        RECT  2.950 -0.115 3.030 0.335 ;
        RECT  2.840 -0.115 2.950 0.115 ;
        RECT  2.760 -0.115 2.840 0.335 ;
        RECT  2.650 -0.115 2.760 0.115 ;
        RECT  2.570 -0.115 2.650 0.335 ;
        RECT  2.425 -0.115 2.570 0.115 ;
        RECT  2.355 -0.115 2.425 0.325 ;
        RECT  2.070 -0.115 2.355 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.310 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.770 1.145 5.040 1.375 ;
        RECT  4.690 0.945 4.770 1.375 ;
        RECT  4.560 1.145 4.690 1.375 ;
        RECT  4.480 0.945 4.560 1.375 ;
        RECT  4.325 1.145 4.480 1.375 ;
        RECT  4.245 0.795 4.325 1.375 ;
        RECT  4.120 1.145 4.245 1.375 ;
        RECT  4.040 0.795 4.120 1.375 ;
        RECT  3.890 1.145 4.040 1.375 ;
        RECT  3.810 0.795 3.890 1.375 ;
        RECT  3.675 1.145 3.810 1.375 ;
        RECT  3.595 0.795 3.675 1.375 ;
        RECT  3.440 1.145 3.595 1.375 ;
        RECT  3.360 0.795 3.440 1.375 ;
        RECT  3.230 1.145 3.360 1.375 ;
        RECT  3.150 0.795 3.230 1.375 ;
        RECT  3.030 1.145 3.150 1.375 ;
        RECT  2.950 0.795 3.030 1.375 ;
        RECT  2.840 1.145 2.950 1.375 ;
        RECT  2.760 0.795 2.840 1.375 ;
        RECT  2.650 1.145 2.760 1.375 ;
        RECT  2.570 0.795 2.650 1.375 ;
        RECT  2.435 1.145 2.570 1.375 ;
        RECT  2.355 0.670 2.435 1.375 ;
        RECT  2.070 1.145 2.355 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.505 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  0.715 0.300 1.015 0.465 ;
        RECT  0.715 0.695 1.015 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        RECT  4.910 0.210 4.990 0.710 ;
        RECT  4.910 0.790 4.990 1.060 ;
        RECT  4.650 0.630 4.910 0.710 ;
        RECT  4.580 0.790 4.910 0.870 ;
        RECT  4.500 0.430 4.580 0.870 ;
        RECT  2.725 0.430 4.500 0.510 ;
    END
END DCCKND12BWP40

MACRO DCCKND14BWP40
    CLASS CORE ;
    FOREIGN DCCKND14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.737800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.595 0.300 1.785 0.465 ;
        RECT  1.595 0.695 1.785 0.885 ;
        RECT  1.505 0.300 1.595 0.885 ;
        RECT  1.475 0.300 1.505 1.045 ;
        RECT  1.405 0.185 1.475 1.045 ;
        RECT  1.225 0.300 1.405 0.885 ;
        RECT  1.095 0.300 1.225 0.465 ;
        RECT  1.095 0.695 1.225 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.380800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.045 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.610 -0.115 5.880 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.170 -0.115 5.320 0.115 ;
        RECT  5.090 -0.115 5.170 0.335 ;
        RECT  4.935 -0.115 5.090 0.115 ;
        RECT  4.855 -0.115 4.935 0.335 ;
        RECT  4.700 -0.115 4.855 0.115 ;
        RECT  4.620 -0.115 4.700 0.335 ;
        RECT  4.490 -0.115 4.620 0.115 ;
        RECT  4.410 -0.115 4.490 0.335 ;
        RECT  4.280 -0.115 4.410 0.115 ;
        RECT  4.200 -0.115 4.280 0.335 ;
        RECT  4.070 -0.115 4.200 0.115 ;
        RECT  3.990 -0.115 4.070 0.335 ;
        RECT  3.860 -0.115 3.990 0.115 ;
        RECT  3.780 -0.115 3.860 0.335 ;
        RECT  3.650 -0.115 3.780 0.115 ;
        RECT  3.570 -0.115 3.650 0.335 ;
        RECT  3.450 -0.115 3.570 0.115 ;
        RECT  3.370 -0.115 3.450 0.335 ;
        RECT  3.260 -0.115 3.370 0.115 ;
        RECT  3.180 -0.115 3.260 0.335 ;
        RECT  3.070 -0.115 3.180 0.115 ;
        RECT  2.990 -0.115 3.070 0.335 ;
        RECT  2.840 -0.115 2.990 0.115 ;
        RECT  2.750 -0.115 2.840 0.350 ;
        RECT  2.450 -0.115 2.750 0.115 ;
        RECT  2.330 -0.115 2.450 0.230 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.315 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.610 1.145 5.880 1.375 ;
        RECT  5.530 0.945 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.945 5.400 1.375 ;
        RECT  5.170 1.145 5.320 1.375 ;
        RECT  5.090 0.795 5.170 1.375 ;
        RECT  4.935 1.145 5.090 1.375 ;
        RECT  4.855 0.795 4.935 1.375 ;
        RECT  4.700 1.145 4.855 1.375 ;
        RECT  4.620 0.795 4.700 1.375 ;
        RECT  4.490 1.145 4.620 1.375 ;
        RECT  4.410 0.795 4.490 1.375 ;
        RECT  4.280 1.145 4.410 1.375 ;
        RECT  4.200 0.795 4.280 1.375 ;
        RECT  4.070 1.145 4.200 1.375 ;
        RECT  3.990 0.795 4.070 1.375 ;
        RECT  3.860 1.145 3.990 1.375 ;
        RECT  3.780 0.795 3.860 1.375 ;
        RECT  3.650 1.145 3.780 1.375 ;
        RECT  3.570 0.795 3.650 1.375 ;
        RECT  3.450 1.145 3.570 1.375 ;
        RECT  3.370 0.795 3.450 1.375 ;
        RECT  3.260 1.145 3.370 1.375 ;
        RECT  3.180 0.795 3.260 1.375 ;
        RECT  3.070 1.145 3.180 1.375 ;
        RECT  2.990 0.795 3.070 1.375 ;
        RECT  2.845 1.145 2.990 1.375 ;
        RECT  2.755 0.685 2.845 1.375 ;
        RECT  2.450 1.145 2.755 1.375 ;
        RECT  2.330 0.955 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.645 0.300 1.785 0.465 ;
        RECT  1.645 0.695 1.785 0.885 ;
        RECT  1.095 0.300 1.155 0.465 ;
        RECT  1.095 0.695 1.155 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        RECT  5.750 0.210 5.830 0.710 ;
        RECT  5.750 0.790 5.830 1.060 ;
        RECT  5.490 0.630 5.750 0.710 ;
        RECT  5.420 0.790 5.750 0.870 ;
        RECT  5.340 0.430 5.420 0.870 ;
        RECT  3.145 0.430 5.340 0.510 ;
    END
END DCCKND14BWP40

MACRO DCCKND16BWP40
    CLASS CORE ;
    FOREIGN DCCKND16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.816000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.715 0.300 1.765 0.465 ;
        RECT  1.715 0.695 1.765 0.885 ;
        RECT  1.505 0.300 1.715 0.885 ;
        RECT  1.455 0.300 1.505 1.045 ;
        RECT  1.385 0.185 1.455 1.045 ;
        RECT  1.365 0.300 1.385 0.885 ;
        RECT  1.075 0.300 1.365 0.465 ;
        RECT  1.075 0.695 1.365 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.435200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.260 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.170 -0.115 6.440 0.115 ;
        RECT  6.090 -0.115 6.170 0.335 ;
        RECT  5.960 -0.115 6.090 0.115 ;
        RECT  5.880 -0.115 5.960 0.335 ;
        RECT  5.760 -0.115 5.880 0.115 ;
        RECT  5.680 -0.115 5.760 0.335 ;
        RECT  5.570 -0.115 5.680 0.115 ;
        RECT  5.490 -0.115 5.570 0.335 ;
        RECT  5.375 -0.115 5.490 0.115 ;
        RECT  5.295 -0.115 5.375 0.335 ;
        RECT  5.180 -0.115 5.295 0.115 ;
        RECT  5.100 -0.115 5.180 0.335 ;
        RECT  4.980 -0.115 5.100 0.115 ;
        RECT  4.900 -0.115 4.980 0.335 ;
        RECT  4.770 -0.115 4.900 0.115 ;
        RECT  4.690 -0.115 4.770 0.335 ;
        RECT  4.560 -0.115 4.690 0.115 ;
        RECT  4.480 -0.115 4.560 0.335 ;
        RECT  4.350 -0.115 4.480 0.115 ;
        RECT  4.270 -0.115 4.350 0.335 ;
        RECT  4.140 -0.115 4.270 0.115 ;
        RECT  4.060 -0.115 4.140 0.335 ;
        RECT  3.930 -0.115 4.060 0.115 ;
        RECT  3.850 -0.115 3.930 0.335 ;
        RECT  3.730 -0.115 3.850 0.115 ;
        RECT  3.650 -0.115 3.730 0.335 ;
        RECT  3.540 -0.115 3.650 0.115 ;
        RECT  3.460 -0.115 3.540 0.335 ;
        RECT  3.350 -0.115 3.460 0.115 ;
        RECT  3.270 -0.115 3.350 0.335 ;
        RECT  3.165 -0.115 3.270 0.115 ;
        RECT  3.095 -0.115 3.165 0.335 ;
        RECT  2.810 -0.115 3.095 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.300 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.145 6.440 1.375 ;
        RECT  6.090 0.945 6.170 1.375 ;
        RECT  5.960 1.145 6.090 1.375 ;
        RECT  5.880 0.945 5.960 1.375 ;
        RECT  5.760 1.145 5.880 1.375 ;
        RECT  5.680 0.795 5.760 1.375 ;
        RECT  5.570 1.145 5.680 1.375 ;
        RECT  5.490 0.795 5.570 1.375 ;
        RECT  5.375 1.145 5.490 1.375 ;
        RECT  5.295 0.795 5.375 1.375 ;
        RECT  5.180 1.145 5.295 1.375 ;
        RECT  5.100 0.795 5.180 1.375 ;
        RECT  4.980 1.145 5.100 1.375 ;
        RECT  4.900 0.795 4.980 1.375 ;
        RECT  4.770 1.145 4.900 1.375 ;
        RECT  4.690 0.795 4.770 1.375 ;
        RECT  4.560 1.145 4.690 1.375 ;
        RECT  4.480 0.795 4.560 1.375 ;
        RECT  4.350 1.145 4.480 1.375 ;
        RECT  4.270 0.795 4.350 1.375 ;
        RECT  4.140 1.145 4.270 1.375 ;
        RECT  4.060 0.795 4.140 1.375 ;
        RECT  3.930 1.145 4.060 1.375 ;
        RECT  3.850 0.795 3.930 1.375 ;
        RECT  3.730 1.145 3.850 1.375 ;
        RECT  3.650 0.795 3.730 1.375 ;
        RECT  3.540 1.145 3.650 1.375 ;
        RECT  3.460 0.795 3.540 1.375 ;
        RECT  3.350 1.145 3.460 1.375 ;
        RECT  3.270 0.795 3.350 1.375 ;
        RECT  3.170 1.145 3.270 1.375 ;
        RECT  3.090 0.685 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.785 0.185 1.835 0.465 ;
        RECT  1.785 0.695 1.835 1.035 ;
        RECT  1.075 0.300 1.295 0.465 ;
        RECT  1.075 0.695 1.295 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        RECT  6.310 0.210 6.390 0.710 ;
        RECT  6.310 0.790 6.390 1.060 ;
        RECT  6.050 0.630 6.310 0.710 ;
        RECT  5.980 0.790 6.310 0.870 ;
        RECT  5.900 0.430 5.980 0.870 ;
        RECT  3.425 0.430 5.900 0.510 ;
    END
END DCCKND16BWP40

MACRO DCCKND18BWP40
    CLASS CORE ;
    FOREIGN DCCKND18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.918000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.995 0.300 2.145 0.465 ;
        RECT  1.995 0.695 2.145 0.885 ;
        RECT  1.835 0.300 1.995 0.885 ;
        RECT  1.765 0.185 1.835 1.045 ;
        RECT  1.715 0.300 1.765 1.045 ;
        RECT  1.645 0.300 1.715 0.885 ;
        RECT  1.455 0.300 1.645 0.465 ;
        RECT  1.505 0.695 1.645 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.489600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.565 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.010 -0.115 7.280 0.115 ;
        RECT  6.930 -0.115 7.010 0.335 ;
        RECT  6.800 -0.115 6.930 0.115 ;
        RECT  6.720 -0.115 6.800 0.335 ;
        RECT  6.590 -0.115 6.720 0.115 ;
        RECT  6.510 -0.115 6.590 0.335 ;
        RECT  6.390 -0.115 6.510 0.115 ;
        RECT  6.310 -0.115 6.390 0.335 ;
        RECT  6.200 -0.115 6.310 0.115 ;
        RECT  6.120 -0.115 6.200 0.335 ;
        RECT  6.010 -0.115 6.120 0.115 ;
        RECT  5.930 -0.115 6.010 0.335 ;
        RECT  5.815 -0.115 5.930 0.115 ;
        RECT  5.735 -0.115 5.815 0.335 ;
        RECT  5.610 -0.115 5.735 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.190 -0.115 5.320 0.115 ;
        RECT  5.110 -0.115 5.190 0.335 ;
        RECT  4.980 -0.115 5.110 0.115 ;
        RECT  4.900 -0.115 4.980 0.335 ;
        RECT  4.770 -0.115 4.900 0.115 ;
        RECT  4.690 -0.115 4.770 0.335 ;
        RECT  4.560 -0.115 4.690 0.115 ;
        RECT  4.480 -0.115 4.560 0.335 ;
        RECT  4.350 -0.115 4.480 0.115 ;
        RECT  4.270 -0.115 4.350 0.335 ;
        RECT  4.150 -0.115 4.270 0.115 ;
        RECT  4.070 -0.115 4.150 0.335 ;
        RECT  3.960 -0.115 4.070 0.115 ;
        RECT  3.880 -0.115 3.960 0.335 ;
        RECT  3.770 -0.115 3.880 0.115 ;
        RECT  3.690 -0.115 3.770 0.335 ;
        RECT  3.585 -0.115 3.690 0.115 ;
        RECT  3.515 -0.115 3.585 0.330 ;
        RECT  3.190 -0.115 3.515 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.310 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.010 1.145 7.280 1.375 ;
        RECT  6.930 0.945 7.010 1.375 ;
        RECT  6.800 1.145 6.930 1.375 ;
        RECT  6.720 0.945 6.800 1.375 ;
        RECT  6.590 1.145 6.720 1.375 ;
        RECT  6.510 0.795 6.590 1.375 ;
        RECT  6.390 1.145 6.510 1.375 ;
        RECT  6.310 0.795 6.390 1.375 ;
        RECT  6.200 1.145 6.310 1.375 ;
        RECT  6.120 0.795 6.200 1.375 ;
        RECT  6.010 1.145 6.120 1.375 ;
        RECT  5.930 0.795 6.010 1.375 ;
        RECT  5.815 1.145 5.930 1.375 ;
        RECT  5.735 0.795 5.815 1.375 ;
        RECT  5.610 1.145 5.735 1.375 ;
        RECT  5.530 0.795 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.795 5.400 1.375 ;
        RECT  5.190 1.145 5.320 1.375 ;
        RECT  5.110 0.795 5.190 1.375 ;
        RECT  4.980 1.145 5.110 1.375 ;
        RECT  4.900 0.795 4.980 1.375 ;
        RECT  4.770 1.145 4.900 1.375 ;
        RECT  4.690 0.795 4.770 1.375 ;
        RECT  4.560 1.145 4.690 1.375 ;
        RECT  4.480 0.795 4.560 1.375 ;
        RECT  4.350 1.145 4.480 1.375 ;
        RECT  4.270 0.795 4.350 1.375 ;
        RECT  4.150 1.145 4.270 1.375 ;
        RECT  4.070 0.795 4.150 1.375 ;
        RECT  3.960 1.145 4.070 1.375 ;
        RECT  3.880 0.795 3.960 1.375 ;
        RECT  3.770 1.145 3.880 1.375 ;
        RECT  3.690 0.795 3.770 1.375 ;
        RECT  3.590 1.145 3.690 1.375 ;
        RECT  3.510 0.685 3.590 1.375 ;
        RECT  3.190 1.145 3.510 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.645 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.645 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.060 0.695 2.145 0.885 ;
        RECT  1.455 0.300 1.575 0.465 ;
        RECT  1.505 0.695 1.575 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        RECT  7.150 0.210 7.230 0.710 ;
        RECT  7.150 0.790 7.230 1.060 ;
        RECT  6.890 0.630 7.150 0.710 ;
        RECT  6.820 0.790 7.150 0.870 ;
        RECT  6.740 0.430 6.820 0.870 ;
        RECT  3.845 0.430 6.740 0.510 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  2.065 0.300 2.145 0.465 ;
    END
END DCCKND18BWP40

MACRO DCCKND20BWP40
    CLASS CORE ;
    FOREIGN DCCKND20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.047200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.275 0.300 2.525 0.465 ;
        RECT  2.275 0.695 2.525 0.885 ;
        RECT  2.215 0.300 2.275 0.885 ;
        RECT  2.135 0.185 2.215 1.045 ;
        RECT  1.925 0.300 2.135 0.885 ;
        RECT  1.835 0.300 1.925 0.465 ;
        RECT  1.835 0.695 1.925 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.505 0.695 1.765 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.544000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.050 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.850 -0.115 8.120 0.115 ;
        RECT  7.770 -0.115 7.850 0.335 ;
        RECT  7.640 -0.115 7.770 0.115 ;
        RECT  7.560 -0.115 7.640 0.335 ;
        RECT  7.430 -0.115 7.560 0.115 ;
        RECT  7.350 -0.115 7.430 0.335 ;
        RECT  7.220 -0.115 7.350 0.115 ;
        RECT  7.140 -0.115 7.220 0.335 ;
        RECT  7.010 -0.115 7.140 0.115 ;
        RECT  6.930 -0.115 7.010 0.335 ;
        RECT  6.810 -0.115 6.930 0.115 ;
        RECT  6.730 -0.115 6.810 0.335 ;
        RECT  6.620 -0.115 6.730 0.115 ;
        RECT  6.540 -0.115 6.620 0.335 ;
        RECT  6.430 -0.115 6.540 0.115 ;
        RECT  6.350 -0.115 6.430 0.335 ;
        RECT  6.235 -0.115 6.350 0.115 ;
        RECT  6.155 -0.115 6.235 0.335 ;
        RECT  6.030 -0.115 6.155 0.115 ;
        RECT  5.950 -0.115 6.030 0.335 ;
        RECT  5.820 -0.115 5.950 0.115 ;
        RECT  5.740 -0.115 5.820 0.335 ;
        RECT  5.610 -0.115 5.740 0.115 ;
        RECT  5.530 -0.115 5.610 0.335 ;
        RECT  5.400 -0.115 5.530 0.115 ;
        RECT  5.320 -0.115 5.400 0.335 ;
        RECT  5.190 -0.115 5.320 0.115 ;
        RECT  5.110 -0.115 5.190 0.335 ;
        RECT  4.980 -0.115 5.110 0.115 ;
        RECT  4.900 -0.115 4.980 0.335 ;
        RECT  4.770 -0.115 4.900 0.115 ;
        RECT  4.690 -0.115 4.770 0.335 ;
        RECT  4.570 -0.115 4.690 0.115 ;
        RECT  4.490 -0.115 4.570 0.335 ;
        RECT  4.380 -0.115 4.490 0.115 ;
        RECT  4.300 -0.115 4.380 0.335 ;
        RECT  4.190 -0.115 4.300 0.115 ;
        RECT  4.110 -0.115 4.190 0.335 ;
        RECT  4.005 -0.115 4.110 0.115 ;
        RECT  3.935 -0.115 4.005 0.320 ;
        RECT  3.570 -0.115 3.935 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.850 1.145 8.120 1.375 ;
        RECT  7.770 0.945 7.850 1.375 ;
        RECT  7.640 1.145 7.770 1.375 ;
        RECT  7.560 0.945 7.640 1.375 ;
        RECT  7.430 1.145 7.560 1.375 ;
        RECT  7.350 0.795 7.430 1.375 ;
        RECT  7.220 1.145 7.350 1.375 ;
        RECT  7.140 0.795 7.220 1.375 ;
        RECT  7.010 1.145 7.140 1.375 ;
        RECT  6.930 0.795 7.010 1.375 ;
        RECT  6.810 1.145 6.930 1.375 ;
        RECT  6.730 0.795 6.810 1.375 ;
        RECT  6.620 1.145 6.730 1.375 ;
        RECT  6.540 0.795 6.620 1.375 ;
        RECT  6.430 1.145 6.540 1.375 ;
        RECT  6.350 0.795 6.430 1.375 ;
        RECT  6.235 1.145 6.350 1.375 ;
        RECT  6.155 0.795 6.235 1.375 ;
        RECT  6.030 1.145 6.155 1.375 ;
        RECT  5.950 0.795 6.030 1.375 ;
        RECT  5.820 1.145 5.950 1.375 ;
        RECT  5.740 0.795 5.820 1.375 ;
        RECT  5.610 1.145 5.740 1.375 ;
        RECT  5.530 0.795 5.610 1.375 ;
        RECT  5.400 1.145 5.530 1.375 ;
        RECT  5.320 0.795 5.400 1.375 ;
        RECT  5.190 1.145 5.320 1.375 ;
        RECT  5.110 0.795 5.190 1.375 ;
        RECT  4.980 1.145 5.110 1.375 ;
        RECT  4.900 0.795 4.980 1.375 ;
        RECT  4.770 1.145 4.900 1.375 ;
        RECT  4.690 0.795 4.770 1.375 ;
        RECT  4.570 1.145 4.690 1.375 ;
        RECT  4.490 0.795 4.570 1.375 ;
        RECT  4.380 1.145 4.490 1.375 ;
        RECT  4.300 0.795 4.380 1.375 ;
        RECT  4.190 1.145 4.300 1.375 ;
        RECT  4.110 0.795 4.190 1.375 ;
        RECT  4.010 1.145 4.110 1.375 ;
        RECT  3.930 0.685 4.010 1.375 ;
        RECT  3.570 1.145 3.930 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        RECT  7.990 0.210 8.070 0.710 ;
        RECT  7.990 0.790 8.070 1.060 ;
        RECT  7.730 0.630 7.990 0.710 ;
        RECT  7.660 0.790 7.990 0.870 ;
        RECT  7.580 0.430 7.660 0.870 ;
        RECT  4.265 0.430 7.580 0.510 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.345 0.300 2.525 0.465 ;
        RECT  2.345 0.695 2.525 0.885 ;
        RECT  1.835 0.300 1.855 0.465 ;
        RECT  1.835 0.695 1.855 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.505 0.695 1.765 0.885 ;
        RECT  1.385 0.695 1.505 1.045 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.075 0.300 1.385 0.465 ;
    END
END DCCKND20BWP40

MACRO DCCKND24BWP40
    CLASS CORE ;
    FOREIGN DCCKND24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.224000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.555 0.185 2.595 0.465 ;
        RECT  2.555 0.695 2.595 1.035 ;
        RECT  2.525 0.185 2.555 1.035 ;
        RECT  2.215 0.300 2.525 0.885 ;
        RECT  2.205 0.185 2.215 1.045 ;
        RECT  2.135 0.185 2.205 0.465 ;
        RECT  2.135 0.695 2.205 1.045 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.652800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.815 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.250 -0.115 9.520 0.115 ;
        RECT  9.170 -0.115 9.250 0.335 ;
        RECT  9.040 -0.115 9.170 0.115 ;
        RECT  8.960 -0.115 9.040 0.335 ;
        RECT  8.830 -0.115 8.960 0.115 ;
        RECT  8.750 -0.115 8.830 0.335 ;
        RECT  8.620 -0.115 8.750 0.115 ;
        RECT  8.540 -0.115 8.620 0.335 ;
        RECT  8.375 -0.115 8.540 0.115 ;
        RECT  8.295 -0.115 8.375 0.335 ;
        RECT  8.130 -0.115 8.295 0.115 ;
        RECT  8.050 -0.115 8.130 0.335 ;
        RECT  7.920 -0.115 8.050 0.115 ;
        RECT  7.840 -0.115 7.920 0.335 ;
        RECT  7.710 -0.115 7.840 0.115 ;
        RECT  7.630 -0.115 7.710 0.335 ;
        RECT  7.510 -0.115 7.630 0.115 ;
        RECT  7.430 -0.115 7.510 0.335 ;
        RECT  7.320 -0.115 7.430 0.115 ;
        RECT  7.240 -0.115 7.320 0.335 ;
        RECT  7.130 -0.115 7.240 0.115 ;
        RECT  7.050 -0.115 7.130 0.335 ;
        RECT  6.935 -0.115 7.050 0.115 ;
        RECT  6.855 -0.115 6.935 0.335 ;
        RECT  6.730 -0.115 6.855 0.115 ;
        RECT  6.650 -0.115 6.730 0.335 ;
        RECT  6.520 -0.115 6.650 0.115 ;
        RECT  6.440 -0.115 6.520 0.335 ;
        RECT  6.310 -0.115 6.440 0.115 ;
        RECT  6.230 -0.115 6.310 0.335 ;
        RECT  6.100 -0.115 6.230 0.115 ;
        RECT  6.020 -0.115 6.100 0.335 ;
        RECT  5.890 -0.115 6.020 0.115 ;
        RECT  5.810 -0.115 5.890 0.335 ;
        RECT  5.680 -0.115 5.810 0.115 ;
        RECT  5.600 -0.115 5.680 0.335 ;
        RECT  5.470 -0.115 5.600 0.115 ;
        RECT  5.390 -0.115 5.470 0.335 ;
        RECT  5.270 -0.115 5.390 0.115 ;
        RECT  5.190 -0.115 5.270 0.335 ;
        RECT  5.080 -0.115 5.190 0.115 ;
        RECT  5.000 -0.115 5.080 0.335 ;
        RECT  4.890 -0.115 5.000 0.115 ;
        RECT  4.810 -0.115 4.890 0.335 ;
        RECT  4.700 -0.115 4.810 0.115 ;
        RECT  4.600 -0.115 4.700 0.360 ;
        RECT  4.330 -0.115 4.600 0.115 ;
        RECT  4.210 -0.115 4.330 0.230 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.230 ;
        RECT  3.570 -0.115 3.830 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.320 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.250 1.145 9.520 1.375 ;
        RECT  9.170 0.945 9.250 1.375 ;
        RECT  9.040 1.145 9.170 1.375 ;
        RECT  8.960 0.945 9.040 1.375 ;
        RECT  8.830 1.145 8.960 1.375 ;
        RECT  8.750 0.795 8.830 1.375 ;
        RECT  8.620 1.145 8.750 1.375 ;
        RECT  8.540 0.795 8.620 1.375 ;
        RECT  8.375 1.145 8.540 1.375 ;
        RECT  8.295 0.795 8.375 1.375 ;
        RECT  8.130 1.145 8.295 1.375 ;
        RECT  8.050 0.795 8.130 1.375 ;
        RECT  7.920 1.145 8.050 1.375 ;
        RECT  7.840 0.795 7.920 1.375 ;
        RECT  7.710 1.145 7.840 1.375 ;
        RECT  7.630 0.795 7.710 1.375 ;
        RECT  7.510 1.145 7.630 1.375 ;
        RECT  7.430 0.795 7.510 1.375 ;
        RECT  7.320 1.145 7.430 1.375 ;
        RECT  7.240 0.795 7.320 1.375 ;
        RECT  7.130 1.145 7.240 1.375 ;
        RECT  7.050 0.795 7.130 1.375 ;
        RECT  6.935 1.145 7.050 1.375 ;
        RECT  6.855 0.795 6.935 1.375 ;
        RECT  6.730 1.145 6.855 1.375 ;
        RECT  6.650 0.795 6.730 1.375 ;
        RECT  6.520 1.145 6.650 1.375 ;
        RECT  6.440 0.795 6.520 1.375 ;
        RECT  6.310 1.145 6.440 1.375 ;
        RECT  6.230 0.795 6.310 1.375 ;
        RECT  6.100 1.145 6.230 1.375 ;
        RECT  6.020 0.795 6.100 1.375 ;
        RECT  5.890 1.145 6.020 1.375 ;
        RECT  5.810 0.795 5.890 1.375 ;
        RECT  5.680 1.145 5.810 1.375 ;
        RECT  5.600 0.795 5.680 1.375 ;
        RECT  5.470 1.145 5.600 1.375 ;
        RECT  5.390 0.795 5.470 1.375 ;
        RECT  5.270 1.145 5.390 1.375 ;
        RECT  5.190 0.795 5.270 1.375 ;
        RECT  5.080 1.145 5.190 1.375 ;
        RECT  5.000 0.795 5.080 1.375 ;
        RECT  4.890 1.145 5.000 1.375 ;
        RECT  4.810 0.795 4.890 1.375 ;
        RECT  4.700 1.145 4.810 1.375 ;
        RECT  4.600 0.695 4.700 1.375 ;
        RECT  4.330 1.145 4.600 1.375 ;
        RECT  4.210 0.955 4.330 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 0.955 3.950 1.375 ;
        RECT  3.570 1.145 3.830 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.955 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.625 0.300 2.905 0.465 ;
        RECT  2.625 0.695 2.905 0.885 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        RECT  9.390 0.210 9.470 0.710 ;
        RECT  9.390 0.790 9.470 1.060 ;
        RECT  9.130 0.630 9.390 0.710 ;
        RECT  9.060 0.790 9.390 0.870 ;
        RECT  8.980 0.430 9.060 0.870 ;
        RECT  4.965 0.430 8.980 0.510 ;
    END
END DCCKND24BWP40

MACRO DCCKND4BWP40
    CLASS CORE ;
    FOREIGN DCCKND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.201000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.660 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.595 0.705 0.665 0.820 ;
        RECT  0.595 0.310 0.660 0.445 ;
        RECT  0.385 0.310 0.595 0.820 ;
        RECT  0.320 0.310 0.385 0.445 ;
        RECT  0.315 0.705 0.385 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.107200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.675 -0.115 1.960 0.115 ;
        RECT  1.595 -0.115 1.675 0.330 ;
        RECT  1.375 -0.115 1.595 0.115 ;
        RECT  1.295 -0.115 1.375 0.330 ;
        RECT  1.130 -0.115 1.295 0.115 ;
        RECT  1.050 -0.115 1.130 0.330 ;
        RECT  0.930 -0.115 1.050 0.115 ;
        RECT  0.850 -0.115 0.930 0.335 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.145 1.960 1.375 ;
        RECT  1.590 0.955 1.670 1.375 ;
        RECT  1.380 1.145 1.590 1.375 ;
        RECT  1.300 0.955 1.380 1.375 ;
        RECT  1.130 1.145 1.300 1.375 ;
        RECT  1.050 0.805 1.130 1.375 ;
        RECT  0.930 1.145 1.050 1.375 ;
        RECT  0.850 0.695 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        RECT  1.815 0.210 1.895 0.710 ;
        RECT  1.815 0.790 1.895 1.050 ;
        RECT  1.580 0.630 1.815 0.710 ;
        RECT  1.510 0.790 1.815 0.870 ;
        RECT  1.430 0.430 1.510 0.870 ;
        RECT  1.215 0.430 1.430 0.510 ;
    END
END DCCKND4BWP40

MACRO DCCKND5BWP40
    CLASS CORE ;
    FOREIGN DCCKND5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.304850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.735 0.705 1.105 0.820 ;
        RECT  0.740 0.310 1.100 0.445 ;
        RECT  0.735 0.185 0.740 0.445 ;
        RECT  0.665 0.185 0.735 1.030 ;
        RECT  0.660 0.185 0.665 0.820 ;
        RECT  0.525 0.310 0.660 0.820 ;
        RECT  0.320 0.310 0.525 0.445 ;
        RECT  0.315 0.705 0.525 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.134000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.445 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.250 0.335 ;
        RECT  2.040 -0.115 2.170 0.115 ;
        RECT  1.960 -0.115 2.040 0.335 ;
        RECT  1.810 -0.115 1.960 0.115 ;
        RECT  1.730 -0.115 1.810 0.335 ;
        RECT  1.580 -0.115 1.730 0.115 ;
        RECT  1.500 -0.115 1.580 0.335 ;
        RECT  1.390 -0.115 1.500 0.115 ;
        RECT  1.310 -0.115 1.390 0.335 ;
        RECT  0.980 -0.115 1.310 0.115 ;
        RECT  0.860 -0.115 0.980 0.240 ;
        RECT  0.560 -0.115 0.860 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.145 2.520 1.375 ;
        RECT  2.170 0.945 2.250 1.375 ;
        RECT  2.040 1.145 2.170 1.375 ;
        RECT  1.960 0.945 2.040 1.375 ;
        RECT  1.810 1.145 1.960 1.375 ;
        RECT  1.730 0.795 1.810 1.375 ;
        RECT  1.580 1.145 1.730 1.375 ;
        RECT  1.500 0.795 1.580 1.375 ;
        RECT  1.390 1.145 1.500 1.375 ;
        RECT  1.310 0.795 1.390 1.375 ;
        RECT  0.970 1.145 1.310 1.375 ;
        RECT  0.850 0.890 0.970 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.805 0.705 1.105 0.820 ;
        RECT  0.805 0.310 1.100 0.445 ;
        RECT  0.320 0.310 0.455 0.445 ;
        RECT  0.315 0.705 0.455 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        RECT  2.390 0.210 2.470 0.710 ;
        RECT  2.390 0.790 2.470 1.060 ;
        RECT  2.130 0.630 2.390 0.710 ;
        RECT  2.060 0.790 2.390 0.870 ;
        RECT  1.980 0.430 2.060 0.870 ;
        RECT  1.465 0.430 1.980 0.510 ;
    END
END DCCKND5BWP40

MACRO DCCKND6BWP40
    CLASS CORE ;
    FOREIGN DCCKND6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.301500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.875 0.705 1.045 0.820 ;
        RECT  0.875 0.310 1.040 0.445 ;
        RECT  0.740 0.310 0.875 0.820 ;
        RECT  0.735 0.185 0.740 0.820 ;
        RECT  0.665 0.185 0.735 1.030 ;
        RECT  0.660 0.185 0.665 0.445 ;
        RECT  0.315 0.705 0.665 0.820 ;
        RECT  0.320 0.310 0.660 0.445 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.160800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.515 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.115 2.800 0.115 ;
        RECT  2.450 -0.115 2.530 0.335 ;
        RECT  2.320 -0.115 2.450 0.115 ;
        RECT  2.240 -0.115 2.320 0.335 ;
        RECT  2.110 -0.115 2.240 0.115 ;
        RECT  2.030 -0.115 2.110 0.335 ;
        RECT  1.910 -0.115 2.030 0.115 ;
        RECT  1.830 -0.115 1.910 0.335 ;
        RECT  1.720 -0.115 1.830 0.115 ;
        RECT  1.640 -0.115 1.720 0.335 ;
        RECT  1.530 -0.115 1.640 0.115 ;
        RECT  1.450 -0.115 1.530 0.335 ;
        RECT  1.330 -0.115 1.450 0.115 ;
        RECT  1.210 -0.115 1.330 0.240 ;
        RECT  0.950 -0.115 1.210 0.115 ;
        RECT  0.830 -0.115 0.950 0.240 ;
        RECT  0.560 -0.115 0.830 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.320 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.145 2.800 1.375 ;
        RECT  2.450 0.945 2.530 1.375 ;
        RECT  2.320 1.145 2.450 1.375 ;
        RECT  2.240 0.945 2.320 1.375 ;
        RECT  2.110 1.145 2.240 1.375 ;
        RECT  2.030 0.795 2.110 1.375 ;
        RECT  1.910 1.145 2.030 1.375 ;
        RECT  1.830 0.795 1.910 1.375 ;
        RECT  1.720 1.145 1.830 1.375 ;
        RECT  1.640 0.795 1.720 1.375 ;
        RECT  1.530 1.145 1.640 1.375 ;
        RECT  1.450 0.795 1.530 1.375 ;
        RECT  1.330 1.145 1.450 1.375 ;
        RECT  1.210 0.750 1.330 1.375 ;
        RECT  0.960 1.145 1.210 1.375 ;
        RECT  0.830 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.830 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.945 0.705 1.045 0.820 ;
        RECT  0.945 0.310 1.040 0.445 ;
        RECT  0.320 0.310 0.595 0.445 ;
        RECT  0.315 0.705 0.595 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        RECT  2.670 0.210 2.750 0.710 ;
        RECT  2.670 0.790 2.750 1.060 ;
        RECT  2.410 0.630 2.670 0.710 ;
        RECT  2.340 0.790 2.670 0.870 ;
        RECT  2.260 0.430 2.340 0.870 ;
        RECT  1.605 0.430 2.260 0.510 ;
    END
END DCCKND6BWP40

MACRO DCCKND8BWP40
    CLASS CORE ;
    FOREIGN DCCKND8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.431800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.015 0.185 1.095 0.445 ;
        RECT  1.020 0.705 1.090 1.030 ;
        RECT  1.015 0.705 1.020 0.820 ;
        RECT  0.700 0.310 1.015 0.820 ;
        RECT  0.695 0.185 0.700 0.820 ;
        RECT  0.665 0.185 0.695 1.030 ;
        RECT  0.620 0.185 0.665 0.445 ;
        RECT  0.625 0.705 0.665 1.030 ;
        RECT  0.315 0.705 0.625 0.820 ;
        RECT  0.320 0.310 0.620 0.445 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.217600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 -0.115 3.640 0.115 ;
        RECT  3.290 -0.115 3.370 0.335 ;
        RECT  3.160 -0.115 3.290 0.115 ;
        RECT  3.080 -0.115 3.160 0.335 ;
        RECT  2.950 -0.115 3.080 0.115 ;
        RECT  2.870 -0.115 2.950 0.335 ;
        RECT  2.740 -0.115 2.870 0.115 ;
        RECT  2.660 -0.115 2.740 0.335 ;
        RECT  2.530 -0.115 2.660 0.115 ;
        RECT  2.450 -0.115 2.530 0.335 ;
        RECT  2.330 -0.115 2.450 0.115 ;
        RECT  2.250 -0.115 2.330 0.335 ;
        RECT  2.140 -0.115 2.250 0.115 ;
        RECT  2.060 -0.115 2.140 0.335 ;
        RECT  1.950 -0.115 2.060 0.115 ;
        RECT  1.870 -0.115 1.950 0.335 ;
        RECT  1.750 -0.115 1.870 0.115 ;
        RECT  1.665 -0.115 1.750 0.345 ;
        RECT  1.305 -0.115 1.665 0.115 ;
        RECT  1.185 -0.115 1.305 0.240 ;
        RECT  0.910 -0.115 1.185 0.115 ;
        RECT  0.790 -0.115 0.910 0.240 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.240 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.145 3.640 1.375 ;
        RECT  3.290 0.945 3.370 1.375 ;
        RECT  3.160 1.145 3.290 1.375 ;
        RECT  3.080 0.945 3.160 1.375 ;
        RECT  2.950 1.145 3.080 1.375 ;
        RECT  2.870 0.795 2.950 1.375 ;
        RECT  2.740 1.145 2.870 1.375 ;
        RECT  2.660 0.795 2.740 1.375 ;
        RECT  2.530 1.145 2.660 1.375 ;
        RECT  2.450 0.795 2.530 1.375 ;
        RECT  2.330 1.145 2.450 1.375 ;
        RECT  2.250 0.795 2.330 1.375 ;
        RECT  2.140 1.145 2.250 1.375 ;
        RECT  2.060 0.795 2.140 1.375 ;
        RECT  1.950 1.145 2.060 1.375 ;
        RECT  1.870 0.795 1.950 1.375 ;
        RECT  1.780 1.145 1.870 1.375 ;
        RECT  1.670 0.725 1.780 1.375 ;
        RECT  1.310 1.145 1.670 1.375 ;
        RECT  1.190 0.890 1.310 1.375 ;
        RECT  0.915 1.145 1.190 1.375 ;
        RECT  0.795 0.890 0.915 1.375 ;
        RECT  0.530 1.145 0.795 1.375 ;
        RECT  0.410 0.890 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.085 0.185 1.095 0.445 ;
        RECT  1.085 0.705 1.090 1.030 ;
        RECT  0.320 0.310 0.595 0.445 ;
        RECT  0.315 0.705 0.595 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        RECT  3.510 0.210 3.590 0.710 ;
        RECT  3.510 0.790 3.590 1.060 ;
        RECT  3.250 0.630 3.510 0.710 ;
        RECT  3.180 0.790 3.510 0.870 ;
        RECT  3.100 0.430 3.180 0.870 ;
        RECT  2.025 0.430 3.100 0.510 ;
    END
END DCCKND8BWP40

MACRO DELAD1BWP40
    CLASS CORE ;
    FOREIGN DELAD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.195 1.225 1.070 ;
        RECT  1.120 0.195 1.155 0.315 ;
        RECT  1.120 0.970 1.155 1.070 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 -0.115 1.260 0.115 ;
        RECT  0.900 -0.115 1.020 0.230 ;
        RECT  0.360 -0.115 0.900 0.115 ;
        RECT  0.240 -0.115 0.360 0.230 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.145 1.260 1.375 ;
        RECT  0.900 1.030 1.020 1.375 ;
        RECT  0.360 1.145 0.900 1.375 ;
        RECT  0.240 1.030 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.010 0.385 1.080 0.855 ;
        RECT  0.805 0.385 1.010 0.455 ;
        RECT  0.800 0.785 1.010 0.855 ;
        RECT  0.605 0.535 0.895 0.640 ;
        RECT  0.695 0.195 0.805 0.455 ;
        RECT  0.695 0.785 0.800 1.060 ;
        RECT  0.535 0.200 0.605 1.045 ;
        RECT  0.455 0.200 0.535 0.270 ;
        RECT  0.455 0.975 0.535 1.045 ;
        RECT  0.345 0.520 0.465 0.640 ;
        RECT  0.275 0.325 0.345 0.935 ;
        RECT  0.145 0.325 0.275 0.395 ;
        RECT  0.145 0.865 0.275 0.935 ;
        RECT  0.035 0.195 0.145 0.395 ;
        RECT  0.035 0.865 0.145 1.060 ;
    END
END DELAD1BWP40

MACRO DELBD1BWP40
    CLASS CORE ;
    FOREIGN DELBD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.096000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.195 1.645 1.065 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 -0.115 1.680 0.115 ;
        RECT  1.365 -0.115 1.435 0.425 ;
        RECT  0.360 -0.115 1.365 0.115 ;
        RECT  0.240 -0.115 0.360 0.250 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 1.145 1.680 1.375 ;
        RECT  1.365 0.790 1.435 1.375 ;
        RECT  0.360 1.145 1.365 1.375 ;
        RECT  0.240 1.010 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.520 1.485 0.640 ;
        RECT  1.225 0.195 1.295 1.065 ;
        RECT  0.940 0.195 1.225 0.265 ;
        RECT  0.940 0.995 1.225 1.065 ;
        RECT  1.055 0.345 1.155 0.915 ;
        RECT  0.860 0.195 0.940 0.315 ;
        RECT  0.860 0.925 0.940 1.065 ;
        RECT  0.745 0.525 0.930 0.640 ;
        RECT  0.675 0.195 0.745 1.055 ;
        RECT  0.535 0.220 0.605 1.030 ;
        RECT  0.455 0.220 0.535 0.290 ;
        RECT  0.455 0.960 0.535 1.030 ;
        RECT  0.345 0.520 0.465 0.640 ;
        RECT  0.275 0.345 0.345 0.915 ;
        RECT  0.145 0.345 0.275 0.415 ;
        RECT  0.145 0.845 0.275 0.915 ;
        RECT  0.035 0.185 0.145 0.415 ;
        RECT  0.035 0.845 0.145 1.075 ;
    END
END DELBD1BWP40

MACRO DELCD1BWP40
    CLASS CORE ;
    FOREIGN DELCD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.116000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 0.185 2.065 1.075 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.015800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.830 -0.115 2.100 0.115 ;
        RECT  1.730 -0.115 1.830 0.415 ;
        RECT  0.360 -0.115 1.730 0.115 ;
        RECT  0.240 -0.115 0.360 0.250 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.145 2.100 1.375 ;
        RECT  1.730 0.745 1.830 1.375 ;
        RECT  0.360 1.145 1.730 1.375 ;
        RECT  0.240 1.010 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.650 0.520 1.880 0.640 ;
        RECT  1.580 0.195 1.650 1.065 ;
        RECT  1.120 0.195 1.580 0.265 ;
        RECT  1.120 0.995 1.580 1.065 ;
        RECT  1.410 0.345 1.510 0.915 ;
        RECT  1.220 0.345 1.320 0.915 ;
        RECT  0.965 0.555 1.140 0.670 ;
        RECT  1.040 0.195 1.120 0.420 ;
        RECT  1.040 0.895 1.120 1.065 ;
        RECT  0.895 0.230 0.965 1.035 ;
        RECT  0.815 0.230 0.895 0.300 ;
        RECT  0.815 0.965 0.895 1.035 ;
        RECT  0.675 0.205 0.745 1.060 ;
        RECT  0.535 0.230 0.605 1.035 ;
        RECT  0.455 0.230 0.535 0.300 ;
        RECT  0.455 0.965 0.535 1.035 ;
        RECT  0.345 0.550 0.465 0.670 ;
        RECT  0.275 0.345 0.345 0.940 ;
        RECT  0.140 0.345 0.275 0.415 ;
        RECT  0.145 0.870 0.275 0.940 ;
        RECT  0.035 0.870 0.145 1.045 ;
        RECT  0.050 0.200 0.140 0.415 ;
    END
END DELCD1BWP40

MACRO DELDD1BWP40
    CLASS CORE ;
    FOREIGN DELDD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.095000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.195 2.905 1.045 ;
        RECT  2.810 0.195 2.825 0.455 ;
        RECT  2.810 0.755 2.825 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.940 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.940 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.650 0.520 2.755 0.640 ;
        RECT  2.580 0.195 2.650 1.065 ;
        RECT  2.290 0.195 2.580 0.265 ;
        RECT  2.290 0.995 2.580 1.065 ;
        RECT  2.400 0.345 2.500 0.915 ;
        RECT  2.120 0.565 2.320 0.655 ;
        RECT  2.220 0.195 2.290 0.455 ;
        RECT  2.220 0.805 2.290 1.065 ;
        RECT  2.040 0.335 2.120 0.925 ;
        RECT  1.840 0.335 1.920 0.925 ;
        RECT  1.680 0.335 1.750 0.925 ;
        RECT  1.640 0.335 1.680 0.460 ;
        RECT  1.640 0.790 1.680 0.925 ;
        RECT  1.450 0.550 1.575 0.670 ;
        RECT  1.380 0.195 1.450 1.065 ;
        RECT  0.900 0.195 1.380 0.265 ;
        RECT  0.900 0.995 1.380 1.065 ;
        RECT  1.210 0.345 1.310 0.915 ;
        RECT  1.010 0.345 1.110 0.915 ;
        RECT  0.720 0.560 0.925 0.660 ;
        RECT  0.830 0.195 0.900 0.455 ;
        RECT  0.830 0.805 0.900 1.065 ;
        RECT  0.650 0.320 0.720 0.940 ;
        RECT  0.510 0.320 0.580 0.940 ;
        RECT  0.445 0.320 0.510 0.440 ;
        RECT  0.445 0.820 0.510 0.940 ;
        RECT  0.345 0.520 0.440 0.640 ;
        RECT  0.275 0.345 0.345 0.915 ;
        RECT  0.035 0.345 0.275 0.415 ;
        RECT  0.035 0.845 0.275 0.915 ;
    END
END DELDD1BWP40

MACRO DELED1BWP40
    CLASS CORE ;
    FOREIGN DELED1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.095000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.200 3.185 1.045 ;
        RECT  3.090 0.200 3.105 0.455 ;
        RECT  3.090 0.770 3.105 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 3.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.940 0.520 3.035 0.640 ;
        RECT  2.870 0.195 2.940 1.065 ;
        RECT  2.390 0.195 2.870 0.265 ;
        RECT  2.390 0.995 2.870 1.065 ;
        RECT  2.690 0.345 2.790 0.915 ;
        RECT  2.500 0.345 2.600 0.915 ;
        RECT  2.320 0.195 2.390 0.455 ;
        RECT  2.320 0.805 2.390 1.065 ;
        RECT  2.220 0.565 2.365 0.655 ;
        RECT  2.140 0.335 2.220 0.925 ;
        RECT  1.950 0.335 2.030 0.925 ;
        RECT  1.785 0.335 1.855 0.925 ;
        RECT  1.730 0.335 1.785 0.455 ;
        RECT  1.730 0.805 1.785 0.925 ;
        RECT  1.620 0.550 1.715 0.670 ;
        RECT  1.550 0.195 1.620 1.065 ;
        RECT  1.080 0.195 1.550 0.265 ;
        RECT  1.080 0.995 1.550 1.065 ;
        RECT  1.370 0.345 1.470 0.915 ;
        RECT  1.180 0.345 1.280 0.915 ;
        RECT  1.010 0.195 1.080 0.455 ;
        RECT  0.930 0.560 1.080 0.660 ;
        RECT  1.010 0.805 1.080 1.065 ;
        RECT  0.860 0.320 0.930 0.940 ;
        RECT  0.795 0.320 0.860 0.440 ;
        RECT  0.795 0.820 0.860 0.940 ;
        RECT  0.640 0.320 0.710 0.940 ;
        RECT  0.500 0.320 0.570 0.940 ;
        RECT  0.435 0.320 0.500 0.440 ;
        RECT  0.435 0.820 0.500 0.940 ;
        RECT  0.345 0.520 0.430 0.640 ;
        RECT  0.275 0.345 0.345 0.915 ;
        RECT  0.035 0.345 0.275 0.415 ;
        RECT  0.035 0.845 0.275 0.915 ;
    END
END DELED1BWP40

MACRO DELFD1BWP40
    CLASS CORE ;
    FOREIGN DELFD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.095000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.085 0.195 4.165 1.045 ;
        RECT  4.070 0.195 4.085 0.455 ;
        RECT  4.070 0.755 4.085 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.015200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 4.200 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.890 0.520 4.015 0.640 ;
        RECT  3.820 0.195 3.890 1.065 ;
        RECT  3.530 0.195 3.820 0.265 ;
        RECT  3.530 0.995 3.820 1.065 ;
        RECT  3.640 0.345 3.740 0.915 ;
        RECT  3.460 0.195 3.530 0.455 ;
        RECT  3.460 0.805 3.530 1.065 ;
        RECT  3.360 0.565 3.505 0.655 ;
        RECT  3.280 0.335 3.360 0.925 ;
        RECT  3.090 0.335 3.170 0.925 ;
        RECT  2.925 0.335 2.995 0.925 ;
        RECT  2.870 0.335 2.925 0.455 ;
        RECT  2.870 0.805 2.925 0.925 ;
        RECT  2.760 0.550 2.855 0.670 ;
        RECT  2.690 0.195 2.760 1.065 ;
        RECT  2.220 0.195 2.690 0.265 ;
        RECT  2.220 0.995 2.690 1.065 ;
        RECT  2.510 0.345 2.610 0.915 ;
        RECT  2.320 0.345 2.420 0.915 ;
        RECT  2.030 0.565 2.240 0.655 ;
        RECT  2.150 0.195 2.220 0.455 ;
        RECT  2.150 0.805 2.220 1.065 ;
        RECT  1.950 0.335 2.030 0.925 ;
        RECT  1.760 0.335 1.840 0.925 ;
        RECT  1.595 0.335 1.665 0.925 ;
        RECT  1.540 0.335 1.595 0.455 ;
        RECT  1.540 0.805 1.595 0.925 ;
        RECT  1.430 0.550 1.525 0.670 ;
        RECT  1.360 0.195 1.430 1.065 ;
        RECT  0.890 0.195 1.360 0.265 ;
        RECT  0.890 0.995 1.360 1.065 ;
        RECT  1.180 0.345 1.280 0.915 ;
        RECT  0.990 0.345 1.090 0.915 ;
        RECT  0.820 0.195 0.890 0.455 ;
        RECT  0.740 0.560 0.890 0.660 ;
        RECT  0.820 0.805 0.890 1.065 ;
        RECT  0.670 0.320 0.740 0.940 ;
        RECT  0.640 0.320 0.670 0.440 ;
        RECT  0.640 0.820 0.670 0.940 ;
        RECT  0.500 0.320 0.570 0.940 ;
        RECT  0.435 0.320 0.500 0.440 ;
        RECT  0.435 0.820 0.500 0.940 ;
        RECT  0.345 0.520 0.430 0.640 ;
        RECT  0.275 0.345 0.345 0.915 ;
        RECT  0.035 0.345 0.275 0.415 ;
        RECT  0.035 0.845 0.275 0.915 ;
    END
END DELFD1BWP40

MACRO DELGD1BWP40
    CLASS CORE ;
    FOREIGN DELGD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.095000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.505 0.195 4.585 1.045 ;
        RECT  4.490 0.195 4.505 0.455 ;
        RECT  4.490 0.760 4.505 1.045 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.520 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.620 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 4.620 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.310 0.520 4.435 0.640 ;
        RECT  4.240 0.195 4.310 1.065 ;
        RECT  3.945 0.195 4.240 0.265 ;
        RECT  3.945 0.995 4.240 1.065 ;
        RECT  4.060 0.345 4.160 0.915 ;
        RECT  3.865 0.195 3.945 0.455 ;
        RECT  3.865 0.805 3.945 1.065 ;
        RECT  3.725 0.335 3.795 0.925 ;
        RECT  3.640 0.335 3.725 0.455 ;
        RECT  3.640 0.805 3.725 0.925 ;
        RECT  3.540 0.550 3.655 0.670 ;
        RECT  3.460 0.335 3.540 0.925 ;
        RECT  3.270 0.335 3.350 0.925 ;
        RECT  3.105 0.335 3.175 0.925 ;
        RECT  3.050 0.335 3.105 0.455 ;
        RECT  3.050 0.805 3.105 0.925 ;
        RECT  2.940 0.550 3.035 0.670 ;
        RECT  2.870 0.195 2.940 1.065 ;
        RECT  2.400 0.195 2.870 0.265 ;
        RECT  2.400 0.995 2.870 1.065 ;
        RECT  2.690 0.345 2.790 0.915 ;
        RECT  2.500 0.345 2.600 0.915 ;
        RECT  2.220 0.565 2.420 0.655 ;
        RECT  2.330 0.195 2.400 0.455 ;
        RECT  2.330 0.805 2.400 1.065 ;
        RECT  2.140 0.335 2.220 0.925 ;
        RECT  1.950 0.335 2.030 0.925 ;
        RECT  1.785 0.335 1.855 0.925 ;
        RECT  1.730 0.335 1.785 0.455 ;
        RECT  1.730 0.805 1.785 0.925 ;
        RECT  1.620 0.550 1.715 0.670 ;
        RECT  1.550 0.195 1.620 1.065 ;
        RECT  1.080 0.195 1.550 0.265 ;
        RECT  1.080 0.995 1.550 1.065 ;
        RECT  1.370 0.345 1.470 0.915 ;
        RECT  1.180 0.345 1.280 0.915 ;
        RECT  1.010 0.195 1.080 0.455 ;
        RECT  0.930 0.560 1.080 0.660 ;
        RECT  1.010 0.805 1.080 1.065 ;
        RECT  0.860 0.320 0.930 0.940 ;
        RECT  0.830 0.320 0.860 0.440 ;
        RECT  0.830 0.820 0.860 0.940 ;
        RECT  0.640 0.320 0.710 0.940 ;
        RECT  0.500 0.320 0.570 0.940 ;
        RECT  0.435 0.320 0.500 0.440 ;
        RECT  0.435 0.820 0.500 0.940 ;
        RECT  0.345 0.520 0.430 0.640 ;
        RECT  0.275 0.345 0.345 0.915 ;
        RECT  0.035 0.345 0.275 0.415 ;
        RECT  0.035 0.845 0.275 0.915 ;
    END
END DELGD1BWP40

MACRO DFCNQD0BWP40
    CLASS CORE ;
    FOREIGN DFCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 1.075 ;
        RECT  3.795 0.185 3.815 0.310 ;
        RECT  3.795 0.905 3.815 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.550 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 -0.115 3.920 0.115 ;
        RECT  3.580 -0.115 3.700 0.235 ;
        RECT  3.100 -0.115 3.580 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.235 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 0.995 3.290 1.375 ;
        RECT  3.115 1.145 3.200 1.375 ;
        RECT  3.015 0.875 3.115 1.375 ;
        RECT  2.335 1.145 3.015 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.925 ;
        RECT  3.185 0.325 3.655 0.395 ;
        RECT  3.480 0.855 3.655 0.925 ;
        RECT  3.390 0.855 3.480 1.025 ;
        RECT  3.300 0.855 3.390 0.925 ;
        RECT  3.230 0.720 3.300 0.925 ;
        RECT  2.705 0.540 3.295 0.610 ;
        RECT  3.005 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.705 0.610 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.810 ;
        RECT  2.010 0.335 2.070 0.810 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.010 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.215 0.625 0.945 ;
        RECT  0.415 0.215 0.555 0.285 ;
        RECT  0.520 0.875 0.555 0.945 ;
        RECT  0.420 0.875 0.520 1.055 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.150 0.345 0.275 0.415 ;
        RECT  0.130 0.840 0.275 0.910 ;
        RECT  0.055 0.195 0.150 0.415 ;
        RECT  0.055 0.840 0.130 1.055 ;
    END
END DFCNQD0BWP40

MACRO DFCNQD1BWP40
    CLASS CORE ;
    FOREIGN DFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.185 3.885 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.024400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.550 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 -0.115 3.920 0.115 ;
        RECT  3.570 -0.115 3.700 0.235 ;
        RECT  3.100 -0.115 3.570 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 0.995 3.290 1.375 ;
        RECT  3.120 1.145 3.200 1.375 ;
        RECT  3.010 0.885 3.120 1.375 ;
        RECT  2.335 1.145 3.010 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.925 ;
        RECT  3.185 0.325 3.655 0.395 ;
        RECT  3.300 0.855 3.655 0.925 ;
        RECT  3.230 0.720 3.300 0.925 ;
        RECT  2.705 0.540 3.295 0.610 ;
        RECT  3.005 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.705 0.610 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.810 ;
        RECT  2.060 0.335 2.070 0.810 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.060 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQD1BWP40

MACRO DFCNQD2BWP40
    CLASS CORE ;
    FOREIGN DFCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.024400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.550 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 -0.115 4.200 0.115 ;
        RECT  4.060 -0.115 4.130 0.480 ;
        RECT  3.700 -0.115 4.060 0.115 ;
        RECT  3.575 -0.115 3.700 0.235 ;
        RECT  3.100 -0.115 3.575 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.130 1.145 4.200 1.375 ;
        RECT  4.060 0.725 4.130 1.375 ;
        RECT  3.690 1.145 4.060 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 0.995 3.290 1.375 ;
        RECT  3.125 1.145 3.200 1.375 ;
        RECT  3.005 0.900 3.125 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.925 ;
        RECT  3.185 0.325 3.655 0.395 ;
        RECT  3.300 0.855 3.655 0.925 ;
        RECT  3.230 0.720 3.300 0.925 ;
        RECT  2.705 0.540 3.295 0.610 ;
        RECT  2.920 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.705 0.610 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.810 ;
        RECT  2.015 0.335 2.070 0.810 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.015 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQD2BWP40

MACRO DFCNQD4BWP40
    CLASS CORE ;
    FOREIGN DFCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.264900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.745 4.880 1.000 ;
        RECT  4.795 0.205 4.870 0.485 ;
        RECT  4.785 0.205 4.795 1.000 ;
        RECT  4.770 0.355 4.785 1.000 ;
        RECT  4.585 0.355 4.770 0.830 ;
        RECT  4.480 0.355 4.585 0.485 ;
        RECT  4.480 0.710 4.585 0.830 ;
        RECT  4.400 0.205 4.480 0.485 ;
        RECT  4.400 0.710 4.480 1.000 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.024400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.050600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.875 0.625 4.055 0.765 ;
        RECT  3.675 0.570 3.875 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 -0.115 5.180 0.115 ;
        RECT  5.040 -0.115 5.110 0.480 ;
        RECT  4.665 -0.115 5.040 0.115 ;
        RECT  4.590 -0.115 4.665 0.275 ;
        RECT  4.275 -0.115 4.590 0.115 ;
        RECT  4.205 -0.115 4.275 0.190 ;
        RECT  3.910 -0.115 4.205 0.115 ;
        RECT  3.775 -0.115 3.910 0.210 ;
        RECT  3.100 -0.115 3.775 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.145 5.180 1.375 ;
        RECT  5.040 0.725 5.110 1.375 ;
        RECT  4.660 1.145 5.040 1.375 ;
        RECT  4.590 0.960 4.660 1.375 ;
        RECT  4.280 1.145 4.590 1.375 ;
        RECT  4.205 1.000 4.280 1.375 ;
        RECT  3.690 1.145 4.205 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 0.995 3.290 1.375 ;
        RECT  3.120 1.145 3.200 1.375 ;
        RECT  3.005 0.895 3.120 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.745 4.880 1.000 ;
        RECT  4.865 0.205 4.870 0.485 ;
        RECT  4.480 0.355 4.515 0.485 ;
        RECT  4.480 0.710 4.515 0.830 ;
        RECT  4.400 0.205 4.480 0.485 ;
        RECT  4.400 0.710 4.480 1.000 ;
        RECT  4.255 0.280 4.330 0.925 ;
        RECT  3.380 0.280 4.255 0.350 ;
        RECT  3.300 0.855 4.255 0.925 ;
        RECT  3.280 0.430 4.090 0.500 ;
        RECT  2.705 0.570 3.495 0.640 ;
        RECT  3.230 0.720 3.300 0.925 ;
        RECT  3.210 0.335 3.280 0.500 ;
        RECT  2.920 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.705 0.640 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.810 ;
        RECT  2.015 0.335 2.070 0.810 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.015 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQD4BWP40

MACRO DFCNQND0BWP40
    CLASS CORE ;
    FOREIGN DFCNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.300 4.025 1.055 ;
        RECT  3.935 0.300 3.955 0.465 ;
        RECT  3.935 0.900 3.955 1.055 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.690 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.810 -0.115 4.060 0.115 ;
        RECT  3.690 -0.115 3.810 0.145 ;
        RECT  3.095 -0.115 3.690 0.115 ;
        RECT  3.005 -0.115 3.095 0.420 ;
        RECT  2.210 -0.115 3.005 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.805 1.145 4.060 1.375 ;
        RECT  3.735 0.940 3.805 1.375 ;
        RECT  3.415 1.145 3.735 1.375 ;
        RECT  3.325 1.095 3.415 1.375 ;
        RECT  3.215 1.145 3.325 1.375 ;
        RECT  3.145 1.095 3.215 1.375 ;
        RECT  2.335 1.145 3.145 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.865 0.605 3.870 0.740 ;
        RECT  3.790 0.220 3.865 0.740 ;
        RECT  3.235 0.220 3.790 0.295 ;
        RECT  3.455 0.925 3.620 1.000 ;
        RECT  3.385 0.375 3.455 1.000 ;
        RECT  3.310 0.375 3.385 0.445 ;
        RECT  3.055 0.630 3.385 0.700 ;
        RECT  3.200 0.815 3.300 0.915 ;
        RECT  3.165 0.220 3.235 0.560 ;
        RECT  2.655 0.845 3.200 0.915 ;
        RECT  2.975 0.490 3.165 0.560 ;
        RECT  2.905 0.490 2.975 0.775 ;
        RECT  2.880 0.490 2.905 0.560 ;
        RECT  2.770 0.995 2.895 1.075 ;
        RECT  2.810 0.315 2.880 0.560 ;
        RECT  2.485 0.995 2.770 1.065 ;
        RECT  2.585 0.335 2.655 0.915 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.810 ;
        RECT  2.015 0.335 2.070 0.810 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.015 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQND0BWP40

MACRO DFCNQND1BWP40
    CLASS CORE ;
    FOREIGN DFCNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.093600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.185 4.025 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.690 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.810 -0.115 4.060 0.115 ;
        RECT  3.690 -0.115 3.810 0.145 ;
        RECT  3.095 -0.115 3.690 0.115 ;
        RECT  3.000 -0.115 3.095 0.425 ;
        RECT  2.210 -0.115 3.000 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.830 1.145 4.060 1.375 ;
        RECT  3.710 0.885 3.830 1.375 ;
        RECT  3.415 1.145 3.710 1.375 ;
        RECT  3.325 1.095 3.415 1.375 ;
        RECT  3.230 1.145 3.325 1.375 ;
        RECT  3.130 0.985 3.230 1.375 ;
        RECT  2.335 1.145 3.130 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.790 0.220 3.865 0.660 ;
        RECT  3.235 0.220 3.790 0.295 ;
        RECT  3.455 0.925 3.620 1.000 ;
        RECT  3.385 0.375 3.455 1.000 ;
        RECT  3.310 0.375 3.385 0.445 ;
        RECT  3.055 0.635 3.385 0.705 ;
        RECT  3.200 0.815 3.300 0.915 ;
        RECT  3.165 0.220 3.235 0.565 ;
        RECT  2.655 0.845 3.200 0.915 ;
        RECT  2.975 0.495 3.165 0.565 ;
        RECT  2.905 0.495 2.975 0.775 ;
        RECT  2.880 0.495 2.905 0.565 ;
        RECT  2.770 0.995 2.895 1.075 ;
        RECT  2.810 0.315 2.880 0.565 ;
        RECT  2.485 0.995 2.770 1.065 ;
        RECT  2.585 0.335 2.655 0.915 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.135 0.820 ;
        RECT  2.015 0.335 2.070 0.820 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.015 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQND1BWP40

MACRO DFCNQND2BWP40
    CLASS CORE ;
    FOREIGN DFCNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.050 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.690 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 -0.115 4.340 0.115 ;
        RECT  4.190 -0.115 4.260 0.475 ;
        RECT  3.810 -0.115 4.190 0.115 ;
        RECT  3.690 -0.115 3.810 0.145 ;
        RECT  3.095 -0.115 3.690 0.115 ;
        RECT  3.025 -0.115 3.095 0.405 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.145 4.340 1.375 ;
        RECT  4.190 0.715 4.260 1.375 ;
        RECT  3.830 1.145 4.190 1.375 ;
        RECT  3.710 1.025 3.830 1.375 ;
        RECT  3.415 1.145 3.710 1.375 ;
        RECT  3.325 1.095 3.415 1.375 ;
        RECT  3.215 1.145 3.325 1.375 ;
        RECT  3.145 0.985 3.215 1.375 ;
        RECT  2.335 1.145 3.145 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.790 0.220 3.870 0.660 ;
        RECT  3.235 0.220 3.790 0.295 ;
        RECT  3.455 0.925 3.620 1.000 ;
        RECT  3.385 0.375 3.455 1.000 ;
        RECT  3.310 0.375 3.385 0.445 ;
        RECT  3.055 0.630 3.385 0.700 ;
        RECT  3.200 0.815 3.300 0.915 ;
        RECT  3.165 0.220 3.235 0.560 ;
        RECT  2.655 0.845 3.200 0.915 ;
        RECT  2.975 0.490 3.165 0.560 ;
        RECT  2.905 0.490 2.975 0.775 ;
        RECT  2.880 0.490 2.905 0.560 ;
        RECT  2.770 0.995 2.895 1.075 ;
        RECT  2.810 0.315 2.880 0.560 ;
        RECT  2.485 0.995 2.770 1.065 ;
        RECT  2.585 0.335 2.655 0.915 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.130 0.815 ;
        RECT  2.010 0.335 2.070 0.815 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.010 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQND2BWP40

MACRO DFCNQND4BWP40
    CLASS CORE ;
    FOREIGN DFCNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.745 4.640 1.000 ;
        RECT  4.545 0.205 4.630 0.485 ;
        RECT  4.515 0.355 4.545 0.485 ;
        RECT  4.515 0.745 4.530 0.830 ;
        RECT  4.305 0.355 4.515 0.830 ;
        RECT  4.250 0.355 4.305 0.455 ;
        RECT  4.250 0.745 4.305 0.830 ;
        RECT  4.165 0.205 4.250 0.455 ;
        RECT  4.165 0.745 4.250 1.035 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.005 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.495 3.895 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 4.900 0.115 ;
        RECT  4.750 -0.115 4.820 0.475 ;
        RECT  4.425 -0.115 4.750 0.115 ;
        RECT  4.355 -0.115 4.425 0.275 ;
        RECT  4.015 -0.115 4.355 0.115 ;
        RECT  3.895 -0.115 4.015 0.145 ;
        RECT  3.095 -0.115 3.895 0.115 ;
        RECT  3.025 -0.115 3.095 0.285 ;
        RECT  2.210 -0.115 3.025 0.115 ;
        RECT  2.140 -0.115 2.210 0.430 ;
        RECT  1.755 -0.115 2.140 0.115 ;
        RECT  1.685 -0.115 1.755 0.335 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.265 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 4.900 1.375 ;
        RECT  4.750 0.710 4.820 1.375 ;
        RECT  4.425 1.145 4.750 1.375 ;
        RECT  4.355 0.915 4.425 1.375 ;
        RECT  4.010 1.145 4.355 1.375 ;
        RECT  3.940 0.835 4.010 1.375 ;
        RECT  3.620 1.145 3.940 1.375 ;
        RECT  3.530 1.095 3.620 1.375 ;
        RECT  3.215 1.145 3.530 1.375 ;
        RECT  3.085 1.035 3.215 1.375 ;
        RECT  2.335 1.145 3.085 1.375 ;
        RECT  2.225 1.040 2.335 1.375 ;
        RECT  1.660 1.145 2.225 1.375 ;
        RECT  1.540 1.070 1.660 1.375 ;
        RECT  0.710 1.145 1.540 1.375 ;
        RECT  0.590 1.020 0.710 1.375 ;
        RECT  0.345 1.145 0.590 1.375 ;
        RECT  0.215 0.990 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.745 4.640 1.000 ;
        RECT  4.585 0.205 4.630 0.485 ;
        RECT  4.165 0.205 4.235 0.455 ;
        RECT  4.165 0.745 4.235 1.035 ;
        RECT  4.075 0.545 4.235 0.615 ;
        RECT  3.995 0.220 4.075 0.615 ;
        RECT  3.325 0.220 3.995 0.295 ;
        RECT  3.660 0.925 3.825 1.000 ;
        RECT  3.590 0.375 3.660 1.000 ;
        RECT  3.515 0.375 3.590 0.445 ;
        RECT  3.135 0.545 3.590 0.615 ;
        RECT  3.415 0.855 3.490 1.005 ;
        RECT  3.045 0.855 3.415 0.925 ;
        RECT  2.975 0.705 3.410 0.775 ;
        RECT  3.255 0.220 3.325 0.425 ;
        RECT  2.975 0.355 3.255 0.425 ;
        RECT  2.975 0.845 3.045 0.925 ;
        RECT  2.905 0.355 2.975 0.775 ;
        RECT  2.655 0.845 2.975 0.915 ;
        RECT  2.785 0.355 2.905 0.425 ;
        RECT  2.770 0.995 2.895 1.075 ;
        RECT  2.485 0.995 2.770 1.065 ;
        RECT  2.585 0.335 2.655 0.915 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.405 0.195 2.415 0.960 ;
        RECT  2.070 0.890 2.405 0.960 ;
        RECT  2.070 0.640 2.145 0.815 ;
        RECT  2.025 0.335 2.070 0.815 ;
        RECT  1.980 0.890 2.070 1.000 ;
        RECT  2.000 0.335 2.025 0.720 ;
        RECT  1.880 0.335 2.000 0.405 ;
        RECT  1.475 0.650 2.000 0.720 ;
        RECT  1.470 0.930 1.980 1.000 ;
        RECT  1.615 0.510 1.920 0.580 ;
        RECT  1.330 0.790 1.835 0.860 ;
        RECT  1.545 0.215 1.615 0.580 ;
        RECT  0.775 0.215 1.545 0.285 ;
        RECT  1.405 0.600 1.475 0.720 ;
        RECT  1.400 0.930 1.470 1.065 ;
        RECT  1.190 0.995 1.400 1.065 ;
        RECT  1.260 0.365 1.330 0.910 ;
        RECT  1.120 0.520 1.190 1.065 ;
        RECT  1.110 0.905 1.120 1.065 ;
        RECT  0.860 0.905 1.110 0.985 ;
        RECT  0.980 0.705 1.050 0.825 ;
        RECT  0.775 0.705 0.980 0.775 ;
        RECT  0.790 0.875 0.860 0.985 ;
        RECT  0.625 0.875 0.790 0.945 ;
        RECT  0.705 0.215 0.775 0.775 ;
        RECT  0.555 0.255 0.625 0.945 ;
        RECT  0.415 0.255 0.555 0.325 ;
        RECT  0.505 0.875 0.555 0.945 ;
        RECT  0.435 0.875 0.505 1.030 ;
        RECT  0.345 0.520 0.385 0.640 ;
        RECT  0.275 0.345 0.345 0.910 ;
        RECT  0.125 0.345 0.275 0.415 ;
        RECT  0.140 0.840 0.275 0.910 ;
        RECT  0.055 0.840 0.140 1.030 ;
        RECT  0.055 0.230 0.125 0.415 ;
    END
END DFCNQND4BWP40

MACRO DFCSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.215 4.585 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.410 -0.115 4.620 0.115 ;
        RECT  4.275 -0.115 4.410 0.350 ;
        RECT  3.380 -0.115 4.275 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.410 ;
        RECT  2.095 -0.115 2.475 0.115 ;
        RECT  1.995 -0.115 2.095 0.425 ;
        RECT  0.730 -0.115 1.995 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.235 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.970 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.565 1.130 0.690 1.375 ;
        RECT  0.370 1.145 0.565 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.060 ;
        RECT  4.080 0.740 4.095 1.060 ;
        RECT  3.950 0.740 4.080 0.810 ;
        RECT  3.805 0.510 4.025 0.630 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.880 0.740 3.950 1.000 ;
        RECT  2.940 0.930 3.880 1.000 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.790 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.365 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.825 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.280 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.395 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.415 0.225 1.915 0.295 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.255 0.850 1.820 0.920 ;
        RECT  1.255 0.365 1.730 0.435 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.325 0.505 1.395 0.730 ;
        RECT  1.185 0.365 1.255 0.920 ;
        RECT  1.095 0.185 1.205 0.285 ;
        RECT  1.035 0.355 1.105 0.910 ;
        RECT  1.090 0.205 1.095 0.285 ;
        RECT  0.955 0.205 1.090 0.275 ;
        RECT  0.960 0.835 1.035 0.910 ;
        RECT  0.885 0.205 0.955 0.420 ;
        RECT  0.760 0.350 0.885 0.420 ;
        RECT  0.750 0.905 0.825 1.060 ;
        RECT  0.685 0.350 0.760 0.800 ;
        RECT  0.360 0.905 0.750 0.975 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.535 0.705 0.685 0.800 ;
        RECT  0.460 0.195 0.540 0.420 ;
        RECT  0.440 0.705 0.535 0.825 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.975 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.140 0.875 0.290 0.975 ;
        RECT  0.080 0.195 0.160 0.410 ;
        RECT  0.060 0.875 0.140 0.995 ;
        LAYER VIA1 ;
        RECT  2.335 0.385 2.405 0.455 ;
        RECT  1.035 0.385 1.105 0.455 ;
        LAYER M2 ;
        RECT  0.985 0.385 2.475 0.455 ;
    END
END DFCSNQD0BWP40

MACRO DFCSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.200 4.585 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.032200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.385 -0.115 4.620 0.115 ;
        RECT  4.295 -0.115 4.385 0.310 ;
        RECT  3.380 -0.115 4.295 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.410 ;
        RECT  2.095 -0.115 2.475 0.115 ;
        RECT  1.995 -0.115 2.095 0.430 ;
        RECT  0.730 -0.115 1.995 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.235 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.955 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.565 1.130 0.690 1.375 ;
        RECT  0.370 1.145 0.565 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.000 ;
        RECT  2.940 0.930 4.095 1.000 ;
        RECT  3.805 0.460 4.025 0.580 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.825 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.300 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.395 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.225 1.915 0.295 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.255 0.850 1.820 0.920 ;
        RECT  1.255 0.365 1.735 0.435 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.325 0.505 1.395 0.730 ;
        RECT  1.185 0.365 1.255 0.920 ;
        RECT  1.095 0.185 1.205 0.285 ;
        RECT  1.035 0.355 1.105 0.910 ;
        RECT  1.090 0.205 1.095 0.285 ;
        RECT  0.955 0.205 1.090 0.275 ;
        RECT  0.960 0.835 1.035 0.910 ;
        RECT  0.885 0.205 0.955 0.420 ;
        RECT  0.760 0.350 0.885 0.420 ;
        RECT  0.750 0.905 0.825 1.060 ;
        RECT  0.685 0.350 0.760 0.800 ;
        RECT  0.360 0.905 0.750 0.975 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.535 0.705 0.685 0.800 ;
        RECT  0.460 0.195 0.540 0.420 ;
        RECT  0.440 0.705 0.535 0.825 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.975 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.140 0.875 0.290 0.975 ;
        RECT  0.080 0.195 0.160 0.410 ;
        RECT  0.060 0.875 0.140 0.995 ;
        LAYER VIA1 ;
        RECT  2.335 0.385 2.405 0.455 ;
        RECT  1.035 0.385 1.105 0.455 ;
        LAYER M2 ;
        RECT  0.985 0.385 2.455 0.455 ;
    END
END DFCSNQD1BWP40

MACRO DFCSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.195 4.585 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.032200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 -0.115 4.900 0.115 ;
        RECT  4.760 -0.115 4.830 0.485 ;
        RECT  4.410 -0.115 4.760 0.115 ;
        RECT  4.275 -0.115 4.410 0.310 ;
        RECT  3.380 -0.115 4.275 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.410 ;
        RECT  2.095 -0.115 2.475 0.115 ;
        RECT  1.995 -0.115 2.095 0.430 ;
        RECT  0.730 -0.115 1.995 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.235 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 1.145 4.900 1.375 ;
        RECT  4.760 0.690 4.830 1.375 ;
        RECT  4.400 1.145 4.760 1.375 ;
        RECT  4.280 0.845 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.565 1.130 0.690 1.375 ;
        RECT  0.370 1.145 0.565 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.000 ;
        RECT  2.940 0.930 4.095 1.000 ;
        RECT  3.805 0.460 4.025 0.580 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.825 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.300 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.395 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.225 1.915 0.295 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.255 0.850 1.820 0.920 ;
        RECT  1.255 0.365 1.725 0.435 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.325 0.505 1.395 0.730 ;
        RECT  1.185 0.365 1.255 0.920 ;
        RECT  1.095 0.185 1.205 0.285 ;
        RECT  1.035 0.355 1.105 0.910 ;
        RECT  1.090 0.205 1.095 0.285 ;
        RECT  0.955 0.205 1.090 0.275 ;
        RECT  0.960 0.835 1.035 0.910 ;
        RECT  0.885 0.205 0.955 0.420 ;
        RECT  0.760 0.350 0.885 0.420 ;
        RECT  0.750 0.905 0.825 1.060 ;
        RECT  0.685 0.350 0.760 0.800 ;
        RECT  0.360 0.905 0.750 0.975 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.535 0.705 0.685 0.800 ;
        RECT  0.460 0.195 0.540 0.420 ;
        RECT  0.440 0.705 0.535 0.825 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.975 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.140 0.875 0.290 0.975 ;
        RECT  0.080 0.195 0.160 0.410 ;
        RECT  0.060 0.875 0.140 0.995 ;
        LAYER VIA1 ;
        RECT  2.335 0.385 2.405 0.455 ;
        RECT  1.035 0.385 1.105 0.455 ;
        LAYER M2 ;
        RECT  0.985 0.385 2.455 0.455 ;
    END
END DFCSNQD2BWP40

MACRO DFCSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.450 4.890 0.765 ;
        RECT  4.785 0.525 4.795 0.635 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.425 0.195 5.520 0.485 ;
        RECT  5.425 0.710 5.520 0.995 ;
        RECT  5.355 0.355 5.425 0.485 ;
        RECT  5.355 0.710 5.425 0.830 ;
        RECT  5.145 0.355 5.355 0.830 ;
        RECT  5.120 0.355 5.145 0.485 ;
        RECT  5.120 0.710 5.145 0.830 ;
        RECT  5.045 0.215 5.120 0.485 ;
        RECT  5.045 0.710 5.120 0.995 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.044600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.335 0.355 3.465 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 -0.115 5.740 0.115 ;
        RECT  5.615 -0.115 5.685 0.440 ;
        RECT  5.310 -0.115 5.615 0.115 ;
        RECT  5.225 -0.115 5.310 0.265 ;
        RECT  4.940 -0.115 5.225 0.115 ;
        RECT  4.850 -0.115 4.940 0.310 ;
        RECT  4.190 -0.115 4.850 0.115 ;
        RECT  4.070 -0.115 4.190 0.140 ;
        RECT  3.390 -0.115 4.070 0.115 ;
        RECT  3.255 -0.115 3.390 0.130 ;
        RECT  2.545 -0.115 3.255 0.115 ;
        RECT  2.475 -0.115 2.545 0.410 ;
        RECT  2.095 -0.115 2.475 0.115 ;
        RECT  1.995 -0.115 2.095 0.430 ;
        RECT  0.730 -0.115 1.995 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.235 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.145 5.740 1.375 ;
        RECT  5.615 0.680 5.685 1.375 ;
        RECT  5.330 1.145 5.615 1.375 ;
        RECT  5.210 0.910 5.330 1.375 ;
        RECT  4.930 1.145 5.210 1.375 ;
        RECT  4.855 0.845 4.930 1.375 ;
        RECT  4.020 1.145 4.855 1.375 ;
        RECT  3.900 1.070 4.020 1.375 ;
        RECT  3.390 1.145 3.900 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.690 1.145 1.530 1.375 ;
        RECT  0.565 1.130 0.690 1.375 ;
        RECT  0.370 1.145 0.565 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.195 5.520 0.485 ;
        RECT  5.425 0.710 5.520 0.995 ;
        RECT  5.045 0.215 5.075 0.485 ;
        RECT  5.045 0.710 5.075 0.995 ;
        RECT  4.645 0.210 4.715 1.000 ;
        RECT  4.065 0.930 4.645 1.000 ;
        RECT  4.535 0.620 4.575 0.740 ;
        RECT  4.465 0.210 4.535 0.860 ;
        RECT  3.785 0.210 4.465 0.280 ;
        RECT  4.350 0.790 4.465 0.860 ;
        RECT  3.865 0.350 4.370 0.420 ;
        RECT  3.985 0.605 4.065 1.000 ;
        RECT  2.940 0.930 3.985 1.000 ;
        RECT  3.715 0.210 3.785 0.860 ;
        RECT  3.710 0.335 3.715 0.860 ;
        RECT  3.695 0.335 3.710 0.445 ;
        RECT  3.225 0.790 3.710 0.860 ;
        RECT  3.605 0.580 3.640 0.700 ;
        RECT  3.535 0.200 3.605 0.700 ;
        RECT  3.000 0.200 3.535 0.270 ;
        RECT  3.155 0.445 3.225 0.860 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 3.000 0.270 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.825 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.300 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.395 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.225 1.915 0.295 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.255 0.850 1.820 0.920 ;
        RECT  1.255 0.365 1.730 0.435 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.325 0.505 1.395 0.730 ;
        RECT  1.185 0.365 1.255 0.920 ;
        RECT  1.095 0.185 1.205 0.285 ;
        RECT  1.035 0.355 1.105 0.910 ;
        RECT  1.090 0.205 1.095 0.285 ;
        RECT  0.955 0.205 1.090 0.275 ;
        RECT  0.960 0.835 1.035 0.910 ;
        RECT  0.885 0.205 0.955 0.420 ;
        RECT  0.760 0.350 0.885 0.420 ;
        RECT  0.750 0.905 0.825 1.060 ;
        RECT  0.685 0.350 0.760 0.800 ;
        RECT  0.360 0.905 0.750 0.975 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.535 0.705 0.685 0.800 ;
        RECT  0.460 0.195 0.540 0.420 ;
        RECT  0.440 0.705 0.535 0.825 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.975 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.140 0.875 0.290 0.975 ;
        RECT  0.080 0.195 0.160 0.410 ;
        RECT  0.060 0.875 0.140 0.995 ;
        LAYER VIA1 ;
        RECT  2.335 0.385 2.405 0.455 ;
        RECT  1.035 0.385 1.105 0.455 ;
        LAYER M2 ;
        RECT  0.985 0.385 2.455 0.455 ;
    END
END DFCSNQD4BWP40

MACRO DFKCNQD0BWP40
    CLASS CORE ;
    FOREIGN DFKCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.050000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.215 3.465 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.010 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.485 0.805 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.115 3.500 0.115 ;
        RECT  3.150 -0.115 3.270 0.280 ;
        RECT  2.855 -0.115 3.150 0.115 ;
        RECT  2.785 -0.115 2.855 0.305 ;
        RECT  2.110 -0.115 2.785 0.115 ;
        RECT  1.990 -0.115 2.110 0.190 ;
        RECT  1.790 -0.115 1.990 0.115 ;
        RECT  1.670 -0.115 1.790 0.190 ;
        RECT  0.730 -0.115 1.670 0.115 ;
        RECT  0.610 -0.115 0.730 0.125 ;
        RECT  0.360 -0.115 0.610 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.245 1.145 3.500 1.375 ;
        RECT  3.175 0.945 3.245 1.375 ;
        RECT  2.870 1.145 3.175 1.375 ;
        RECT  2.800 0.950 2.870 1.375 ;
        RECT  2.125 1.145 2.800 1.375 ;
        RECT  2.050 0.785 2.125 1.375 ;
        RECT  1.725 1.145 2.050 1.375 ;
        RECT  1.655 0.860 1.725 1.375 ;
        RECT  0.910 1.145 1.655 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.370 1.145 0.790 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.375 3.300 0.805 ;
        RECT  3.045 0.375 3.230 0.445 ;
        RECT  3.050 0.735 3.230 0.805 ;
        RECT  2.910 0.545 3.150 0.615 ;
        RECT  2.980 0.735 3.050 1.065 ;
        RECT  2.975 0.240 3.045 0.445 ;
        RECT  2.770 0.375 2.975 0.445 ;
        RECT  2.840 0.545 2.910 0.805 ;
        RECT  2.730 0.735 2.840 0.805 ;
        RECT  2.690 0.375 2.770 0.640 ;
        RECT  2.660 0.735 2.730 1.060 ;
        RECT  2.400 0.990 2.660 1.060 ;
        RECT  2.585 0.200 2.615 0.640 ;
        RECT  2.545 0.200 2.585 0.910 ;
        RECT  2.410 0.200 2.545 0.270 ;
        RECT  2.515 0.570 2.545 0.910 ;
        RECT  2.400 0.355 2.475 0.475 ;
        RECT  2.290 0.185 2.410 0.270 ;
        RECT  2.330 0.355 2.400 1.060 ;
        RECT  1.885 0.345 1.955 0.960 ;
        RECT  1.855 0.345 1.885 0.455 ;
        RECT  1.865 0.700 1.885 0.960 ;
        RECT  1.640 0.700 1.865 0.770 ;
        RECT  1.785 0.515 1.815 0.625 ;
        RECT  1.715 0.260 1.785 0.625 ;
        RECT  1.360 0.260 1.715 0.330 ;
        RECT  1.570 0.650 1.640 0.770 ;
        RECT  1.500 0.400 1.580 0.470 ;
        RECT  1.500 0.840 1.550 0.910 ;
        RECT  1.430 0.400 1.500 0.910 ;
        RECT  1.290 0.980 1.420 1.075 ;
        RECT  1.290 0.260 1.360 0.910 ;
        RECT  1.190 0.840 1.290 0.910 ;
        RECT  0.340 0.980 1.290 1.050 ;
        RECT  1.130 0.195 1.205 0.490 ;
        RECT  1.125 0.570 1.205 0.770 ;
        RECT  0.340 0.195 1.130 0.265 ;
        RECT  0.520 0.700 1.125 0.770 ;
        RECT  0.590 0.840 1.110 0.910 ;
        RECT  0.520 0.345 0.580 0.415 ;
        RECT  0.505 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.505 0.910 ;
        RECT  0.435 0.695 0.450 0.910 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.195 0.340 1.050 ;
        RECT  0.055 0.280 0.270 0.400 ;
        RECT  0.055 0.840 0.270 0.960 ;
    END
END DFKCNQD0BWP40

MACRO DFKCNQD1BWP40
    CLASS CORE ;
    FOREIGN DFKCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.185 3.465 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.990 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.485 0.805 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.245 -0.115 3.500 0.115 ;
        RECT  3.175 -0.115 3.245 0.305 ;
        RECT  2.855 -0.115 3.175 0.115 ;
        RECT  2.785 -0.115 2.855 0.325 ;
        RECT  2.105 -0.115 2.785 0.115 ;
        RECT  1.985 -0.115 2.105 0.125 ;
        RECT  1.740 -0.115 1.985 0.115 ;
        RECT  1.620 -0.115 1.740 0.125 ;
        RECT  0.720 -0.115 1.620 0.115 ;
        RECT  0.600 -0.115 0.720 0.125 ;
        RECT  0.360 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.245 1.145 3.500 1.375 ;
        RECT  3.175 0.860 3.245 1.375 ;
        RECT  2.870 1.145 3.175 1.375 ;
        RECT  2.800 0.950 2.870 1.375 ;
        RECT  2.125 1.145 2.800 1.375 ;
        RECT  2.050 0.690 2.125 1.375 ;
        RECT  1.725 1.145 2.050 1.375 ;
        RECT  1.655 0.860 1.725 1.375 ;
        RECT  0.910 1.145 1.655 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.370 1.145 0.790 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.395 3.300 0.775 ;
        RECT  3.045 0.395 3.230 0.465 ;
        RECT  3.050 0.705 3.230 0.775 ;
        RECT  2.910 0.545 3.150 0.615 ;
        RECT  2.980 0.705 3.050 1.000 ;
        RECT  2.975 0.215 3.045 0.465 ;
        RECT  2.770 0.395 2.975 0.465 ;
        RECT  2.840 0.545 2.910 0.805 ;
        RECT  2.720 0.735 2.840 0.805 ;
        RECT  2.690 0.395 2.770 0.640 ;
        RECT  2.650 0.735 2.720 1.065 ;
        RECT  2.430 0.995 2.650 1.065 ;
        RECT  2.580 0.195 2.615 0.640 ;
        RECT  2.545 0.195 2.580 0.915 ;
        RECT  1.400 0.195 2.545 0.265 ;
        RECT  2.510 0.570 2.545 0.915 ;
        RECT  2.430 0.355 2.475 0.475 ;
        RECT  2.360 0.355 2.430 1.065 ;
        RECT  1.885 0.340 1.955 0.960 ;
        RECT  1.855 0.340 1.885 0.450 ;
        RECT  1.865 0.700 1.885 0.960 ;
        RECT  1.640 0.700 1.865 0.770 ;
        RECT  1.785 0.515 1.815 0.625 ;
        RECT  1.715 0.345 1.785 0.625 ;
        RECT  1.330 0.345 1.715 0.415 ;
        RECT  1.570 0.650 1.640 0.770 ;
        RECT  1.500 0.485 1.560 0.555 ;
        RECT  1.500 0.840 1.550 0.910 ;
        RECT  1.430 0.485 1.500 0.910 ;
        RECT  1.290 0.980 1.420 1.075 ;
        RECT  1.260 0.195 1.330 0.910 ;
        RECT  0.340 0.980 1.290 1.050 ;
        RECT  1.200 0.195 1.260 0.295 ;
        RECT  1.190 0.840 1.260 0.910 ;
        RECT  1.130 0.380 1.190 0.500 ;
        RECT  1.100 0.570 1.190 0.770 ;
        RECT  1.060 0.195 1.130 0.500 ;
        RECT  0.590 0.840 1.110 0.910 ;
        RECT  0.520 0.700 1.100 0.770 ;
        RECT  0.340 0.195 1.060 0.265 ;
        RECT  0.520 0.345 0.580 0.415 ;
        RECT  0.505 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.505 0.910 ;
        RECT  0.435 0.695 0.450 0.910 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.195 0.340 1.050 ;
        RECT  0.055 0.280 0.270 0.400 ;
        RECT  0.055 0.840 0.270 0.960 ;
    END
END DFKCNQD1BWP40

MACRO DFKCNQD2BWP40
    CLASS CORE ;
    FOREIGN DFKCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.385 0.185 3.475 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.990 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.485 0.805 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.710 -0.115 3.780 0.115 ;
        RECT  3.625 -0.115 3.710 0.470 ;
        RECT  3.245 -0.115 3.625 0.115 ;
        RECT  3.175 -0.115 3.245 0.300 ;
        RECT  2.855 -0.115 3.175 0.115 ;
        RECT  2.785 -0.115 2.855 0.325 ;
        RECT  2.105 -0.115 2.785 0.115 ;
        RECT  1.985 -0.115 2.105 0.125 ;
        RECT  1.740 -0.115 1.985 0.115 ;
        RECT  1.620 -0.115 1.740 0.125 ;
        RECT  0.720 -0.115 1.620 0.115 ;
        RECT  0.600 -0.115 0.720 0.125 ;
        RECT  0.360 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.710 1.145 3.780 1.375 ;
        RECT  3.625 0.670 3.710 1.375 ;
        RECT  3.245 1.145 3.625 1.375 ;
        RECT  3.175 0.860 3.245 1.375 ;
        RECT  2.870 1.145 3.175 1.375 ;
        RECT  2.800 0.950 2.870 1.375 ;
        RECT  2.125 1.145 2.800 1.375 ;
        RECT  2.050 0.690 2.125 1.375 ;
        RECT  1.725 1.145 2.050 1.375 ;
        RECT  1.655 0.860 1.725 1.375 ;
        RECT  0.910 1.145 1.655 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.370 1.145 0.790 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.240 0.395 3.310 0.775 ;
        RECT  3.045 0.395 3.240 0.465 ;
        RECT  3.050 0.705 3.240 0.775 ;
        RECT  2.910 0.545 3.150 0.615 ;
        RECT  2.980 0.705 3.050 1.000 ;
        RECT  2.975 0.215 3.045 0.465 ;
        RECT  2.770 0.395 2.975 0.465 ;
        RECT  2.840 0.545 2.910 0.805 ;
        RECT  2.720 0.735 2.840 0.805 ;
        RECT  2.690 0.395 2.770 0.640 ;
        RECT  2.650 0.735 2.720 1.065 ;
        RECT  2.430 0.995 2.650 1.065 ;
        RECT  2.580 0.195 2.615 0.640 ;
        RECT  2.545 0.195 2.580 0.915 ;
        RECT  1.400 0.195 2.545 0.265 ;
        RECT  2.510 0.570 2.545 0.915 ;
        RECT  2.430 0.355 2.475 0.475 ;
        RECT  2.360 0.355 2.430 1.065 ;
        RECT  1.885 0.340 1.955 0.960 ;
        RECT  1.855 0.340 1.885 0.450 ;
        RECT  1.865 0.700 1.885 0.960 ;
        RECT  1.640 0.700 1.865 0.770 ;
        RECT  1.785 0.515 1.815 0.625 ;
        RECT  1.715 0.345 1.785 0.625 ;
        RECT  1.330 0.345 1.715 0.415 ;
        RECT  1.570 0.650 1.640 0.770 ;
        RECT  1.500 0.485 1.560 0.555 ;
        RECT  1.500 0.840 1.550 0.910 ;
        RECT  1.430 0.485 1.500 0.910 ;
        RECT  1.290 0.980 1.420 1.075 ;
        RECT  1.260 0.195 1.330 0.910 ;
        RECT  0.340 0.980 1.290 1.050 ;
        RECT  1.200 0.195 1.260 0.295 ;
        RECT  1.190 0.840 1.260 0.910 ;
        RECT  1.130 0.380 1.190 0.500 ;
        RECT  1.100 0.570 1.190 0.770 ;
        RECT  1.060 0.195 1.130 0.500 ;
        RECT  0.590 0.840 1.110 0.910 ;
        RECT  0.520 0.700 1.100 0.770 ;
        RECT  0.340 0.195 1.060 0.265 ;
        RECT  0.520 0.345 0.580 0.415 ;
        RECT  0.505 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.505 0.910 ;
        RECT  0.435 0.695 0.450 0.910 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.195 0.340 1.050 ;
        RECT  0.055 0.280 0.270 0.400 ;
        RECT  0.055 0.840 0.270 0.960 ;
    END
END DFKCNQD2BWP40

MACRO DFKCNQD4BWP40
    CLASS CORE ;
    FOREIGN DFKCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.005 0.205 4.095 0.470 ;
        RECT  4.005 0.685 4.095 1.075 ;
        RECT  3.955 0.385 4.005 0.470 ;
        RECT  3.955 0.685 4.005 0.770 ;
        RECT  3.745 0.385 3.955 0.770 ;
        RECT  3.735 0.385 3.745 0.470 ;
        RECT  3.735 0.685 3.745 0.770 ;
        RECT  3.645 0.210 3.735 0.470 ;
        RECT  3.645 0.685 3.735 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.990 0.630 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.485 0.805 0.630 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 -0.115 4.340 0.115 ;
        RECT  4.215 -0.115 4.290 0.445 ;
        RECT  3.905 -0.115 4.215 0.115 ;
        RECT  3.835 -0.115 3.905 0.255 ;
        RECT  3.505 -0.115 3.835 0.115 ;
        RECT  3.435 -0.115 3.505 0.265 ;
        RECT  3.100 -0.115 3.435 0.115 ;
        RECT  3.030 -0.115 3.100 0.265 ;
        RECT  2.920 -0.115 3.030 0.115 ;
        RECT  2.850 -0.115 2.920 0.400 ;
        RECT  2.160 -0.115 2.850 0.115 ;
        RECT  2.040 -0.115 2.160 0.125 ;
        RECT  1.740 -0.115 2.040 0.115 ;
        RECT  1.620 -0.115 1.740 0.125 ;
        RECT  0.720 -0.115 1.620 0.115 ;
        RECT  0.600 -0.115 0.720 0.125 ;
        RECT  0.360 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.360 0.125 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.215 0.715 4.290 1.375 ;
        RECT  3.905 1.145 4.215 1.375 ;
        RECT  3.835 0.885 3.905 1.375 ;
        RECT  3.505 1.145 3.835 1.375 ;
        RECT  3.435 1.020 3.505 1.375 ;
        RECT  3.100 1.145 3.435 1.375 ;
        RECT  3.030 0.865 3.100 1.375 ;
        RECT  2.925 1.145 3.030 1.375 ;
        RECT  2.855 0.835 2.925 1.375 ;
        RECT  2.160 1.145 2.855 1.375 ;
        RECT  2.090 0.670 2.160 1.375 ;
        RECT  1.725 1.145 2.090 1.375 ;
        RECT  1.655 0.860 1.725 1.375 ;
        RECT  0.910 1.145 1.655 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.370 1.145 0.790 1.375 ;
        RECT  0.250 1.130 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.025 0.205 4.095 0.470 ;
        RECT  4.025 0.685 4.095 1.075 ;
        RECT  3.645 0.210 3.675 0.470 ;
        RECT  3.645 0.685 3.675 1.075 ;
        RECT  3.575 0.545 3.615 0.615 ;
        RECT  3.505 0.365 3.575 0.895 ;
        RECT  3.290 0.365 3.505 0.435 ;
        RECT  3.290 0.825 3.505 0.895 ;
        RECT  3.220 0.205 3.290 0.435 ;
        RECT  3.220 0.525 3.290 0.755 ;
        RECT  3.220 0.825 3.290 1.075 ;
        RECT  3.070 0.365 3.220 0.435 ;
        RECT  2.785 0.685 3.220 0.755 ;
        RECT  3.000 0.365 3.070 0.575 ;
        RECT  2.830 0.505 3.000 0.575 ;
        RECT  2.760 0.505 2.830 0.615 ;
        RECT  2.715 0.685 2.785 1.015 ;
        RECT  2.495 0.945 2.715 1.015 ;
        RECT  2.645 0.195 2.680 0.620 ;
        RECT  2.610 0.195 2.645 0.795 ;
        RECT  1.400 0.195 2.610 0.265 ;
        RECT  2.575 0.550 2.610 0.795 ;
        RECT  2.495 0.350 2.540 0.470 ;
        RECT  2.425 0.350 2.495 1.015 ;
        RECT  1.885 0.340 1.955 0.960 ;
        RECT  1.855 0.340 1.885 0.450 ;
        RECT  1.865 0.700 1.885 0.960 ;
        RECT  1.640 0.700 1.865 0.770 ;
        RECT  1.785 0.515 1.815 0.625 ;
        RECT  1.715 0.345 1.785 0.625 ;
        RECT  1.330 0.345 1.715 0.415 ;
        RECT  1.570 0.650 1.640 0.770 ;
        RECT  1.500 0.485 1.560 0.555 ;
        RECT  1.500 0.840 1.550 0.910 ;
        RECT  1.430 0.485 1.500 0.910 ;
        RECT  1.290 0.980 1.420 1.075 ;
        RECT  1.260 0.195 1.330 0.910 ;
        RECT  0.340 0.980 1.290 1.050 ;
        RECT  1.200 0.195 1.260 0.295 ;
        RECT  1.190 0.840 1.260 0.910 ;
        RECT  1.130 0.380 1.190 0.500 ;
        RECT  1.100 0.570 1.190 0.770 ;
        RECT  1.060 0.195 1.130 0.500 ;
        RECT  0.590 0.840 1.110 0.910 ;
        RECT  0.520 0.700 1.100 0.770 ;
        RECT  0.340 0.195 1.060 0.265 ;
        RECT  0.520 0.345 0.580 0.415 ;
        RECT  0.505 0.345 0.520 0.770 ;
        RECT  0.450 0.345 0.505 0.910 ;
        RECT  0.435 0.695 0.450 0.910 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.195 0.340 1.050 ;
        RECT  0.055 0.280 0.270 0.400 ;
        RECT  0.055 0.840 0.270 0.960 ;
    END
END DFKCNQD4BWP40

MACRO DFKCSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFKCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.190 0.675 ;
        RECT  0.035 0.495 0.130 0.770 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.680 0.575 0.800 ;
        RECT  0.455 0.680 0.545 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.225 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.011800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.985 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.305 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.305 ;
        RECT  2.675 -0.115 3.375 0.115 ;
        RECT  2.605 -0.115 2.675 0.445 ;
        RECT  2.300 -0.115 2.605 0.115 ;
        RECT  2.180 -0.115 2.300 0.210 ;
        RECT  1.300 -0.115 2.180 0.115 ;
        RECT  1.180 -0.115 1.300 0.125 ;
        RECT  0.340 -0.115 1.180 0.115 ;
        RECT  0.180 -0.115 0.340 0.125 ;
        RECT  0.000 -0.115 0.180 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.950 3.815 1.375 ;
        RECT  3.450 1.145 3.745 1.375 ;
        RECT  3.380 0.895 3.450 1.375 ;
        RECT  2.675 1.145 3.380 1.375 ;
        RECT  2.605 0.785 2.675 1.375 ;
        RECT  2.295 1.145 2.605 1.375 ;
        RECT  2.185 0.890 2.295 1.375 ;
        RECT  1.300 1.145 2.185 1.375 ;
        RECT  1.180 1.135 1.300 1.375 ;
        RECT  0.950 1.145 1.180 1.375 ;
        RECT  0.830 1.135 0.950 1.375 ;
        RECT  0.340 1.145 0.830 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.405 3.855 0.820 ;
        RECT  3.635 0.405 3.785 0.475 ;
        RECT  3.635 0.750 3.785 0.820 ;
        RECT  3.565 0.185 3.635 0.475 ;
        RECT  3.565 0.750 3.635 1.015 ;
        RECT  3.310 0.545 3.585 0.615 ;
        RECT  3.270 0.405 3.565 0.475 ;
        RECT  3.240 0.545 3.310 1.045 ;
        RECT  3.180 0.545 3.240 0.615 ;
        RECT  2.960 0.975 3.240 1.045 ;
        RECT  3.110 0.240 3.180 0.615 ;
        RECT  3.100 0.770 3.170 0.890 ;
        RECT  2.960 0.240 3.110 0.310 ;
        RECT  2.985 0.770 3.100 0.840 ;
        RECT  2.915 0.440 2.985 0.840 ;
        RECT  2.410 0.300 2.480 0.980 ;
        RECT  2.195 0.745 2.410 0.815 ;
        RECT  2.270 0.280 2.340 0.640 ;
        RECT  1.875 0.280 2.270 0.350 ;
        RECT  2.125 0.695 2.195 0.815 ;
        RECT  2.035 0.420 2.110 0.490 ;
        RECT  2.035 0.885 2.105 0.955 ;
        RECT  1.965 0.420 2.035 0.955 ;
        RECT  1.805 0.205 1.875 0.925 ;
        RECT  1.665 0.395 1.735 0.785 ;
        RECT  1.615 0.195 1.690 0.320 ;
        RECT  1.615 0.865 1.685 1.065 ;
        RECT  1.510 0.395 1.665 0.465 ;
        RECT  1.510 0.715 1.665 0.785 ;
        RECT  0.595 0.195 1.615 0.265 ;
        RECT  0.695 0.995 1.615 1.065 ;
        RECT  1.440 0.345 1.510 0.465 ;
        RECT  1.440 0.715 1.510 0.915 ;
        RECT  1.370 0.545 1.430 0.615 ;
        RECT  1.300 0.345 1.370 0.915 ;
        RECT  1.010 0.345 1.300 0.415 ;
        RECT  0.990 0.845 1.300 0.915 ;
        RECT  0.505 0.335 0.930 0.405 ;
        RECT  0.690 0.530 0.790 0.630 ;
        RECT  0.625 0.955 0.695 1.065 ;
        RECT  0.385 0.530 0.690 0.600 ;
        RECT  0.435 0.335 0.505 0.445 ;
        RECT  0.365 0.530 0.385 0.940 ;
        RECT  0.295 0.355 0.365 0.940 ;
        RECT  0.125 0.355 0.295 0.425 ;
        RECT  0.125 0.870 0.295 0.940 ;
        RECT  0.055 0.305 0.125 0.425 ;
        RECT  0.055 0.870 0.125 1.075 ;
    END
END DFKCSNQD0BWP40

MACRO DFKCSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFKCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.190 0.675 ;
        RECT  0.035 0.495 0.130 0.770 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.680 0.575 0.800 ;
        RECT  0.455 0.680 0.545 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.225 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.985 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.305 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.325 ;
        RECT  2.675 -0.115 3.375 0.115 ;
        RECT  2.605 -0.115 2.675 0.435 ;
        RECT  2.300 -0.115 2.605 0.115 ;
        RECT  2.180 -0.115 2.300 0.210 ;
        RECT  1.300 -0.115 2.180 0.115 ;
        RECT  1.180 -0.115 1.300 0.125 ;
        RECT  0.320 -0.115 1.180 0.115 ;
        RECT  0.200 -0.115 0.320 0.125 ;
        RECT  0.000 -0.115 0.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.860 3.815 1.375 ;
        RECT  3.450 1.145 3.745 1.375 ;
        RECT  3.380 0.720 3.450 1.375 ;
        RECT  2.675 1.145 3.380 1.375 ;
        RECT  2.605 0.690 2.675 1.375 ;
        RECT  2.275 1.145 2.605 1.375 ;
        RECT  2.205 0.865 2.275 1.375 ;
        RECT  1.300 1.145 2.205 1.375 ;
        RECT  1.180 1.135 1.300 1.375 ;
        RECT  0.950 1.145 1.180 1.375 ;
        RECT  0.830 1.135 0.950 1.375 ;
        RECT  0.340 1.145 0.830 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.780 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.710 3.775 0.780 ;
        RECT  3.565 0.205 3.635 0.465 ;
        RECT  3.565 0.710 3.635 1.075 ;
        RECT  3.310 0.545 3.585 0.615 ;
        RECT  3.230 0.395 3.565 0.465 ;
        RECT  3.240 0.545 3.310 1.045 ;
        RECT  3.160 0.545 3.240 0.615 ;
        RECT  2.960 0.975 3.240 1.045 ;
        RECT  3.100 0.770 3.170 0.890 ;
        RECT  3.090 0.240 3.160 0.615 ;
        RECT  2.990 0.770 3.100 0.840 ;
        RECT  2.960 0.240 3.090 0.310 ;
        RECT  2.920 0.440 2.990 0.840 ;
        RECT  2.410 0.300 2.480 0.980 ;
        RECT  2.395 0.300 2.410 0.415 ;
        RECT  2.395 0.720 2.410 0.980 ;
        RECT  2.205 0.720 2.395 0.790 ;
        RECT  2.325 0.470 2.340 0.590 ;
        RECT  2.255 0.280 2.325 0.590 ;
        RECT  1.900 0.280 2.255 0.350 ;
        RECT  2.135 0.670 2.205 0.790 ;
        RECT  2.045 0.885 2.105 0.955 ;
        RECT  2.045 0.420 2.100 0.490 ;
        RECT  1.975 0.420 2.045 0.955 ;
        RECT  1.830 0.195 1.900 0.960 ;
        RECT  1.785 0.195 1.830 0.265 ;
        RECT  1.690 0.395 1.760 0.785 ;
        RECT  0.615 0.195 1.705 0.265 ;
        RECT  1.600 0.855 1.700 1.065 ;
        RECT  1.510 0.395 1.690 0.465 ;
        RECT  1.510 0.715 1.690 0.785 ;
        RECT  0.695 0.995 1.600 1.065 ;
        RECT  1.440 0.345 1.510 0.465 ;
        RECT  1.440 0.715 1.510 0.910 ;
        RECT  1.370 0.545 1.440 0.615 ;
        RECT  1.300 0.355 1.370 0.925 ;
        RECT  1.010 0.355 1.300 0.425 ;
        RECT  0.990 0.855 1.300 0.925 ;
        RECT  0.410 0.355 0.930 0.425 ;
        RECT  0.385 0.535 0.795 0.605 ;
        RECT  0.625 0.925 0.695 1.065 ;
        RECT  0.340 0.535 0.385 0.940 ;
        RECT  0.270 0.355 0.340 0.940 ;
        RECT  0.125 0.355 0.270 0.425 ;
        RECT  0.125 0.870 0.270 0.940 ;
        RECT  0.055 0.305 0.125 0.425 ;
        RECT  0.055 0.870 0.125 1.075 ;
    END
END DFKCSNQD1BWP40

MACRO DFKCSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFKCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.190 0.675 ;
        RECT  0.035 0.495 0.130 0.770 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.945 0.195 4.035 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.680 0.575 0.800 ;
        RECT  0.455 0.680 0.545 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.225 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.985 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.275 -0.115 4.340 0.115 ;
        RECT  4.195 -0.115 4.275 0.460 ;
        RECT  3.815 -0.115 4.195 0.115 ;
        RECT  3.745 -0.115 3.815 0.305 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.325 ;
        RECT  2.675 -0.115 3.375 0.115 ;
        RECT  2.605 -0.115 2.675 0.435 ;
        RECT  2.300 -0.115 2.605 0.115 ;
        RECT  2.180 -0.115 2.300 0.210 ;
        RECT  1.300 -0.115 2.180 0.115 ;
        RECT  1.180 -0.115 1.300 0.125 ;
        RECT  0.320 -0.115 1.180 0.115 ;
        RECT  0.200 -0.115 0.320 0.125 ;
        RECT  0.000 -0.115 0.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.275 1.145 4.340 1.375 ;
        RECT  4.195 0.700 4.275 1.375 ;
        RECT  3.815 1.145 4.195 1.375 ;
        RECT  3.745 0.860 3.815 1.375 ;
        RECT  3.450 1.145 3.745 1.375 ;
        RECT  3.380 0.720 3.450 1.375 ;
        RECT  2.675 1.145 3.380 1.375 ;
        RECT  2.605 0.690 2.675 1.375 ;
        RECT  2.275 1.145 2.605 1.375 ;
        RECT  2.205 0.865 2.275 1.375 ;
        RECT  1.300 1.145 2.205 1.375 ;
        RECT  1.180 1.135 1.300 1.375 ;
        RECT  0.950 1.145 1.180 1.375 ;
        RECT  0.830 1.135 0.950 1.375 ;
        RECT  0.340 1.145 0.830 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.780 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.710 3.775 0.780 ;
        RECT  3.565 0.205 3.635 0.465 ;
        RECT  3.565 0.710 3.635 1.075 ;
        RECT  3.310 0.545 3.585 0.615 ;
        RECT  3.230 0.395 3.565 0.465 ;
        RECT  3.240 0.545 3.310 1.045 ;
        RECT  3.160 0.545 3.240 0.615 ;
        RECT  2.960 0.975 3.240 1.045 ;
        RECT  3.100 0.770 3.170 0.890 ;
        RECT  3.090 0.240 3.160 0.615 ;
        RECT  2.990 0.770 3.100 0.840 ;
        RECT  2.960 0.240 3.090 0.310 ;
        RECT  2.920 0.440 2.990 0.840 ;
        RECT  2.410 0.300 2.480 0.980 ;
        RECT  2.395 0.300 2.410 0.415 ;
        RECT  2.395 0.720 2.410 0.980 ;
        RECT  2.205 0.720 2.395 0.790 ;
        RECT  2.325 0.470 2.340 0.590 ;
        RECT  2.255 0.280 2.325 0.590 ;
        RECT  1.900 0.280 2.255 0.350 ;
        RECT  2.135 0.670 2.205 0.790 ;
        RECT  2.045 0.885 2.105 0.955 ;
        RECT  2.045 0.420 2.100 0.490 ;
        RECT  1.975 0.420 2.045 0.955 ;
        RECT  1.830 0.195 1.900 0.960 ;
        RECT  1.785 0.195 1.830 0.265 ;
        RECT  1.690 0.395 1.760 0.785 ;
        RECT  0.615 0.195 1.705 0.265 ;
        RECT  1.600 0.855 1.700 1.065 ;
        RECT  1.510 0.395 1.690 0.465 ;
        RECT  1.510 0.715 1.690 0.785 ;
        RECT  0.695 0.995 1.600 1.065 ;
        RECT  1.440 0.345 1.510 0.465 ;
        RECT  1.440 0.715 1.510 0.910 ;
        RECT  1.370 0.545 1.440 0.615 ;
        RECT  1.300 0.355 1.370 0.925 ;
        RECT  1.010 0.355 1.300 0.425 ;
        RECT  0.990 0.855 1.300 0.925 ;
        RECT  0.410 0.355 0.930 0.425 ;
        RECT  0.385 0.535 0.795 0.605 ;
        RECT  0.625 0.925 0.695 1.065 ;
        RECT  0.340 0.535 0.385 0.940 ;
        RECT  0.270 0.355 0.340 0.940 ;
        RECT  0.125 0.355 0.270 0.425 ;
        RECT  0.125 0.870 0.270 0.940 ;
        RECT  0.055 0.305 0.125 0.425 ;
        RECT  0.055 0.870 0.125 1.075 ;
    END
END DFKCSNQD2BWP40

MACRO DFKCSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFKCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.190 0.675 ;
        RECT  0.035 0.495 0.130 0.770 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.705 0.205 4.795 0.470 ;
        RECT  4.705 0.685 4.795 1.075 ;
        RECT  4.655 0.385 4.705 0.470 ;
        RECT  4.655 0.685 4.705 0.770 ;
        RECT  4.445 0.385 4.655 0.770 ;
        RECT  4.435 0.385 4.445 0.470 ;
        RECT  4.435 0.685 4.445 0.770 ;
        RECT  4.345 0.205 4.435 0.470 ;
        RECT  4.345 0.685 4.435 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.680 0.575 0.800 ;
        RECT  0.455 0.680 0.545 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.225 0.765 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.985 0.765 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.990 0.445 ;
        RECT  4.605 -0.115 4.915 0.115 ;
        RECT  4.535 -0.115 4.605 0.255 ;
        RECT  4.225 -0.115 4.535 0.115 ;
        RECT  4.155 -0.115 4.225 0.305 ;
        RECT  3.845 -0.115 4.155 0.115 ;
        RECT  3.775 -0.115 3.845 0.305 ;
        RECT  3.060 -0.115 3.775 0.115 ;
        RECT  2.980 -0.115 3.060 0.445 ;
        RECT  2.670 -0.115 2.980 0.115 ;
        RECT  2.590 -0.115 2.670 0.445 ;
        RECT  2.300 -0.115 2.590 0.115 ;
        RECT  2.180 -0.115 2.300 0.210 ;
        RECT  1.300 -0.115 2.180 0.115 ;
        RECT  1.180 -0.115 1.300 0.125 ;
        RECT  0.320 -0.115 1.180 0.115 ;
        RECT  0.200 -0.115 0.320 0.125 ;
        RECT  0.000 -0.115 0.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.915 0.715 4.990 1.375 ;
        RECT  4.605 1.145 4.915 1.375 ;
        RECT  4.535 0.885 4.605 1.375 ;
        RECT  4.245 1.145 4.535 1.375 ;
        RECT  4.135 0.970 4.245 1.375 ;
        RECT  3.850 1.145 4.135 1.375 ;
        RECT  3.780 0.695 3.850 1.375 ;
        RECT  3.060 1.145 3.780 1.375 ;
        RECT  2.980 0.810 3.060 1.375 ;
        RECT  2.670 1.145 2.980 1.375 ;
        RECT  2.590 0.795 2.670 1.375 ;
        RECT  2.275 1.145 2.590 1.375 ;
        RECT  2.205 0.865 2.275 1.375 ;
        RECT  1.300 1.145 2.205 1.375 ;
        RECT  1.180 1.135 1.300 1.375 ;
        RECT  0.950 1.145 1.180 1.375 ;
        RECT  0.830 1.135 0.950 1.375 ;
        RECT  0.340 1.145 0.830 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.205 4.795 0.470 ;
        RECT  4.725 0.685 4.795 1.075 ;
        RECT  4.345 0.205 4.375 0.470 ;
        RECT  4.345 0.685 4.375 1.075 ;
        RECT  4.265 0.545 4.325 0.615 ;
        RECT  4.195 0.395 4.265 0.820 ;
        RECT  4.035 0.395 4.195 0.465 ;
        RECT  4.035 0.750 4.195 0.820 ;
        RECT  3.710 0.545 4.055 0.615 ;
        RECT  3.965 0.185 4.035 0.465 ;
        RECT  3.965 0.750 4.035 1.075 ;
        RECT  3.635 0.395 3.965 0.465 ;
        RECT  3.640 0.545 3.710 1.060 ;
        RECT  3.530 0.545 3.640 0.615 ;
        RECT  3.350 0.990 3.640 1.060 ;
        RECT  3.490 0.800 3.560 0.920 ;
        RECT  3.460 0.240 3.530 0.615 ;
        RECT  3.390 0.800 3.490 0.870 ;
        RECT  3.350 0.240 3.460 0.310 ;
        RECT  3.320 0.430 3.390 0.870 ;
        RECT  3.180 0.215 3.250 0.585 ;
        RECT  3.175 0.665 3.250 1.065 ;
        RECT  2.860 0.515 3.180 0.585 ;
        RECT  2.860 0.665 3.175 0.740 ;
        RECT  2.780 0.335 2.860 0.585 ;
        RECT  2.780 0.665 2.860 0.910 ;
        RECT  2.410 0.300 2.480 0.980 ;
        RECT  2.395 0.300 2.410 0.415 ;
        RECT  2.395 0.720 2.410 0.980 ;
        RECT  2.205 0.720 2.395 0.790 ;
        RECT  2.325 0.470 2.340 0.590 ;
        RECT  2.255 0.280 2.325 0.590 ;
        RECT  1.900 0.280 2.255 0.350 ;
        RECT  2.135 0.670 2.205 0.790 ;
        RECT  2.045 0.885 2.105 0.955 ;
        RECT  2.045 0.420 2.100 0.490 ;
        RECT  1.975 0.420 2.045 0.955 ;
        RECT  1.830 0.195 1.900 0.960 ;
        RECT  1.785 0.195 1.830 0.265 ;
        RECT  1.690 0.395 1.760 0.785 ;
        RECT  0.615 0.195 1.705 0.265 ;
        RECT  1.600 0.855 1.700 1.065 ;
        RECT  1.510 0.395 1.690 0.465 ;
        RECT  1.510 0.715 1.690 0.785 ;
        RECT  0.695 0.995 1.600 1.065 ;
        RECT  1.440 0.345 1.510 0.465 ;
        RECT  1.440 0.715 1.510 0.910 ;
        RECT  1.370 0.545 1.440 0.615 ;
        RECT  1.300 0.355 1.370 0.925 ;
        RECT  1.010 0.355 1.300 0.425 ;
        RECT  0.990 0.855 1.300 0.925 ;
        RECT  0.410 0.355 0.930 0.425 ;
        RECT  0.385 0.535 0.795 0.605 ;
        RECT  0.625 0.925 0.695 1.065 ;
        RECT  0.340 0.535 0.385 0.940 ;
        RECT  0.270 0.355 0.340 0.940 ;
        RECT  0.125 0.355 0.270 0.425 ;
        RECT  0.125 0.870 0.270 0.940 ;
        RECT  0.055 0.305 0.125 0.425 ;
        RECT  0.055 0.870 0.125 1.075 ;
    END
END DFKCSNQD4BWP40

MACRO DFKSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFKSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.735 0.765 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.050000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.195 3.885 1.060 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 -0.115 3.920 0.115 ;
        RECT  3.570 -0.115 3.690 0.260 ;
        RECT  3.275 -0.115 3.570 0.115 ;
        RECT  3.205 -0.115 3.275 0.305 ;
        RECT  2.590 -0.115 3.205 0.115 ;
        RECT  2.460 -0.115 2.590 0.120 ;
        RECT  2.160 -0.115 2.460 0.115 ;
        RECT  2.040 -0.115 2.160 0.120 ;
        RECT  1.305 -0.115 2.040 0.115 ;
        RECT  1.185 -0.115 1.305 0.120 ;
        RECT  0.950 -0.115 1.185 0.115 ;
        RECT  0.830 -0.115 0.950 0.120 ;
        RECT  0.345 -0.115 0.830 0.115 ;
        RECT  0.220 -0.115 0.345 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.665 1.145 3.920 1.375 ;
        RECT  3.595 0.945 3.665 1.375 ;
        RECT  3.290 1.145 3.595 1.375 ;
        RECT  3.220 0.950 3.290 1.375 ;
        RECT  2.540 1.145 3.220 1.375 ;
        RECT  2.465 0.775 2.540 1.375 ;
        RECT  2.150 1.145 2.465 1.375 ;
        RECT  2.080 0.840 2.150 1.375 ;
        RECT  0.930 1.145 2.080 1.375 ;
        RECT  0.810 1.140 0.930 1.375 ;
        RECT  0.370 1.145 0.810 1.375 ;
        RECT  0.250 1.140 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.375 3.720 0.805 ;
        RECT  3.465 0.375 3.650 0.445 ;
        RECT  3.470 0.735 3.650 0.805 ;
        RECT  3.330 0.545 3.570 0.615 ;
        RECT  3.400 0.735 3.470 1.065 ;
        RECT  3.395 0.195 3.465 0.445 ;
        RECT  3.185 0.375 3.395 0.445 ;
        RECT  3.260 0.545 3.330 0.805 ;
        RECT  3.150 0.735 3.260 0.805 ;
        RECT  3.115 0.375 3.185 0.640 ;
        RECT  3.080 0.735 3.150 1.055 ;
        RECT  2.850 0.985 3.080 1.055 ;
        RECT  3.005 0.195 3.035 0.620 ;
        RECT  2.965 0.195 3.005 0.905 ;
        RECT  2.835 0.195 2.965 0.265 ;
        RECT  2.935 0.550 2.965 0.905 ;
        RECT  2.850 0.350 2.895 0.470 ;
        RECT  2.780 0.350 2.850 1.055 ;
        RECT  2.705 0.185 2.835 0.265 ;
        RECT  0.505 0.195 2.705 0.265 ;
        RECT  2.295 0.355 2.365 0.950 ;
        RECT  2.285 0.355 2.295 0.465 ;
        RECT  2.285 0.700 2.295 0.950 ;
        RECT  2.055 0.700 2.285 0.770 ;
        RECT  2.205 0.510 2.225 0.630 ;
        RECT  2.135 0.355 2.205 0.630 ;
        RECT  1.750 0.355 2.135 0.425 ;
        RECT  1.985 0.655 2.055 0.770 ;
        RECT  1.890 0.840 1.985 0.910 ;
        RECT  1.890 0.495 1.940 0.565 ;
        RECT  1.785 0.995 1.905 1.075 ;
        RECT  1.820 0.495 1.890 0.910 ;
        RECT  0.340 0.995 1.785 1.065 ;
        RECT  1.680 0.355 1.750 0.905 ;
        RECT  1.600 0.355 1.680 0.425 ;
        RECT  1.200 0.835 1.565 0.905 ;
        RECT  1.010 0.350 1.505 0.420 ;
        RECT  0.930 0.520 0.950 0.640 ;
        RECT  0.860 0.335 0.930 0.925 ;
        RECT  0.590 0.335 0.860 0.405 ;
        RECT  0.590 0.855 0.860 0.925 ;
        RECT  0.435 0.195 0.505 0.915 ;
        RECT  0.270 0.345 0.340 1.065 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.055 0.835 0.270 0.950 ;
        RECT  0.055 0.195 0.125 0.415 ;
    END
END DFKSNQD0BWP40

MACRO DFKSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFKSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.735 0.765 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.100000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.185 3.885 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 -0.115 3.920 0.115 ;
        RECT  3.570 -0.115 3.690 0.280 ;
        RECT  3.275 -0.115 3.570 0.115 ;
        RECT  3.205 -0.115 3.275 0.305 ;
        RECT  2.580 -0.115 3.205 0.115 ;
        RECT  2.460 -0.115 2.580 0.120 ;
        RECT  2.160 -0.115 2.460 0.115 ;
        RECT  2.040 -0.115 2.160 0.120 ;
        RECT  1.305 -0.115 2.040 0.115 ;
        RECT  1.185 -0.115 1.305 0.120 ;
        RECT  0.950 -0.115 1.185 0.115 ;
        RECT  0.830 -0.115 0.950 0.120 ;
        RECT  0.345 -0.115 0.830 0.115 ;
        RECT  0.220 -0.115 0.345 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.665 1.145 3.920 1.375 ;
        RECT  3.595 0.860 3.665 1.375 ;
        RECT  3.285 1.145 3.595 1.375 ;
        RECT  3.215 0.950 3.285 1.375 ;
        RECT  2.545 1.145 3.215 1.375 ;
        RECT  2.470 0.685 2.545 1.375 ;
        RECT  2.150 1.145 2.470 1.375 ;
        RECT  2.080 0.840 2.150 1.375 ;
        RECT  0.890 1.145 2.080 1.375 ;
        RECT  0.770 1.140 0.890 1.375 ;
        RECT  0.370 1.145 0.770 1.375 ;
        RECT  0.250 1.140 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.375 3.720 0.765 ;
        RECT  3.465 0.375 3.650 0.445 ;
        RECT  3.470 0.695 3.650 0.765 ;
        RECT  3.330 0.545 3.555 0.615 ;
        RECT  3.400 0.695 3.470 1.000 ;
        RECT  3.395 0.195 3.465 0.445 ;
        RECT  3.190 0.375 3.395 0.445 ;
        RECT  3.260 0.545 3.330 0.805 ;
        RECT  3.140 0.735 3.260 0.805 ;
        RECT  3.110 0.375 3.190 0.640 ;
        RECT  3.070 0.735 3.140 1.060 ;
        RECT  2.850 0.990 3.070 1.060 ;
        RECT  3.000 0.195 3.035 0.620 ;
        RECT  2.965 0.195 3.000 0.910 ;
        RECT  2.835 0.195 2.965 0.265 ;
        RECT  2.930 0.550 2.965 0.910 ;
        RECT  2.850 0.350 2.895 0.470 ;
        RECT  2.780 0.350 2.850 1.060 ;
        RECT  2.705 0.185 2.835 0.265 ;
        RECT  0.505 0.195 2.705 0.265 ;
        RECT  2.355 0.375 2.395 0.770 ;
        RECT  2.325 0.375 2.355 0.950 ;
        RECT  2.285 0.375 2.325 0.485 ;
        RECT  2.285 0.700 2.325 0.950 ;
        RECT  2.040 0.700 2.285 0.770 ;
        RECT  2.205 0.550 2.255 0.620 ;
        RECT  2.135 0.335 2.205 0.620 ;
        RECT  1.750 0.335 2.135 0.405 ;
        RECT  1.970 0.650 2.040 0.770 ;
        RECT  1.890 0.840 1.985 0.910 ;
        RECT  1.890 0.475 1.940 0.545 ;
        RECT  1.785 0.995 1.905 1.075 ;
        RECT  1.820 0.475 1.890 0.910 ;
        RECT  0.340 0.995 1.785 1.065 ;
        RECT  1.680 0.335 1.750 0.905 ;
        RECT  1.610 0.335 1.680 0.445 ;
        RECT  1.205 0.835 1.560 0.905 ;
        RECT  1.010 0.335 1.505 0.405 ;
        RECT  0.930 0.520 0.950 0.640 ;
        RECT  0.860 0.335 0.930 0.925 ;
        RECT  0.590 0.335 0.860 0.405 ;
        RECT  0.590 0.855 0.860 0.925 ;
        RECT  0.435 0.195 0.505 0.915 ;
        RECT  0.270 0.345 0.340 1.065 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.055 0.835 0.270 0.950 ;
        RECT  0.055 0.195 0.125 0.415 ;
    END
END DFKSNQD1BWP40

MACRO DFKSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFKSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.735 0.765 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.805 0.185 3.895 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.115 4.200 0.115 ;
        RECT  4.055 -0.115 4.125 0.450 ;
        RECT  3.690 -0.115 4.055 0.115 ;
        RECT  3.570 -0.115 3.690 0.280 ;
        RECT  3.275 -0.115 3.570 0.115 ;
        RECT  3.205 -0.115 3.275 0.305 ;
        RECT  2.580 -0.115 3.205 0.115 ;
        RECT  2.460 -0.115 2.580 0.120 ;
        RECT  2.160 -0.115 2.460 0.115 ;
        RECT  2.040 -0.115 2.160 0.120 ;
        RECT  1.305 -0.115 2.040 0.115 ;
        RECT  1.185 -0.115 1.305 0.120 ;
        RECT  0.950 -0.115 1.185 0.115 ;
        RECT  0.830 -0.115 0.950 0.120 ;
        RECT  0.345 -0.115 0.830 0.115 ;
        RECT  0.220 -0.115 0.345 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.145 4.200 1.375 ;
        RECT  4.055 0.710 4.125 1.375 ;
        RECT  3.665 1.145 4.055 1.375 ;
        RECT  3.595 0.860 3.665 1.375 ;
        RECT  3.285 1.145 3.595 1.375 ;
        RECT  3.215 0.950 3.285 1.375 ;
        RECT  2.545 1.145 3.215 1.375 ;
        RECT  2.470 0.685 2.545 1.375 ;
        RECT  2.150 1.145 2.470 1.375 ;
        RECT  2.080 0.840 2.150 1.375 ;
        RECT  0.890 1.145 2.080 1.375 ;
        RECT  0.770 1.140 0.890 1.375 ;
        RECT  0.370 1.145 0.770 1.375 ;
        RECT  0.250 1.140 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.665 0.375 3.735 0.765 ;
        RECT  3.465 0.375 3.665 0.445 ;
        RECT  3.470 0.695 3.665 0.765 ;
        RECT  3.330 0.545 3.555 0.615 ;
        RECT  3.400 0.695 3.470 1.000 ;
        RECT  3.395 0.195 3.465 0.445 ;
        RECT  3.190 0.375 3.395 0.445 ;
        RECT  3.260 0.545 3.330 0.805 ;
        RECT  3.140 0.735 3.260 0.805 ;
        RECT  3.110 0.375 3.190 0.640 ;
        RECT  3.070 0.735 3.140 1.060 ;
        RECT  2.850 0.990 3.070 1.060 ;
        RECT  3.000 0.195 3.035 0.620 ;
        RECT  2.965 0.195 3.000 0.910 ;
        RECT  2.835 0.195 2.965 0.265 ;
        RECT  2.930 0.550 2.965 0.910 ;
        RECT  2.850 0.350 2.895 0.470 ;
        RECT  2.780 0.350 2.850 1.060 ;
        RECT  2.705 0.185 2.835 0.265 ;
        RECT  0.505 0.195 2.705 0.265 ;
        RECT  2.355 0.375 2.395 0.770 ;
        RECT  2.325 0.375 2.355 0.950 ;
        RECT  2.285 0.375 2.325 0.485 ;
        RECT  2.285 0.700 2.325 0.950 ;
        RECT  2.040 0.700 2.285 0.770 ;
        RECT  2.205 0.550 2.255 0.620 ;
        RECT  2.135 0.335 2.205 0.620 ;
        RECT  1.750 0.335 2.135 0.405 ;
        RECT  1.970 0.650 2.040 0.770 ;
        RECT  1.890 0.840 1.985 0.910 ;
        RECT  1.890 0.475 1.940 0.545 ;
        RECT  1.785 0.995 1.905 1.075 ;
        RECT  1.820 0.475 1.890 0.910 ;
        RECT  0.340 0.995 1.785 1.065 ;
        RECT  1.680 0.335 1.750 0.905 ;
        RECT  1.610 0.335 1.680 0.445 ;
        RECT  1.205 0.835 1.560 0.905 ;
        RECT  1.010 0.335 1.505 0.405 ;
        RECT  0.930 0.520 0.950 0.640 ;
        RECT  0.860 0.335 0.930 0.925 ;
        RECT  0.590 0.335 0.860 0.405 ;
        RECT  0.590 0.855 0.860 0.925 ;
        RECT  0.435 0.195 0.505 0.915 ;
        RECT  0.270 0.345 0.340 1.065 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.055 0.835 0.270 0.950 ;
        RECT  0.055 0.195 0.125 0.415 ;
    END
END DFKSNQD2BWP40

MACRO DFKSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFKSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.735 0.765 ;
        END
    END SN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.425 0.205 4.515 0.470 ;
        RECT  4.425 0.685 4.515 1.075 ;
        RECT  4.375 0.385 4.425 0.470 ;
        RECT  4.375 0.685 4.425 0.770 ;
        RECT  4.165 0.385 4.375 0.770 ;
        RECT  4.155 0.385 4.165 0.470 ;
        RECT  4.155 0.685 4.165 0.770 ;
        RECT  4.065 0.210 4.155 0.470 ;
        RECT  4.065 0.685 4.155 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.365 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.635 -0.115 4.710 0.445 ;
        RECT  4.325 -0.115 4.635 0.115 ;
        RECT  4.255 -0.115 4.325 0.255 ;
        RECT  3.925 -0.115 4.255 0.115 ;
        RECT  3.855 -0.115 3.925 0.265 ;
        RECT  3.520 -0.115 3.855 0.115 ;
        RECT  3.450 -0.115 3.520 0.265 ;
        RECT  3.340 -0.115 3.450 0.115 ;
        RECT  3.270 -0.115 3.340 0.400 ;
        RECT  2.540 -0.115 3.270 0.115 ;
        RECT  2.420 -0.115 2.540 0.120 ;
        RECT  2.160 -0.115 2.420 0.115 ;
        RECT  2.040 -0.115 2.160 0.120 ;
        RECT  1.305 -0.115 2.040 0.115 ;
        RECT  1.185 -0.115 1.305 0.120 ;
        RECT  0.950 -0.115 1.185 0.115 ;
        RECT  0.830 -0.115 0.950 0.120 ;
        RECT  0.345 -0.115 0.830 0.115 ;
        RECT  0.220 -0.115 0.345 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.635 0.715 4.710 1.375 ;
        RECT  4.325 1.145 4.635 1.375 ;
        RECT  4.255 0.885 4.325 1.375 ;
        RECT  3.925 1.145 4.255 1.375 ;
        RECT  3.855 1.020 3.925 1.375 ;
        RECT  3.520 1.145 3.855 1.375 ;
        RECT  3.450 0.865 3.520 1.375 ;
        RECT  3.345 1.145 3.450 1.375 ;
        RECT  3.275 0.835 3.345 1.375 ;
        RECT  2.535 1.145 3.275 1.375 ;
        RECT  2.465 0.685 2.535 1.375 ;
        RECT  2.150 1.145 2.465 1.375 ;
        RECT  2.080 0.840 2.150 1.375 ;
        RECT  0.890 1.145 2.080 1.375 ;
        RECT  0.770 1.140 0.890 1.375 ;
        RECT  0.370 1.145 0.770 1.375 ;
        RECT  0.250 1.140 0.370 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.205 4.515 0.470 ;
        RECT  4.445 0.685 4.515 1.075 ;
        RECT  4.065 0.210 4.095 0.470 ;
        RECT  4.065 0.685 4.095 1.075 ;
        RECT  3.995 0.545 4.035 0.615 ;
        RECT  3.925 0.365 3.995 0.895 ;
        RECT  3.710 0.365 3.925 0.435 ;
        RECT  3.710 0.825 3.925 0.895 ;
        RECT  3.640 0.205 3.710 0.435 ;
        RECT  3.640 0.525 3.710 0.755 ;
        RECT  3.640 0.825 3.710 1.075 ;
        RECT  3.490 0.365 3.640 0.435 ;
        RECT  3.205 0.685 3.640 0.755 ;
        RECT  3.420 0.365 3.490 0.575 ;
        RECT  3.250 0.505 3.420 0.575 ;
        RECT  3.180 0.505 3.250 0.615 ;
        RECT  3.135 0.685 3.205 1.015 ;
        RECT  2.915 0.945 3.135 1.015 ;
        RECT  3.065 0.195 3.100 0.620 ;
        RECT  3.030 0.195 3.065 0.795 ;
        RECT  0.505 0.195 3.030 0.265 ;
        RECT  2.995 0.550 3.030 0.795 ;
        RECT  2.915 0.350 2.960 0.470 ;
        RECT  2.845 0.350 2.915 1.015 ;
        RECT  2.355 0.375 2.395 0.770 ;
        RECT  2.325 0.375 2.355 0.950 ;
        RECT  2.285 0.375 2.325 0.485 ;
        RECT  2.285 0.700 2.325 0.950 ;
        RECT  2.040 0.700 2.285 0.770 ;
        RECT  2.205 0.550 2.255 0.620 ;
        RECT  2.135 0.335 2.205 0.620 ;
        RECT  1.750 0.335 2.135 0.405 ;
        RECT  1.970 0.650 2.040 0.770 ;
        RECT  1.890 0.840 1.985 0.910 ;
        RECT  1.890 0.475 1.940 0.545 ;
        RECT  1.785 0.995 1.905 1.075 ;
        RECT  1.820 0.475 1.890 0.910 ;
        RECT  0.340 0.995 1.785 1.065 ;
        RECT  1.680 0.335 1.750 0.905 ;
        RECT  1.610 0.335 1.680 0.445 ;
        RECT  1.205 0.835 1.560 0.905 ;
        RECT  1.010 0.335 1.505 0.405 ;
        RECT  0.930 0.520 0.950 0.640 ;
        RECT  0.860 0.335 0.930 0.925 ;
        RECT  0.590 0.335 0.860 0.405 ;
        RECT  0.590 0.855 0.860 0.925 ;
        RECT  0.435 0.195 0.505 0.915 ;
        RECT  0.270 0.345 0.340 1.065 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.055 0.835 0.270 0.950 ;
        RECT  0.055 0.195 0.125 0.415 ;
    END
END DFKSNQD4BWP40

MACRO DFMQD0BWP40
    CLASS CORE ;
    FOREIGN DFMQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.640 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.045 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.895 0.635 1.015 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.675 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.705 -0.115 3.375 0.115 ;
        RECT  2.560 -0.115 2.705 0.125 ;
        RECT  2.035 -0.115 2.560 0.115 ;
        RECT  1.915 -0.115 2.035 0.125 ;
        RECT  1.120 -0.115 1.915 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.250 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.660 1.145 3.310 1.375 ;
        RECT  2.540 0.970 2.660 1.375 ;
        RECT  2.050 1.145 2.540 1.375 ;
        RECT  1.930 0.805 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.810 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.740 3.775 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.960 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.005 0.860 3.415 0.930 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.115 0.195 3.185 0.780 ;
        RECT  2.940 0.195 3.115 0.265 ;
        RECT  2.935 0.350 3.005 0.930 ;
        RECT  2.830 0.185 2.940 0.265 ;
        RECT  2.915 0.350 2.935 0.470 ;
        RECT  2.810 0.185 2.830 0.875 ;
        RECT  2.760 0.195 2.810 0.875 ;
        RECT  1.660 0.195 2.760 0.265 ;
        RECT  2.440 0.785 2.760 0.875 ;
        RECT  2.290 0.520 2.690 0.640 ;
        RECT  2.360 0.785 2.440 0.995 ;
        RECT  2.150 0.335 2.220 0.900 ;
        RECT  1.890 0.540 2.150 0.660 ;
        RECT  1.820 0.370 1.860 0.460 ;
        RECT  1.740 0.370 1.820 0.925 ;
        RECT  1.660 0.995 1.760 1.065 ;
        RECT  1.590 0.845 1.660 1.065 ;
        RECT  1.575 0.350 1.645 0.765 ;
        RECT  1.450 0.845 1.590 0.915 ;
        RECT  1.530 0.690 1.575 0.765 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  0.590 0.985 1.460 1.055 ;
        RECT  1.380 0.345 1.450 0.915 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.145 0.845 1.380 0.915 ;
        RECT  0.815 0.845 0.910 0.915 ;
        RECT  0.820 0.335 0.890 0.525 ;
        RECT  0.815 0.455 0.820 0.525 ;
        RECT  0.745 0.455 0.815 0.915 ;
        RECT  0.540 0.695 0.620 0.915 ;
        RECT  0.140 0.845 0.540 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.395 0.525 2.465 0.595 ;
        RECT  1.575 0.525 1.645 0.595 ;
        LAYER M2 ;
        RECT  1.525 0.525 2.515 0.595 ;
    END
END DFMQD0BWP40

MACRO DFMQD1BWP40
    CLASS CORE ;
    FOREIGN DFMQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.640 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.895 0.635 1.015 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.675 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.715 -0.115 3.375 0.115 ;
        RECT  2.570 -0.115 2.715 0.125 ;
        RECT  2.025 -0.115 2.570 0.115 ;
        RECT  1.905 -0.115 2.025 0.125 ;
        RECT  1.120 -0.115 1.905 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.250 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.660 1.145 3.310 1.375 ;
        RECT  2.540 0.970 2.660 1.375 ;
        RECT  2.055 1.145 2.540 1.375 ;
        RECT  1.935 0.730 2.055 1.375 ;
        RECT  1.120 1.145 1.935 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.810 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.740 3.775 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.960 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.015 0.860 3.415 0.930 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.115 0.195 3.185 0.780 ;
        RECT  2.940 0.195 3.115 0.265 ;
        RECT  2.945 0.350 3.015 0.930 ;
        RECT  2.910 0.350 2.945 0.470 ;
        RECT  2.840 0.185 2.940 0.265 ;
        RECT  2.810 0.185 2.840 0.875 ;
        RECT  2.770 0.195 2.810 0.875 ;
        RECT  1.650 0.195 2.770 0.265 ;
        RECT  2.450 0.785 2.770 0.875 ;
        RECT  2.290 0.520 2.690 0.640 ;
        RECT  2.355 0.785 2.450 1.015 ;
        RECT  2.150 0.335 2.220 0.950 ;
        RECT  1.890 0.530 2.150 0.650 ;
        RECT  1.750 0.345 1.820 0.925 ;
        RECT  1.640 0.995 1.765 1.065 ;
        RECT  1.635 0.690 1.655 0.765 ;
        RECT  1.570 0.845 1.640 1.065 ;
        RECT  1.565 0.350 1.635 0.765 ;
        RECT  1.450 0.845 1.570 0.915 ;
        RECT  1.545 0.690 1.565 0.765 ;
        RECT  0.585 0.195 1.480 0.265 ;
        RECT  0.605 0.985 1.465 1.055 ;
        RECT  1.380 0.345 1.450 0.915 ;
        RECT  1.160 0.345 1.380 0.415 ;
        RECT  1.155 0.845 1.380 0.915 ;
        RECT  0.815 0.845 0.910 0.915 ;
        RECT  0.820 0.335 0.890 0.525 ;
        RECT  0.815 0.455 0.820 0.525 ;
        RECT  0.745 0.455 0.815 0.915 ;
        RECT  0.540 0.695 0.620 0.915 ;
        RECT  0.140 0.845 0.540 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.385 0.525 2.455 0.595 ;
        RECT  1.565 0.525 1.635 0.595 ;
        LAYER M2 ;
        RECT  1.515 0.525 2.505 0.595 ;
    END
END DFMQD1BWP40

MACRO DFMQD2BWP40
    CLASS CORE ;
    FOREIGN DFMQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.640 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.195 4.035 1.075 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.895 0.635 1.015 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.675 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.250 -0.115 4.340 0.115 ;
        RECT  4.180 -0.115 4.250 0.495 ;
        RECT  3.815 -0.115 4.180 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.715 -0.115 3.375 0.115 ;
        RECT  2.570 -0.115 2.715 0.125 ;
        RECT  2.025 -0.115 2.570 0.115 ;
        RECT  1.905 -0.115 2.025 0.125 ;
        RECT  1.120 -0.115 1.905 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.250 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.145 4.340 1.375 ;
        RECT  4.180 0.700 4.250 1.375 ;
        RECT  3.815 1.145 4.180 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.660 1.145 3.310 1.375 ;
        RECT  2.540 0.970 2.660 1.375 ;
        RECT  2.055 1.145 2.540 1.375 ;
        RECT  1.935 0.730 2.055 1.375 ;
        RECT  1.120 1.145 1.935 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.810 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.740 3.785 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.960 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.015 0.860 3.415 0.930 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.115 0.195 3.185 0.780 ;
        RECT  2.940 0.195 3.115 0.265 ;
        RECT  2.945 0.350 3.015 0.930 ;
        RECT  2.910 0.350 2.945 0.470 ;
        RECT  2.840 0.185 2.940 0.265 ;
        RECT  2.810 0.185 2.840 0.875 ;
        RECT  2.770 0.195 2.810 0.875 ;
        RECT  1.650 0.195 2.770 0.265 ;
        RECT  2.455 0.785 2.770 0.875 ;
        RECT  2.290 0.520 2.690 0.640 ;
        RECT  2.355 0.785 2.455 1.045 ;
        RECT  2.150 0.335 2.220 0.955 ;
        RECT  1.890 0.530 2.150 0.650 ;
        RECT  1.745 0.350 1.820 0.925 ;
        RECT  1.660 0.995 1.765 1.065 ;
        RECT  1.590 0.845 1.660 1.065 ;
        RECT  1.635 0.690 1.655 0.765 ;
        RECT  1.565 0.350 1.635 0.765 ;
        RECT  1.450 0.845 1.590 0.915 ;
        RECT  1.545 0.690 1.565 0.765 ;
        RECT  0.585 0.195 1.480 0.265 ;
        RECT  0.605 0.985 1.465 1.055 ;
        RECT  1.380 0.345 1.450 0.915 ;
        RECT  1.160 0.345 1.380 0.415 ;
        RECT  1.155 0.845 1.380 0.915 ;
        RECT  0.815 0.845 0.910 0.915 ;
        RECT  0.820 0.335 0.890 0.525 ;
        RECT  0.815 0.455 0.820 0.525 ;
        RECT  0.745 0.455 0.815 0.915 ;
        RECT  0.540 0.695 0.620 0.915 ;
        RECT  0.140 0.845 0.540 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.365 0.525 2.435 0.595 ;
        RECT  1.565 0.525 1.635 0.595 ;
        LAYER M2 ;
        RECT  1.515 0.525 2.485 0.595 ;
    END
END DFMQD2BWP40

MACRO DFMQD4BWP40
    CLASS CORE ;
    FOREIGN DFMQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SA
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.640 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.865 0.195 4.960 0.440 ;
        RECT  4.865 0.745 4.960 0.995 ;
        RECT  4.795 0.355 4.865 0.440 ;
        RECT  4.795 0.745 4.865 0.830 ;
        RECT  4.585 0.355 4.795 0.830 ;
        RECT  4.560 0.355 4.585 0.485 ;
        RECT  4.565 0.705 4.585 0.830 ;
        RECT  4.490 0.705 4.565 0.995 ;
        RECT  4.490 0.210 4.560 0.485 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.895 0.635 1.015 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.675 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.115 5.180 0.115 ;
        RECT  5.050 -0.115 5.125 0.445 ;
        RECT  4.750 -0.115 5.050 0.115 ;
        RECT  4.670 -0.115 4.750 0.265 ;
        RECT  4.365 -0.115 4.670 0.115 ;
        RECT  4.295 -0.115 4.365 0.315 ;
        RECT  3.995 -0.115 4.295 0.115 ;
        RECT  3.925 -0.115 3.995 0.315 ;
        RECT  3.160 -0.115 3.925 0.115 ;
        RECT  3.040 -0.115 3.160 0.125 ;
        RECT  2.735 -0.115 3.040 0.115 ;
        RECT  2.605 -0.115 2.735 0.125 ;
        RECT  2.040 -0.115 2.605 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.120 -0.115 1.920 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.250 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.145 5.180 1.375 ;
        RECT  5.050 0.700 5.125 1.375 ;
        RECT  4.765 1.145 5.050 1.375 ;
        RECT  4.655 0.905 4.765 1.375 ;
        RECT  4.390 1.145 4.655 1.375 ;
        RECT  4.275 0.880 4.390 1.375 ;
        RECT  4.000 1.145 4.275 1.375 ;
        RECT  3.870 1.130 4.000 1.375 ;
        RECT  3.180 1.145 3.870 1.375 ;
        RECT  3.060 1.010 3.180 1.375 ;
        RECT  2.750 1.145 3.060 1.375 ;
        RECT  2.630 0.900 2.750 1.375 ;
        RECT  2.090 1.145 2.630 1.375 ;
        RECT  1.965 0.730 2.090 1.375 ;
        RECT  1.120 1.145 1.965 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.195 4.960 0.440 ;
        RECT  4.865 0.745 4.960 0.995 ;
        RECT  4.490 0.210 4.515 0.485 ;
        RECT  4.490 0.705 4.515 0.995 ;
        RECT  4.350 0.395 4.420 0.810 ;
        RECT  4.185 0.395 4.350 0.465 ;
        RECT  4.185 0.740 4.350 0.810 ;
        RECT  4.115 0.195 4.185 0.465 ;
        RECT  4.115 0.740 4.185 0.980 ;
        RECT  4.035 0.545 4.135 0.615 ;
        RECT  3.885 0.395 4.115 0.465 ;
        RECT  3.965 0.545 4.035 0.930 ;
        RECT  3.565 0.860 3.965 0.930 ;
        RECT  3.815 0.395 3.885 0.600 ;
        RECT  3.665 0.195 3.745 0.780 ;
        RECT  3.425 0.195 3.665 0.265 ;
        RECT  3.495 0.350 3.565 0.930 ;
        RECT  3.355 0.195 3.425 0.625 ;
        RECT  2.830 0.850 3.400 0.920 ;
        RECT  1.700 0.195 3.355 0.265 ;
        RECT  3.190 0.555 3.355 0.625 ;
        RECT  3.215 0.345 3.285 0.465 ;
        RECT  2.830 0.345 3.215 0.420 ;
        RECT  3.110 0.555 3.190 0.780 ;
        RECT  2.505 0.710 3.110 0.780 ;
        RECT  2.345 0.510 2.935 0.630 ;
        RECT  2.415 0.710 2.505 1.000 ;
        RECT  2.185 0.335 2.255 0.945 ;
        RECT  1.920 0.530 2.185 0.650 ;
        RECT  1.840 0.370 1.905 0.450 ;
        RECT  1.760 0.370 1.840 0.925 ;
        RECT  1.665 0.995 1.765 1.065 ;
        RECT  1.595 0.350 1.685 0.760 ;
        RECT  1.595 0.845 1.665 1.065 ;
        RECT  1.535 0.690 1.595 0.760 ;
        RECT  1.465 0.845 1.595 0.915 ;
        RECT  1.465 0.345 1.515 0.505 ;
        RECT  0.585 0.195 1.480 0.265 ;
        RECT  1.395 0.345 1.465 0.915 ;
        RECT  0.605 0.985 1.465 1.055 ;
        RECT  1.160 0.345 1.395 0.415 ;
        RECT  1.155 0.845 1.395 0.915 ;
        RECT  0.815 0.845 0.910 0.915 ;
        RECT  0.820 0.335 0.890 0.525 ;
        RECT  0.815 0.455 0.820 0.525 ;
        RECT  0.745 0.455 0.815 0.915 ;
        RECT  0.540 0.695 0.620 0.915 ;
        RECT  0.140 0.845 0.540 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.490 0.525 2.560 0.595 ;
        RECT  1.615 0.525 1.685 0.595 ;
        LAYER M2 ;
        RECT  1.565 0.525 2.610 0.595 ;
    END
END DFMQD4BWP40

MACRO DFNCNQD0BWP40
    CLASS CORE ;
    FOREIGN DFNCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 1.075 ;
        RECT  3.795 0.185 3.815 0.325 ;
        RECT  3.795 0.905 3.815 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.040 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.530 0.525 3.555 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 -0.115 3.920 0.115 ;
        RECT  3.570 -0.115 3.700 0.255 ;
        RECT  3.100 -0.115 3.570 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.195 -0.115 3.025 0.115 ;
        RECT  2.075 -0.115 2.195 0.310 ;
        RECT  1.765 -0.115 2.075 0.115 ;
        RECT  1.695 -0.115 1.765 0.260 ;
        RECT  0.710 -0.115 1.695 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.250 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 1.005 3.290 1.375 ;
        RECT  3.125 1.145 3.200 1.375 ;
        RECT  3.005 0.885 3.125 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 0.940 2.335 1.375 ;
        RECT  1.640 1.145 2.225 1.375 ;
        RECT  1.520 1.070 1.640 1.375 ;
        RECT  0.730 1.145 1.520 1.375 ;
        RECT  0.610 1.055 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.040 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.935 ;
        RECT  3.285 0.325 3.655 0.395 ;
        RECT  3.475 0.865 3.655 0.935 ;
        RECT  3.395 0.495 3.550 0.765 ;
        RECT  3.390 0.865 3.475 1.000 ;
        RECT  3.300 0.865 3.390 0.935 ;
        RECT  2.715 0.530 3.315 0.600 ;
        RECT  3.230 0.710 3.300 0.935 ;
        RECT  3.205 0.195 3.285 0.395 ;
        RECT  3.005 0.710 3.230 0.780 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.715 0.600 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.250 0.390 2.320 0.850 ;
        RECT  1.890 0.390 2.250 0.460 ;
        RECT  1.490 0.780 2.250 0.850 ;
        RECT  1.820 0.545 2.165 0.615 ;
        RECT  1.350 0.930 1.845 1.000 ;
        RECT  1.750 0.330 1.820 0.615 ;
        RECT  1.585 0.330 1.750 0.400 ;
        RECT  1.560 0.480 1.680 0.700 ;
        RECT  1.515 0.215 1.585 0.400 ;
        RECT  0.795 0.215 1.515 0.285 ;
        RECT  1.420 0.620 1.490 0.850 ;
        RECT  1.280 0.355 1.350 1.000 ;
        RECT  1.225 0.355 1.280 0.430 ;
        RECT  1.140 0.510 1.210 0.985 ;
        RECT  0.870 0.905 1.140 0.985 ;
        RECT  1.000 0.705 1.070 0.825 ;
        RECT  0.795 0.705 1.000 0.775 ;
        RECT  0.800 0.885 0.870 0.985 ;
        RECT  0.345 0.885 0.800 0.955 ;
        RECT  0.725 0.215 0.795 0.775 ;
        RECT  0.555 0.215 0.625 0.805 ;
        RECT  0.415 0.215 0.555 0.285 ;
        RECT  0.415 0.735 0.555 0.805 ;
        RECT  0.345 0.525 0.385 0.645 ;
        RECT  0.275 0.345 0.345 0.955 ;
        RECT  0.130 0.345 0.275 0.415 ;
        RECT  0.125 0.885 0.275 0.955 ;
        RECT  0.055 0.190 0.130 0.415 ;
        RECT  0.055 0.885 0.125 1.045 ;
        LAYER VIA1 ;
        RECT  3.435 0.525 3.505 0.595 ;
        RECT  1.590 0.525 1.660 0.595 ;
    END
END DFNCNQD0BWP40

MACRO DFNCNQD1BWP40
    CLASS CORE ;
    FOREIGN DFNCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.795 0.185 3.885 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.040 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.525 3.540 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 -0.115 3.920 0.115 ;
        RECT  3.575 -0.115 3.700 0.255 ;
        RECT  3.100 -0.115 3.575 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.195 -0.115 3.025 0.115 ;
        RECT  2.075 -0.115 2.195 0.235 ;
        RECT  1.750 -0.115 2.075 0.115 ;
        RECT  1.680 -0.115 1.750 0.260 ;
        RECT  0.710 -0.115 1.680 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.215 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.145 3.920 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 1.005 3.290 1.375 ;
        RECT  3.125 1.145 3.200 1.375 ;
        RECT  3.005 0.895 3.125 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 0.930 2.335 1.375 ;
        RECT  1.640 1.145 2.225 1.375 ;
        RECT  1.520 1.070 1.640 1.375 ;
        RECT  0.730 1.145 1.520 1.375 ;
        RECT  0.610 1.055 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.040 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.935 ;
        RECT  3.285 0.325 3.655 0.395 ;
        RECT  3.300 0.865 3.655 0.935 ;
        RECT  3.395 0.495 3.550 0.765 ;
        RECT  2.710 0.540 3.315 0.610 ;
        RECT  3.230 0.720 3.300 0.935 ;
        RECT  3.200 0.205 3.285 0.395 ;
        RECT  2.920 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.710 0.610 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.405 0.195 2.485 1.065 ;
        RECT  2.240 0.335 2.310 0.850 ;
        RECT  1.880 0.335 2.240 0.405 ;
        RECT  1.495 0.780 2.240 0.850 ;
        RECT  1.810 0.545 2.160 0.615 ;
        RECT  1.355 0.930 1.830 1.000 ;
        RECT  1.740 0.340 1.810 0.615 ;
        RECT  1.610 0.340 1.740 0.410 ;
        RECT  1.565 0.490 1.670 0.700 ;
        RECT  1.540 0.215 1.610 0.410 ;
        RECT  0.795 0.215 1.540 0.285 ;
        RECT  1.425 0.560 1.495 0.850 ;
        RECT  1.285 0.355 1.355 1.000 ;
        RECT  1.225 0.355 1.285 0.425 ;
        RECT  1.140 0.505 1.215 0.985 ;
        RECT  1.110 0.505 1.140 0.625 ;
        RECT  0.850 0.905 1.140 0.985 ;
        RECT  1.000 0.705 1.070 0.825 ;
        RECT  0.795 0.705 1.000 0.775 ;
        RECT  0.790 0.875 0.850 0.985 ;
        RECT  0.725 0.215 0.795 0.775 ;
        RECT  0.345 0.875 0.790 0.960 ;
        RECT  0.555 0.225 0.625 0.790 ;
        RECT  0.415 0.225 0.555 0.295 ;
        RECT  0.415 0.720 0.555 0.790 ;
        RECT  0.345 0.525 0.385 0.645 ;
        RECT  0.275 0.295 0.345 0.960 ;
        RECT  0.130 0.295 0.275 0.375 ;
        RECT  0.135 0.875 0.275 0.960 ;
        RECT  0.055 0.875 0.135 1.065 ;
        RECT  0.055 0.195 0.130 0.375 ;
        LAYER VIA1 ;
        RECT  3.420 0.525 3.490 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
    END
END DFNCNQD1BWP40

MACRO DFNCNQD2BWP40
    CLASS CORE ;
    FOREIGN DFNCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.140400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.810 0.185 3.885 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.040 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.520 0.525 3.550 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.105 -0.115 4.200 0.115 ;
        RECT  4.035 -0.115 4.105 0.480 ;
        RECT  3.700 -0.115 4.035 0.115 ;
        RECT  3.575 -0.115 3.700 0.255 ;
        RECT  3.100 -0.115 3.575 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.195 -0.115 3.025 0.115 ;
        RECT  2.075 -0.115 2.195 0.315 ;
        RECT  1.750 -0.115 2.075 0.115 ;
        RECT  1.680 -0.115 1.750 0.260 ;
        RECT  0.710 -0.115 1.680 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.215 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.105 1.145 4.200 1.375 ;
        RECT  4.035 0.680 4.105 1.375 ;
        RECT  3.690 1.145 4.035 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 1.005 3.290 1.375 ;
        RECT  3.125 1.145 3.200 1.375 ;
        RECT  3.005 0.895 3.125 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 0.940 2.335 1.375 ;
        RECT  1.640 1.145 2.225 1.375 ;
        RECT  1.520 1.070 1.640 1.375 ;
        RECT  0.730 1.145 1.520 1.375 ;
        RECT  0.610 1.055 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.040 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.655 0.325 3.725 0.935 ;
        RECT  3.295 0.325 3.655 0.395 ;
        RECT  3.300 0.865 3.655 0.935 ;
        RECT  3.395 0.495 3.550 0.765 ;
        RECT  2.710 0.540 3.315 0.610 ;
        RECT  3.230 0.720 3.300 0.935 ;
        RECT  3.205 0.205 3.295 0.395 ;
        RECT  2.925 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.710 0.610 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.405 0.195 2.485 1.065 ;
        RECT  2.245 0.395 2.315 0.850 ;
        RECT  1.880 0.395 2.245 0.465 ;
        RECT  1.490 0.780 2.245 0.850 ;
        RECT  1.810 0.545 2.160 0.615 ;
        RECT  1.350 0.930 1.850 1.000 ;
        RECT  1.740 0.340 1.810 0.615 ;
        RECT  1.575 0.340 1.740 0.410 ;
        RECT  1.560 0.485 1.670 0.700 ;
        RECT  1.505 0.215 1.575 0.410 ;
        RECT  0.795 0.215 1.505 0.285 ;
        RECT  1.420 0.620 1.490 0.850 ;
        RECT  1.280 0.355 1.350 1.000 ;
        RECT  1.205 0.355 1.280 0.425 ;
        RECT  1.140 0.505 1.210 0.985 ;
        RECT  0.850 0.905 1.140 0.985 ;
        RECT  1.000 0.705 1.070 0.825 ;
        RECT  0.795 0.705 1.000 0.775 ;
        RECT  0.790 0.875 0.850 0.985 ;
        RECT  0.725 0.215 0.795 0.775 ;
        RECT  0.345 0.875 0.790 0.960 ;
        RECT  0.555 0.350 0.625 0.790 ;
        RECT  0.415 0.350 0.555 0.420 ;
        RECT  0.415 0.720 0.555 0.790 ;
        RECT  0.345 0.525 0.385 0.645 ;
        RECT  0.275 0.335 0.345 0.960 ;
        RECT  0.130 0.335 0.275 0.415 ;
        RECT  0.130 0.875 0.275 0.960 ;
        RECT  0.055 0.195 0.130 0.415 ;
        RECT  0.055 0.875 0.130 1.065 ;
        LAYER VIA1 ;
        RECT  3.430 0.525 3.500 0.595 ;
        RECT  1.580 0.525 1.650 0.595 ;
    END
END DFNCNQD2BWP40

MACRO DFNCNQD4BWP40
    CLASS CORE ;
    FOREIGN DFNCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.264900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.745 4.880 1.000 ;
        RECT  4.795 0.205 4.870 0.485 ;
        RECT  4.785 0.205 4.795 1.000 ;
        RECT  4.770 0.355 4.785 1.000 ;
        RECT  4.585 0.355 4.770 0.830 ;
        RECT  4.480 0.355 4.585 0.485 ;
        RECT  4.480 0.710 4.585 0.830 ;
        RECT  4.400 0.205 4.480 0.485 ;
        RECT  4.400 0.710 4.480 1.000 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.040 0.625 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.050600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.525 3.860 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 -0.115 5.180 0.115 ;
        RECT  5.040 -0.115 5.110 0.480 ;
        RECT  4.665 -0.115 5.040 0.115 ;
        RECT  4.590 -0.115 4.665 0.275 ;
        RECT  4.310 -0.115 4.590 0.115 ;
        RECT  4.175 -0.115 4.310 0.140 ;
        RECT  3.910 -0.115 4.175 0.115 ;
        RECT  3.775 -0.115 3.910 0.140 ;
        RECT  3.100 -0.115 3.775 0.115 ;
        RECT  3.025 -0.115 3.100 0.425 ;
        RECT  2.195 -0.115 3.025 0.115 ;
        RECT  2.075 -0.115 2.195 0.235 ;
        RECT  1.755 -0.115 2.075 0.115 ;
        RECT  1.685 -0.115 1.755 0.260 ;
        RECT  0.710 -0.115 1.685 0.115 ;
        RECT  0.590 -0.115 0.710 0.145 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.145 5.180 1.375 ;
        RECT  5.040 0.705 5.110 1.375 ;
        RECT  4.660 1.145 5.040 1.375 ;
        RECT  4.590 0.960 4.660 1.375 ;
        RECT  4.280 1.145 4.590 1.375 ;
        RECT  4.205 1.000 4.280 1.375 ;
        RECT  3.690 1.145 4.205 1.375 ;
        RECT  3.570 1.025 3.690 1.375 ;
        RECT  3.290 1.145 3.570 1.375 ;
        RECT  3.200 0.995 3.290 1.375 ;
        RECT  3.125 1.145 3.200 1.375 ;
        RECT  3.005 0.895 3.125 1.375 ;
        RECT  2.335 1.145 3.005 1.375 ;
        RECT  2.225 0.930 2.335 1.375 ;
        RECT  1.640 1.145 2.225 1.375 ;
        RECT  1.520 1.070 1.640 1.375 ;
        RECT  0.730 1.145 1.520 1.375 ;
        RECT  0.610 1.055 0.730 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.220 1.040 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.745 4.880 1.000 ;
        RECT  4.865 0.205 4.870 0.485 ;
        RECT  4.480 0.355 4.515 0.485 ;
        RECT  4.480 0.710 4.515 0.830 ;
        RECT  4.400 0.205 4.480 0.485 ;
        RECT  4.400 0.710 4.480 1.000 ;
        RECT  4.255 0.210 4.330 0.925 ;
        RECT  3.380 0.210 4.255 0.280 ;
        RECT  3.300 0.855 4.255 0.925 ;
        RECT  3.185 0.360 4.090 0.430 ;
        RECT  3.675 0.515 3.925 0.675 ;
        RECT  2.705 0.570 3.495 0.640 ;
        RECT  3.230 0.720 3.300 0.925 ;
        RECT  2.930 0.720 3.230 0.790 ;
        RECT  2.730 0.995 2.880 1.075 ;
        RECT  2.695 0.815 2.765 0.885 ;
        RECT  2.485 0.995 2.730 1.065 ;
        RECT  2.695 0.310 2.705 0.640 ;
        RECT  2.625 0.310 2.695 0.885 ;
        RECT  2.485 0.195 2.550 0.265 ;
        RECT  2.405 0.195 2.485 1.065 ;
        RECT  2.235 0.335 2.305 0.850 ;
        RECT  1.880 0.335 2.235 0.405 ;
        RECT  1.490 0.780 2.235 0.850 ;
        RECT  1.810 0.545 2.150 0.615 ;
        RECT  1.350 0.930 1.845 1.000 ;
        RECT  1.740 0.330 1.810 0.615 ;
        RECT  1.575 0.330 1.740 0.400 ;
        RECT  1.560 0.480 1.670 0.700 ;
        RECT  1.505 0.215 1.575 0.400 ;
        RECT  0.795 0.215 1.505 0.285 ;
        RECT  1.420 0.610 1.490 0.850 ;
        RECT  1.280 0.355 1.350 1.000 ;
        RECT  1.230 0.355 1.280 0.425 ;
        RECT  1.140 0.505 1.210 0.985 ;
        RECT  0.850 0.905 1.140 0.985 ;
        RECT  1.000 0.705 1.070 0.825 ;
        RECT  0.795 0.705 1.000 0.775 ;
        RECT  0.790 0.875 0.850 0.985 ;
        RECT  0.725 0.215 0.795 0.775 ;
        RECT  0.345 0.875 0.790 0.960 ;
        RECT  0.555 0.350 0.625 0.790 ;
        RECT  0.415 0.350 0.555 0.420 ;
        RECT  0.415 0.720 0.555 0.790 ;
        RECT  0.345 0.525 0.385 0.645 ;
        RECT  0.275 0.340 0.345 0.960 ;
        RECT  0.125 0.340 0.275 0.415 ;
        RECT  0.130 0.875 0.275 0.960 ;
        RECT  0.055 0.875 0.130 1.065 ;
        RECT  0.055 0.195 0.125 0.415 ;
        LAYER VIA1 ;
        RECT  3.740 0.525 3.810 0.595 ;
        RECT  1.580 0.525 1.650 0.595 ;
    END
END DFNCNQD4BWP40

MACRO DFNCSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFNCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.215 4.585 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.021400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.410 -0.115 4.620 0.115 ;
        RECT  4.275 -0.115 4.410 0.350 ;
        RECT  3.380 -0.115 4.275 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.400 ;
        RECT  0.730 -0.115 2.475 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.260 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.955 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.715 1.145 1.530 1.375 ;
        RECT  0.590 1.045 0.715 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.000 ;
        RECT  2.940 0.930 4.095 1.000 ;
        RECT  3.805 0.510 4.025 0.630 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.790 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.365 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.880 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.205 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  1.110 0.205 2.335 0.275 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.390 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.355 1.920 0.425 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.250 0.850 1.820 0.920 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.320 0.505 1.390 0.715 ;
        RECT  1.250 0.355 1.330 0.425 ;
        RECT  1.180 0.355 1.250 0.920 ;
        RECT  1.040 0.205 1.110 0.915 ;
        RECT  0.960 0.840 1.040 0.915 ;
        RECT  0.810 0.875 0.880 1.060 ;
        RECT  0.760 0.875 0.810 0.955 ;
        RECT  0.685 0.350 0.760 0.955 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.515 0.875 0.685 0.955 ;
        RECT  0.460 0.205 0.540 0.420 ;
        RECT  0.440 0.875 0.515 1.065 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.915 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.135 0.845 0.290 0.915 ;
        RECT  0.080 0.205 0.160 0.410 ;
        RECT  0.060 0.845 0.135 1.065 ;
    END
END DFNCSNQD0BWP40

MACRO DFNCSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFNCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.205 4.585 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.020800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.022400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.385 -0.115 4.620 0.115 ;
        RECT  4.295 -0.115 4.385 0.310 ;
        RECT  3.380 -0.115 4.295 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.400 ;
        RECT  0.730 -0.115 2.475 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.260 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.145 4.620 1.375 ;
        RECT  4.280 0.855 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.715 1.145 1.530 1.375 ;
        RECT  0.590 1.045 0.715 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.000 ;
        RECT  2.940 0.930 4.095 1.000 ;
        RECT  3.805 0.460 4.025 0.580 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.880 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.205 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  1.110 0.205 2.335 0.275 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.390 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.355 1.920 0.425 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.250 0.850 1.820 0.920 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.320 0.505 1.390 0.710 ;
        RECT  1.250 0.355 1.330 0.425 ;
        RECT  1.180 0.355 1.250 0.920 ;
        RECT  1.040 0.205 1.110 0.915 ;
        RECT  0.960 0.840 1.040 0.915 ;
        RECT  0.810 0.875 0.880 1.060 ;
        RECT  0.760 0.875 0.810 0.945 ;
        RECT  0.685 0.350 0.760 0.945 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.510 0.875 0.685 0.945 ;
        RECT  0.460 0.205 0.540 0.420 ;
        RECT  0.440 0.875 0.510 1.065 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.915 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.135 0.845 0.290 0.915 ;
        RECT  0.080 0.205 0.160 0.410 ;
        RECT  0.060 0.845 0.135 1.065 ;
    END
END DFNCSNQD1BWP40

MACRO DFNCSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFNCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.450 4.340 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.195 4.585 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.020800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.022400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.490 3.485 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 -0.115 4.900 0.115 ;
        RECT  4.760 -0.115 4.830 0.485 ;
        RECT  4.410 -0.115 4.760 0.115 ;
        RECT  4.275 -0.115 4.410 0.310 ;
        RECT  3.380 -0.115 4.275 0.115 ;
        RECT  3.245 -0.115 3.380 0.250 ;
        RECT  2.545 -0.115 3.245 0.115 ;
        RECT  2.475 -0.115 2.545 0.400 ;
        RECT  0.730 -0.115 2.475 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.260 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 1.145 4.900 1.375 ;
        RECT  4.760 0.690 4.830 1.375 ;
        RECT  4.400 1.145 4.760 1.375 ;
        RECT  4.280 0.955 4.400 1.375 ;
        RECT  3.995 1.145 4.280 1.375 ;
        RECT  3.865 1.095 3.995 1.375 ;
        RECT  3.390 1.145 3.865 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.715 1.145 1.530 1.375 ;
        RECT  0.590 1.045 0.715 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.095 0.285 4.165 1.000 ;
        RECT  2.940 0.930 4.095 1.000 ;
        RECT  3.805 0.460 4.025 0.580 ;
        RECT  3.480 0.195 3.995 0.265 ;
        RECT  3.730 0.335 3.805 0.860 ;
        RECT  3.695 0.335 3.730 0.445 ;
        RECT  3.470 0.790 3.730 0.860 ;
        RECT  3.625 0.520 3.650 0.700 ;
        RECT  3.555 0.340 3.625 0.700 ;
        RECT  3.050 0.340 3.555 0.410 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.980 0.195 3.050 0.410 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.705 0.195 2.980 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.880 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.205 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  1.110 0.205 2.335 0.275 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.390 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.355 1.920 0.425 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.250 0.850 1.820 0.920 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.320 0.505 1.390 0.710 ;
        RECT  1.250 0.355 1.325 0.425 ;
        RECT  1.180 0.355 1.250 0.920 ;
        RECT  1.040 0.205 1.110 0.915 ;
        RECT  0.960 0.840 1.040 0.915 ;
        RECT  0.810 0.875 0.880 1.060 ;
        RECT  0.760 0.875 0.810 0.945 ;
        RECT  0.685 0.350 0.760 0.945 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.600 0.825 0.685 0.945 ;
        RECT  0.515 0.875 0.600 0.955 ;
        RECT  0.460 0.205 0.540 0.420 ;
        RECT  0.440 0.875 0.515 1.065 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.915 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.135 0.845 0.290 0.915 ;
        RECT  0.080 0.205 0.160 0.410 ;
        RECT  0.060 0.845 0.135 1.065 ;
    END
END DFNCSNQD2BWP40

MACRO DFNCSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFNCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.450 4.890 0.765 ;
        RECT  4.785 0.525 4.795 0.635 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.425 0.195 5.520 0.485 ;
        RECT  5.425 0.710 5.520 0.995 ;
        RECT  5.355 0.355 5.425 0.485 ;
        RECT  5.355 0.710 5.425 0.830 ;
        RECT  5.145 0.355 5.355 0.830 ;
        RECT  5.120 0.355 5.145 0.485 ;
        RECT  5.120 0.710 5.145 0.830 ;
        RECT  5.045 0.215 5.120 0.485 ;
        RECT  5.045 0.710 5.120 0.995 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.020800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.960 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.210 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.044600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.335 0.355 3.465 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 -0.115 5.740 0.115 ;
        RECT  5.615 -0.115 5.685 0.440 ;
        RECT  5.310 -0.115 5.615 0.115 ;
        RECT  5.225 -0.115 5.310 0.265 ;
        RECT  4.940 -0.115 5.225 0.115 ;
        RECT  4.850 -0.115 4.940 0.310 ;
        RECT  4.190 -0.115 4.850 0.115 ;
        RECT  4.070 -0.115 4.190 0.140 ;
        RECT  3.390 -0.115 4.070 0.115 ;
        RECT  3.255 -0.115 3.390 0.130 ;
        RECT  2.545 -0.115 3.255 0.115 ;
        RECT  2.475 -0.115 2.545 0.400 ;
        RECT  0.730 -0.115 2.475 0.115 ;
        RECT  0.620 -0.115 0.730 0.270 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.260 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.145 5.740 1.375 ;
        RECT  5.615 0.680 5.685 1.375 ;
        RECT  5.330 1.145 5.615 1.375 ;
        RECT  5.210 0.910 5.330 1.375 ;
        RECT  4.930 1.145 5.210 1.375 ;
        RECT  4.855 0.860 4.930 1.375 ;
        RECT  4.020 1.145 4.855 1.375 ;
        RECT  3.900 1.070 4.020 1.375 ;
        RECT  3.390 1.145 3.900 1.375 ;
        RECT  3.270 1.070 3.390 1.375 ;
        RECT  1.690 1.145 3.270 1.375 ;
        RECT  1.530 1.130 1.690 1.375 ;
        RECT  0.715 1.145 1.530 1.375 ;
        RECT  0.590 1.045 0.715 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.005 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.195 5.520 0.485 ;
        RECT  5.425 0.710 5.520 0.995 ;
        RECT  5.045 0.215 5.075 0.485 ;
        RECT  5.045 0.710 5.075 0.995 ;
        RECT  4.645 0.210 4.715 1.000 ;
        RECT  4.065 0.930 4.645 1.000 ;
        RECT  4.535 0.620 4.575 0.740 ;
        RECT  4.465 0.210 4.535 0.860 ;
        RECT  3.785 0.210 4.465 0.280 ;
        RECT  4.350 0.790 4.465 0.860 ;
        RECT  3.865 0.350 4.370 0.420 ;
        RECT  3.985 0.605 4.065 1.000 ;
        RECT  2.940 0.930 3.985 1.000 ;
        RECT  3.715 0.210 3.785 0.860 ;
        RECT  3.710 0.335 3.715 0.860 ;
        RECT  3.695 0.335 3.710 0.445 ;
        RECT  3.225 0.790 3.710 0.860 ;
        RECT  3.605 0.580 3.640 0.700 ;
        RECT  3.535 0.200 3.605 0.700 ;
        RECT  3.000 0.200 3.535 0.270 ;
        RECT  3.155 0.445 3.225 0.860 ;
        RECT  3.010 0.535 3.085 0.785 ;
        RECT  2.900 0.535 3.010 0.605 ;
        RECT  2.955 0.195 3.000 0.270 ;
        RECT  2.705 0.195 2.955 0.265 ;
        RECT  2.865 0.825 2.940 1.000 ;
        RECT  2.705 0.685 2.930 0.755 ;
        RECT  2.785 0.355 2.900 0.605 ;
        RECT  2.475 0.825 2.865 0.900 ;
        RECT  2.620 0.970 2.775 1.060 ;
        RECT  2.635 0.195 2.705 0.755 ;
        RECT  0.880 0.990 2.620 1.060 ;
        RECT  2.405 0.825 2.475 0.915 ;
        RECT  2.405 0.485 2.415 0.625 ;
        RECT  2.335 0.205 2.405 0.625 ;
        RECT  2.045 0.840 2.405 0.915 ;
        RECT  1.110 0.205 2.335 0.275 ;
        RECT  2.205 0.355 2.265 0.575 ;
        RECT  2.185 0.355 2.205 0.760 ;
        RECT  2.115 0.505 2.185 0.760 ;
        RECT  1.390 0.505 2.115 0.575 ;
        RECT  1.975 0.645 2.045 0.915 ;
        RECT  1.670 0.645 1.975 0.715 ;
        RECT  1.425 0.355 1.920 0.425 ;
        RECT  1.820 0.800 1.895 0.920 ;
        RECT  1.250 0.850 1.820 0.920 ;
        RECT  1.575 0.645 1.670 0.770 ;
        RECT  1.320 0.505 1.390 0.710 ;
        RECT  1.250 0.355 1.330 0.425 ;
        RECT  1.180 0.355 1.250 0.920 ;
        RECT  1.040 0.205 1.110 0.915 ;
        RECT  0.960 0.840 1.040 0.915 ;
        RECT  0.810 0.875 0.880 1.060 ;
        RECT  0.760 0.875 0.810 0.945 ;
        RECT  0.685 0.350 0.760 0.945 ;
        RECT  0.540 0.350 0.685 0.420 ;
        RECT  0.515 0.865 0.685 0.945 ;
        RECT  0.460 0.205 0.540 0.420 ;
        RECT  0.440 0.865 0.515 1.065 ;
        RECT  0.360 0.520 0.410 0.640 ;
        RECT  0.290 0.340 0.360 0.915 ;
        RECT  0.160 0.340 0.290 0.410 ;
        RECT  0.135 0.845 0.290 0.915 ;
        RECT  0.080 0.205 0.160 0.410 ;
        RECT  0.060 0.845 0.135 1.065 ;
    END
END DFNCSNQD4BWP40

MACRO DFNQD0BWP40
    CLASS CORE ;
    FOREIGN DFNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.195 3.325 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.115 3.360 0.115 ;
        RECT  3.040 -0.115 3.110 0.295 ;
        RECT  2.740 -0.115 3.040 0.115 ;
        RECT  2.670 -0.115 2.740 0.325 ;
        RECT  1.935 -0.115 2.670 0.115 ;
        RECT  1.815 -0.115 1.935 0.125 ;
        RECT  1.275 -0.115 1.815 0.115 ;
        RECT  1.145 -0.115 1.275 0.125 ;
        RECT  0.370 -0.115 1.145 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 1.145 3.360 1.375 ;
        RECT  3.040 0.945 3.110 1.375 ;
        RECT  2.735 1.145 3.040 1.375 ;
        RECT  2.605 1.130 2.735 1.375 ;
        RECT  1.935 1.145 2.605 1.375 ;
        RECT  1.815 1.135 1.935 1.375 ;
        RECT  1.275 1.145 1.815 1.375 ;
        RECT  1.155 1.135 1.275 1.375 ;
        RECT  0.395 1.145 1.155 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.085 0.405 3.155 0.815 ;
        RECT  2.930 0.405 3.085 0.475 ;
        RECT  2.930 0.745 3.085 0.815 ;
        RECT  2.860 0.195 2.930 0.475 ;
        RECT  2.860 0.745 2.930 0.955 ;
        RECT  2.610 0.405 2.860 0.475 ;
        RECT  2.780 0.545 2.845 0.615 ;
        RECT  2.710 0.545 2.780 0.910 ;
        RECT  2.255 0.840 2.710 0.910 ;
        RECT  2.540 0.405 2.610 0.580 ;
        RECT  2.395 0.685 2.505 0.755 ;
        RECT  2.325 0.195 2.395 0.755 ;
        RECT  2.225 0.195 2.325 0.265 ;
        RECT  2.175 0.345 2.255 0.910 ;
        RECT  2.105 0.985 2.235 1.075 ;
        RECT  2.075 0.185 2.225 0.265 ;
        RECT  0.470 0.985 2.105 1.055 ;
        RECT  1.815 0.195 2.075 0.265 ;
        RECT  1.885 0.520 1.960 0.905 ;
        RECT  1.295 0.835 1.885 0.905 ;
        RECT  1.745 0.195 1.815 0.765 ;
        RECT  0.975 0.195 1.745 0.265 ;
        RECT  1.595 0.695 1.745 0.765 ;
        RECT  1.435 0.345 1.505 0.765 ;
        RECT  1.155 0.345 1.435 0.415 ;
        RECT  1.395 0.695 1.435 0.765 ;
        RECT  1.295 0.520 1.350 0.635 ;
        RECT  1.225 0.520 1.295 0.905 ;
        RECT  0.855 0.835 1.225 0.905 ;
        RECT  1.085 0.345 1.155 0.625 ;
        RECT  1.065 0.535 1.085 0.625 ;
        RECT  0.995 0.695 1.075 0.765 ;
        RECT  0.995 0.350 1.015 0.470 ;
        RECT  0.925 0.350 0.995 0.765 ;
        RECT  0.845 0.185 0.975 0.265 ;
        RECT  0.775 0.350 0.855 0.905 ;
        RECT  0.295 0.195 0.845 0.265 ;
        RECT  0.665 0.350 0.775 0.420 ;
        RECT  0.635 0.835 0.775 0.905 ;
        RECT  0.380 0.390 0.470 1.055 ;
        RECT  0.155 0.985 0.380 1.055 ;
        RECT  0.225 0.195 0.295 0.715 ;
        RECT  0.085 0.205 0.155 1.055 ;
        RECT  0.055 0.205 0.085 0.325 ;
        RECT  0.035 0.985 0.085 1.055 ;
    END
END DFNQD0BWP40

MACRO DFNQD1BWP40
    CLASS CORE ;
    FOREIGN DFNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.195 3.325 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.115 3.360 0.115 ;
        RECT  3.040 -0.115 3.110 0.325 ;
        RECT  2.740 -0.115 3.040 0.115 ;
        RECT  2.670 -0.115 2.740 0.325 ;
        RECT  1.935 -0.115 2.670 0.115 ;
        RECT  1.815 -0.115 1.935 0.125 ;
        RECT  1.275 -0.115 1.815 0.115 ;
        RECT  1.145 -0.115 1.275 0.125 ;
        RECT  0.370 -0.115 1.145 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 1.145 3.360 1.375 ;
        RECT  3.040 0.845 3.110 1.375 ;
        RECT  2.770 1.145 3.040 1.375 ;
        RECT  2.640 1.010 2.770 1.375 ;
        RECT  1.935 1.145 2.640 1.375 ;
        RECT  1.815 1.135 1.935 1.375 ;
        RECT  1.275 1.145 1.815 1.375 ;
        RECT  1.155 1.135 1.275 1.375 ;
        RECT  0.395 1.145 1.155 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.085 0.405 3.155 0.765 ;
        RECT  2.930 0.405 3.085 0.475 ;
        RECT  2.930 0.695 3.085 0.765 ;
        RECT  2.860 0.195 2.930 0.475 ;
        RECT  2.860 0.695 2.930 0.955 ;
        RECT  2.780 0.545 2.890 0.615 ;
        RECT  2.610 0.405 2.860 0.475 ;
        RECT  2.710 0.545 2.780 0.910 ;
        RECT  2.255 0.840 2.710 0.910 ;
        RECT  2.540 0.405 2.610 0.580 ;
        RECT  2.395 0.685 2.505 0.755 ;
        RECT  2.325 0.195 2.395 0.755 ;
        RECT  2.225 0.195 2.325 0.265 ;
        RECT  2.175 0.345 2.255 0.910 ;
        RECT  2.105 0.985 2.235 1.075 ;
        RECT  2.075 0.185 2.225 0.265 ;
        RECT  0.470 0.985 2.105 1.055 ;
        RECT  1.815 0.195 2.075 0.265 ;
        RECT  1.885 0.520 1.960 0.905 ;
        RECT  1.295 0.835 1.885 0.905 ;
        RECT  1.745 0.195 1.815 0.765 ;
        RECT  0.975 0.195 1.745 0.265 ;
        RECT  1.600 0.695 1.745 0.765 ;
        RECT  1.435 0.345 1.505 0.765 ;
        RECT  1.155 0.345 1.435 0.415 ;
        RECT  1.395 0.695 1.435 0.765 ;
        RECT  1.295 0.520 1.350 0.635 ;
        RECT  1.225 0.520 1.295 0.905 ;
        RECT  0.855 0.835 1.225 0.905 ;
        RECT  1.085 0.345 1.155 0.625 ;
        RECT  1.065 0.535 1.085 0.625 ;
        RECT  0.995 0.695 1.075 0.765 ;
        RECT  0.995 0.350 1.015 0.470 ;
        RECT  0.925 0.350 0.995 0.765 ;
        RECT  0.845 0.185 0.975 0.265 ;
        RECT  0.775 0.350 0.855 0.905 ;
        RECT  0.305 0.195 0.845 0.265 ;
        RECT  0.665 0.350 0.775 0.420 ;
        RECT  0.635 0.835 0.775 0.905 ;
        RECT  0.380 0.390 0.470 1.055 ;
        RECT  0.160 0.985 0.380 1.055 ;
        RECT  0.235 0.195 0.305 0.715 ;
        RECT  0.090 0.205 0.160 1.055 ;
        RECT  0.055 0.205 0.090 0.325 ;
        RECT  0.035 0.985 0.090 1.055 ;
    END
END DFNQD1BWP40

MACRO DFNQD2BWP40
    CLASS CORE ;
    FOREIGN DFNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.195 3.340 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 -0.115 3.640 0.115 ;
        RECT  3.515 -0.115 3.585 0.430 ;
        RECT  3.110 -0.115 3.515 0.115 ;
        RECT  3.040 -0.115 3.110 0.315 ;
        RECT  2.740 -0.115 3.040 0.115 ;
        RECT  2.670 -0.115 2.740 0.315 ;
        RECT  1.935 -0.115 2.670 0.115 ;
        RECT  1.815 -0.115 1.935 0.125 ;
        RECT  1.275 -0.115 1.815 0.115 ;
        RECT  1.145 -0.115 1.275 0.125 ;
        RECT  0.370 -0.115 1.145 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 1.145 3.640 1.375 ;
        RECT  3.515 0.700 3.585 1.375 ;
        RECT  3.110 1.145 3.515 1.375 ;
        RECT  3.040 0.845 3.110 1.375 ;
        RECT  2.765 1.145 3.040 1.375 ;
        RECT  2.645 1.030 2.765 1.375 ;
        RECT  1.935 1.145 2.645 1.375 ;
        RECT  1.815 1.135 1.935 1.375 ;
        RECT  1.275 1.145 1.815 1.375 ;
        RECT  1.155 1.135 1.275 1.375 ;
        RECT  0.395 1.145 1.155 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.095 0.395 3.165 0.765 ;
        RECT  2.930 0.395 3.095 0.465 ;
        RECT  2.930 0.695 3.095 0.765 ;
        RECT  2.860 0.195 2.930 0.465 ;
        RECT  2.860 0.695 2.930 0.955 ;
        RECT  2.780 0.545 2.885 0.615 ;
        RECT  2.610 0.395 2.860 0.465 ;
        RECT  2.710 0.545 2.780 0.910 ;
        RECT  2.255 0.840 2.710 0.910 ;
        RECT  2.540 0.395 2.610 0.580 ;
        RECT  2.395 0.685 2.505 0.755 ;
        RECT  2.325 0.195 2.395 0.755 ;
        RECT  2.225 0.195 2.325 0.265 ;
        RECT  2.175 0.345 2.255 0.910 ;
        RECT  2.105 0.985 2.235 1.075 ;
        RECT  2.075 0.185 2.225 0.265 ;
        RECT  0.470 0.985 2.105 1.055 ;
        RECT  1.815 0.195 2.075 0.265 ;
        RECT  1.885 0.520 1.960 0.905 ;
        RECT  1.295 0.835 1.885 0.905 ;
        RECT  1.745 0.195 1.815 0.765 ;
        RECT  0.975 0.195 1.745 0.265 ;
        RECT  1.600 0.695 1.745 0.765 ;
        RECT  1.435 0.345 1.505 0.765 ;
        RECT  1.155 0.345 1.435 0.415 ;
        RECT  1.395 0.695 1.435 0.765 ;
        RECT  1.295 0.520 1.350 0.635 ;
        RECT  1.225 0.520 1.295 0.905 ;
        RECT  0.855 0.835 1.225 0.905 ;
        RECT  1.085 0.345 1.155 0.625 ;
        RECT  1.065 0.535 1.085 0.625 ;
        RECT  0.995 0.695 1.075 0.765 ;
        RECT  0.995 0.350 1.015 0.470 ;
        RECT  0.925 0.350 0.995 0.765 ;
        RECT  0.845 0.185 0.975 0.265 ;
        RECT  0.775 0.350 0.855 0.905 ;
        RECT  0.305 0.195 0.845 0.265 ;
        RECT  0.665 0.350 0.775 0.420 ;
        RECT  0.635 0.835 0.775 0.905 ;
        RECT  0.380 0.390 0.470 1.055 ;
        RECT  0.160 0.985 0.380 1.055 ;
        RECT  0.235 0.195 0.305 0.715 ;
        RECT  0.090 0.205 0.160 1.055 ;
        RECT  0.055 0.205 0.090 0.325 ;
        RECT  0.035 0.985 0.090 1.055 ;
    END
END DFNQD2BWP40

MACRO DFNQD4BWP40
    CLASS CORE ;
    FOREIGN DFNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.885 0.195 3.980 0.475 ;
        RECT  3.885 0.665 3.980 1.065 ;
        RECT  3.815 0.355 3.885 0.475 ;
        RECT  3.815 0.665 3.885 0.785 ;
        RECT  3.605 0.355 3.815 0.785 ;
        RECT  3.575 0.355 3.605 0.480 ;
        RECT  3.575 0.665 3.605 0.785 ;
        RECT  3.505 0.215 3.575 0.480 ;
        RECT  3.505 0.665 3.575 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.675 0.625 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.075 -0.115 4.150 0.420 ;
        RECT  3.770 -0.115 4.075 0.115 ;
        RECT  3.690 -0.115 3.770 0.275 ;
        RECT  3.380 -0.115 3.690 0.115 ;
        RECT  3.310 -0.115 3.380 0.325 ;
        RECT  3.175 -0.115 3.310 0.115 ;
        RECT  3.105 -0.115 3.175 0.320 ;
        RECT  2.730 -0.115 3.105 0.115 ;
        RECT  2.660 -0.115 2.730 0.325 ;
        RECT  1.935 -0.115 2.660 0.115 ;
        RECT  1.815 -0.115 1.935 0.125 ;
        RECT  1.275 -0.115 1.815 0.115 ;
        RECT  1.145 -0.115 1.275 0.125 ;
        RECT  0.370 -0.115 1.145 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.075 0.685 4.150 1.375 ;
        RECT  3.785 1.145 4.075 1.375 ;
        RECT  3.675 0.905 3.785 1.375 ;
        RECT  3.380 1.145 3.675 1.375 ;
        RECT  3.310 0.845 3.380 1.375 ;
        RECT  3.175 1.145 3.310 1.375 ;
        RECT  3.105 0.845 3.175 1.375 ;
        RECT  2.735 1.145 3.105 1.375 ;
        RECT  2.605 1.130 2.735 1.375 ;
        RECT  1.910 1.145 2.605 1.375 ;
        RECT  1.790 1.045 1.910 1.375 ;
        RECT  1.275 1.145 1.790 1.375 ;
        RECT  1.155 1.135 1.275 1.375 ;
        RECT  0.395 1.145 1.155 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.195 3.980 0.475 ;
        RECT  3.885 0.665 3.980 1.065 ;
        RECT  3.505 0.215 3.535 0.480 ;
        RECT  3.505 0.665 3.535 1.065 ;
        RECT  3.335 0.405 3.405 0.765 ;
        RECT  2.920 0.405 3.335 0.475 ;
        RECT  2.920 0.695 3.335 0.765 ;
        RECT  2.770 0.545 2.970 0.615 ;
        RECT  2.850 0.195 2.920 0.475 ;
        RECT  2.850 0.695 2.920 1.030 ;
        RECT  2.610 0.405 2.850 0.475 ;
        RECT  2.700 0.545 2.770 0.910 ;
        RECT  2.255 0.840 2.700 0.910 ;
        RECT  2.540 0.405 2.610 0.580 ;
        RECT  2.395 0.690 2.505 0.760 ;
        RECT  2.325 0.195 2.395 0.760 ;
        RECT  2.225 0.195 2.325 0.265 ;
        RECT  2.175 0.345 2.255 0.910 ;
        RECT  2.075 0.185 2.225 0.265 ;
        RECT  1.825 0.195 2.075 0.265 ;
        RECT  1.895 0.505 1.970 0.905 ;
        RECT  1.295 0.835 1.895 0.905 ;
        RECT  1.755 0.195 1.825 0.765 ;
        RECT  0.975 0.195 1.755 0.265 ;
        RECT  1.580 0.695 1.755 0.765 ;
        RECT  1.510 0.985 1.630 1.075 ;
        RECT  0.470 0.985 1.510 1.055 ;
        RECT  1.425 0.345 1.500 0.765 ;
        RECT  1.155 0.345 1.425 0.415 ;
        RECT  1.390 0.695 1.425 0.765 ;
        RECT  1.295 0.520 1.350 0.635 ;
        RECT  1.225 0.520 1.295 0.905 ;
        RECT  0.855 0.835 1.225 0.905 ;
        RECT  1.085 0.345 1.155 0.625 ;
        RECT  1.065 0.535 1.085 0.625 ;
        RECT  0.995 0.695 1.075 0.765 ;
        RECT  0.995 0.350 1.015 0.470 ;
        RECT  0.925 0.350 0.995 0.765 ;
        RECT  0.845 0.185 0.975 0.265 ;
        RECT  0.775 0.350 0.855 0.905 ;
        RECT  0.310 0.195 0.845 0.265 ;
        RECT  0.665 0.350 0.775 0.420 ;
        RECT  0.635 0.835 0.775 0.905 ;
        RECT  0.380 0.390 0.470 1.055 ;
        RECT  0.160 0.985 0.380 1.055 ;
        RECT  0.240 0.195 0.310 0.705 ;
        RECT  0.090 0.205 0.160 1.055 ;
        RECT  0.055 0.205 0.090 0.325 ;
        RECT  0.035 0.985 0.090 1.055 ;
    END
END DFNQD4BWP40

MACRO DFNSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFNSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.685 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.075 ;
        RECT  4.075 0.185 4.095 0.310 ;
        RECT  4.075 0.950 4.095 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.705 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.790 0.670 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.935 -0.115 4.200 0.115 ;
        RECT  3.865 -0.115 3.935 0.290 ;
        RECT  2.965 -0.115 3.865 0.115 ;
        RECT  2.890 -0.115 2.965 0.240 ;
        RECT  2.310 -0.115 2.890 0.115 ;
        RECT  2.195 -0.115 2.310 0.215 ;
        RECT  1.285 -0.115 2.195 0.115 ;
        RECT  1.155 -0.115 1.285 0.125 ;
        RECT  0.370 -0.115 1.155 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.145 4.200 1.375 ;
        RECT  3.860 1.045 3.980 1.375 ;
        RECT  3.085 1.145 3.860 1.375 ;
        RECT  2.965 1.015 3.085 1.375 ;
        RECT  2.255 1.145 2.965 1.375 ;
        RECT  2.135 1.140 2.255 1.375 ;
        RECT  1.755 1.145 2.135 1.375 ;
        RECT  1.625 1.140 1.755 1.375 ;
        RECT  1.285 1.145 1.625 1.375 ;
        RECT  1.165 1.135 1.285 1.375 ;
        RECT  0.375 1.145 1.165 1.375 ;
        RECT  0.295 1.015 0.375 1.375 ;
        RECT  0.000 1.145 0.295 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.930 0.520 4.005 0.975 ;
        RECT  3.455 0.905 3.930 0.975 ;
        RECT  3.595 0.750 3.770 0.825 ;
        RECT  3.595 0.195 3.755 0.275 ;
        RECT  3.525 0.195 3.595 0.825 ;
        RECT  3.105 0.195 3.525 0.275 ;
        RECT  3.385 0.355 3.455 0.975 ;
        RECT  3.255 0.355 3.385 0.425 ;
        RECT  3.215 0.620 3.315 0.740 ;
        RECT  3.180 0.355 3.255 0.540 ;
        RECT  3.145 0.620 3.215 0.935 ;
        RECT  2.935 0.470 3.180 0.540 ;
        RECT  2.610 0.865 3.145 0.935 ;
        RECT  3.035 0.195 3.105 0.390 ;
        RECT  2.750 0.320 3.035 0.390 ;
        RECT  2.865 0.470 2.935 0.645 ;
        RECT  2.750 0.710 2.825 0.785 ;
        RECT  2.680 0.195 2.750 0.785 ;
        RECT  2.460 0.195 2.680 0.265 ;
        RECT  2.535 0.345 2.610 0.935 ;
        RECT  2.385 1.005 2.550 1.075 ;
        RECT  2.390 0.195 2.460 0.365 ;
        RECT  2.125 0.295 2.390 0.365 ;
        RECT  2.315 0.990 2.385 1.075 ;
        RECT  0.555 0.990 2.315 1.060 ;
        RECT  2.220 0.490 2.290 0.920 ;
        RECT  1.305 0.850 2.220 0.920 ;
        RECT  2.055 0.195 2.125 0.365 ;
        RECT  0.985 0.195 2.055 0.265 ;
        RECT  1.900 0.350 1.970 0.775 ;
        RECT  1.890 0.520 1.900 0.775 ;
        RECT  1.835 0.520 1.890 0.640 ;
        RECT  1.495 0.345 1.745 0.415 ;
        RECT  1.425 0.345 1.495 0.780 ;
        RECT  1.165 0.345 1.425 0.415 ;
        RECT  1.305 0.520 1.355 0.640 ;
        RECT  1.235 0.520 1.305 0.920 ;
        RECT  0.865 0.850 1.235 0.920 ;
        RECT  1.095 0.345 1.165 0.625 ;
        RECT  1.075 0.535 1.095 0.625 ;
        RECT  1.005 0.695 1.085 0.765 ;
        RECT  1.005 0.350 1.025 0.470 ;
        RECT  0.935 0.350 1.005 0.765 ;
        RECT  0.855 0.185 0.985 0.265 ;
        RECT  0.785 0.350 0.865 0.920 ;
        RECT  0.290 0.195 0.855 0.265 ;
        RECT  0.675 0.350 0.785 0.420 ;
        RECT  0.655 0.850 0.785 0.920 ;
        RECT  0.465 0.855 0.555 1.060 ;
        RECT  0.375 0.390 0.465 0.925 ;
        RECT  0.155 0.855 0.375 0.925 ;
        RECT  0.220 0.195 0.290 0.705 ;
        RECT  0.150 0.855 0.155 1.045 ;
        RECT  0.080 0.205 0.150 1.045 ;
        RECT  0.055 0.205 0.080 0.325 ;
    END
END DFNSNQD0BWP40

MACRO DFNSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFNSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.685 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.185 4.165 1.075 ;
        RECT  4.075 0.185 4.095 0.465 ;
        RECT  4.075 0.685 4.095 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.705 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.790 0.670 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.935 -0.115 4.200 0.115 ;
        RECT  3.865 -0.115 3.935 0.420 ;
        RECT  2.965 -0.115 3.865 0.115 ;
        RECT  2.890 -0.115 2.965 0.240 ;
        RECT  2.310 -0.115 2.890 0.115 ;
        RECT  2.195 -0.115 2.310 0.215 ;
        RECT  1.285 -0.115 2.195 0.115 ;
        RECT  1.155 -0.115 1.285 0.125 ;
        RECT  0.370 -0.115 1.155 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.145 4.200 1.375 ;
        RECT  3.860 1.045 3.980 1.375 ;
        RECT  3.085 1.145 3.860 1.375 ;
        RECT  2.965 1.015 3.085 1.375 ;
        RECT  2.255 1.145 2.965 1.375 ;
        RECT  2.135 1.140 2.255 1.375 ;
        RECT  1.755 1.145 2.135 1.375 ;
        RECT  1.625 1.140 1.755 1.375 ;
        RECT  1.285 1.145 1.625 1.375 ;
        RECT  1.165 1.135 1.285 1.375 ;
        RECT  0.375 1.145 1.165 1.375 ;
        RECT  0.300 1.015 0.375 1.375 ;
        RECT  0.000 1.145 0.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.930 0.520 4.005 0.975 ;
        RECT  3.455 0.905 3.930 0.975 ;
        RECT  3.595 0.750 3.770 0.825 ;
        RECT  3.595 0.195 3.755 0.275 ;
        RECT  3.525 0.195 3.595 0.825 ;
        RECT  3.105 0.195 3.525 0.275 ;
        RECT  3.385 0.355 3.455 0.975 ;
        RECT  3.255 0.355 3.385 0.425 ;
        RECT  3.215 0.620 3.315 0.740 ;
        RECT  3.180 0.355 3.255 0.540 ;
        RECT  3.145 0.620 3.215 0.935 ;
        RECT  2.935 0.470 3.180 0.540 ;
        RECT  2.610 0.865 3.145 0.935 ;
        RECT  3.035 0.195 3.105 0.390 ;
        RECT  2.750 0.320 3.035 0.390 ;
        RECT  2.865 0.470 2.935 0.645 ;
        RECT  2.750 0.710 2.825 0.785 ;
        RECT  2.680 0.195 2.750 0.785 ;
        RECT  2.460 0.195 2.680 0.265 ;
        RECT  2.535 0.345 2.610 0.935 ;
        RECT  2.385 1.005 2.550 1.075 ;
        RECT  2.390 0.195 2.460 0.365 ;
        RECT  2.125 0.295 2.390 0.365 ;
        RECT  2.315 0.990 2.385 1.075 ;
        RECT  0.555 0.990 2.315 1.060 ;
        RECT  2.220 0.490 2.290 0.920 ;
        RECT  1.305 0.850 2.220 0.920 ;
        RECT  2.055 0.195 2.125 0.365 ;
        RECT  0.985 0.195 2.055 0.265 ;
        RECT  1.900 0.350 1.970 0.775 ;
        RECT  1.890 0.520 1.900 0.775 ;
        RECT  1.835 0.520 1.890 0.640 ;
        RECT  1.495 0.345 1.745 0.415 ;
        RECT  1.425 0.345 1.495 0.780 ;
        RECT  1.165 0.345 1.425 0.415 ;
        RECT  1.305 0.520 1.355 0.640 ;
        RECT  1.235 0.520 1.305 0.920 ;
        RECT  0.865 0.850 1.235 0.920 ;
        RECT  1.095 0.345 1.165 0.625 ;
        RECT  1.075 0.535 1.095 0.625 ;
        RECT  1.005 0.695 1.085 0.765 ;
        RECT  1.005 0.350 1.025 0.470 ;
        RECT  0.935 0.350 1.005 0.765 ;
        RECT  0.855 0.185 0.985 0.265 ;
        RECT  0.785 0.350 0.865 0.920 ;
        RECT  0.290 0.195 0.855 0.265 ;
        RECT  0.675 0.350 0.785 0.420 ;
        RECT  0.655 0.850 0.785 0.920 ;
        RECT  0.465 0.865 0.555 1.060 ;
        RECT  0.375 0.390 0.465 0.935 ;
        RECT  0.150 0.865 0.375 0.935 ;
        RECT  0.220 0.195 0.290 0.705 ;
        RECT  0.080 0.205 0.150 0.935 ;
        RECT  0.055 0.205 0.080 0.325 ;
    END
END DFNSNQD1BWP40

MACRO DFNSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFNSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.685 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.124000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.370 4.165 0.880 ;
        RECT  4.020 0.195 4.095 0.445 ;
        RECT  4.020 0.805 4.095 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.705 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.355 3.790 0.670 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.115 4.340 0.115 ;
        RECT  4.215 -0.115 4.285 0.255 ;
        RECT  3.900 -0.115 4.215 0.115 ;
        RECT  3.830 -0.115 3.900 0.265 ;
        RECT  2.965 -0.115 3.830 0.115 ;
        RECT  2.890 -0.115 2.965 0.240 ;
        RECT  2.310 -0.115 2.890 0.115 ;
        RECT  2.195 -0.115 2.310 0.215 ;
        RECT  1.285 -0.115 2.195 0.115 ;
        RECT  1.155 -0.115 1.285 0.125 ;
        RECT  0.370 -0.115 1.155 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 1.145 4.340 1.375 ;
        RECT  4.215 0.950 4.285 1.375 ;
        RECT  3.925 1.145 4.215 1.375 ;
        RECT  3.805 1.045 3.925 1.375 ;
        RECT  3.085 1.145 3.805 1.375 ;
        RECT  2.965 1.015 3.085 1.375 ;
        RECT  2.255 1.145 2.965 1.375 ;
        RECT  2.135 1.140 2.255 1.375 ;
        RECT  1.755 1.145 2.135 1.375 ;
        RECT  1.625 1.140 1.755 1.375 ;
        RECT  1.285 1.145 1.625 1.375 ;
        RECT  1.165 1.135 1.285 1.375 ;
        RECT  0.375 1.145 1.165 1.375 ;
        RECT  0.300 1.015 0.375 1.375 ;
        RECT  0.000 1.145 0.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.950 0.525 4.025 0.635 ;
        RECT  3.875 0.525 3.950 0.975 ;
        RECT  3.455 0.905 3.875 0.975 ;
        RECT  3.595 0.195 3.755 0.275 ;
        RECT  3.595 0.750 3.710 0.825 ;
        RECT  3.525 0.195 3.595 0.825 ;
        RECT  3.105 0.195 3.525 0.275 ;
        RECT  3.385 0.355 3.455 0.975 ;
        RECT  3.255 0.355 3.385 0.425 ;
        RECT  3.215 0.620 3.315 0.740 ;
        RECT  3.180 0.355 3.255 0.540 ;
        RECT  3.145 0.620 3.215 0.935 ;
        RECT  2.935 0.470 3.180 0.540 ;
        RECT  2.610 0.865 3.145 0.935 ;
        RECT  3.035 0.195 3.105 0.390 ;
        RECT  2.750 0.320 3.035 0.390 ;
        RECT  2.865 0.470 2.935 0.645 ;
        RECT  2.750 0.710 2.825 0.785 ;
        RECT  2.680 0.195 2.750 0.785 ;
        RECT  2.460 0.195 2.680 0.265 ;
        RECT  2.535 0.345 2.610 0.935 ;
        RECT  2.385 1.005 2.550 1.075 ;
        RECT  2.390 0.195 2.460 0.365 ;
        RECT  2.125 0.295 2.390 0.365 ;
        RECT  2.315 0.990 2.385 1.075 ;
        RECT  0.555 0.990 2.315 1.060 ;
        RECT  2.220 0.490 2.290 0.920 ;
        RECT  1.305 0.850 2.220 0.920 ;
        RECT  2.055 0.195 2.125 0.365 ;
        RECT  0.985 0.195 2.055 0.265 ;
        RECT  1.900 0.350 1.970 0.775 ;
        RECT  1.890 0.520 1.900 0.775 ;
        RECT  1.835 0.520 1.890 0.640 ;
        RECT  1.495 0.345 1.745 0.415 ;
        RECT  1.425 0.345 1.495 0.780 ;
        RECT  1.165 0.345 1.425 0.415 ;
        RECT  1.305 0.520 1.355 0.640 ;
        RECT  1.235 0.520 1.305 0.920 ;
        RECT  0.865 0.850 1.235 0.920 ;
        RECT  1.095 0.345 1.165 0.625 ;
        RECT  1.075 0.535 1.095 0.625 ;
        RECT  1.005 0.695 1.085 0.765 ;
        RECT  1.005 0.350 1.025 0.470 ;
        RECT  0.935 0.350 1.005 0.765 ;
        RECT  0.855 0.185 0.985 0.265 ;
        RECT  0.785 0.350 0.865 0.920 ;
        RECT  0.290 0.195 0.855 0.265 ;
        RECT  0.675 0.350 0.785 0.420 ;
        RECT  0.655 0.850 0.785 0.920 ;
        RECT  0.465 0.865 0.555 1.060 ;
        RECT  0.375 0.390 0.465 0.935 ;
        RECT  0.150 0.865 0.375 0.935 ;
        RECT  0.220 0.195 0.290 0.705 ;
        RECT  0.080 0.205 0.150 0.935 ;
        RECT  0.055 0.205 0.080 0.325 ;
    END
END DFNSNQD2BWP40

MACRO DFNSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFNSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.685 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.185 4.820 0.460 ;
        RECT  4.725 0.785 4.810 1.075 ;
        RECT  4.655 0.330 4.725 0.460 ;
        RECT  4.655 0.785 4.725 0.905 ;
        RECT  4.445 0.330 4.655 0.905 ;
        RECT  4.435 0.330 4.445 0.460 ;
        RECT  4.435 0.785 4.445 0.905 ;
        RECT  4.345 0.185 4.435 0.460 ;
        RECT  4.345 0.785 4.435 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.705 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.355 4.115 0.670 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.985 0.410 ;
        RECT  4.605 -0.115 4.915 0.115 ;
        RECT  4.535 -0.115 4.605 0.255 ;
        RECT  4.225 -0.115 4.535 0.115 ;
        RECT  4.155 -0.115 4.225 0.265 ;
        RECT  3.490 -0.115 4.155 0.115 ;
        RECT  3.370 -0.115 3.490 0.130 ;
        RECT  2.970 -0.115 3.370 0.115 ;
        RECT  2.895 -0.115 2.970 0.240 ;
        RECT  2.310 -0.115 2.895 0.115 ;
        RECT  2.195 -0.115 2.310 0.215 ;
        RECT  1.285 -0.115 2.195 0.115 ;
        RECT  1.155 -0.115 1.285 0.125 ;
        RECT  0.370 -0.115 1.155 0.115 ;
        RECT  0.250 -0.115 0.370 0.125 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 1.145 5.040 1.375 ;
        RECT  4.915 0.725 4.985 1.375 ;
        RECT  4.605 1.145 4.915 1.375 ;
        RECT  4.535 0.995 4.605 1.375 ;
        RECT  4.250 1.145 4.535 1.375 ;
        RECT  4.130 1.045 4.250 1.375 ;
        RECT  3.880 1.145 4.130 1.375 ;
        RECT  3.760 1.045 3.880 1.375 ;
        RECT  3.085 1.145 3.760 1.375 ;
        RECT  2.965 1.015 3.085 1.375 ;
        RECT  2.215 1.145 2.965 1.375 ;
        RECT  2.095 1.140 2.215 1.375 ;
        RECT  1.755 1.145 2.095 1.375 ;
        RECT  1.625 1.140 1.755 1.375 ;
        RECT  1.285 1.145 1.625 1.375 ;
        RECT  1.165 1.135 1.285 1.375 ;
        RECT  0.375 1.145 1.165 1.375 ;
        RECT  0.300 1.015 0.375 1.375 ;
        RECT  0.000 1.145 0.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.185 4.820 0.460 ;
        RECT  4.725 0.785 4.810 1.075 ;
        RECT  4.345 0.185 4.375 0.460 ;
        RECT  4.345 0.785 4.375 1.075 ;
        RECT  4.275 0.545 4.375 0.615 ;
        RECT  4.200 0.545 4.275 0.965 ;
        RECT  3.700 0.895 4.200 0.965 ;
        RECT  3.870 0.200 4.080 0.275 ;
        RECT  3.870 0.750 4.055 0.825 ;
        RECT  3.800 0.200 3.870 0.825 ;
        RECT  3.110 0.200 3.800 0.280 ;
        RECT  3.630 0.380 3.700 0.965 ;
        RECT  3.250 0.380 3.630 0.450 ;
        RECT  3.370 0.820 3.630 0.895 ;
        RECT  3.230 0.610 3.490 0.680 ;
        RECT  3.180 0.380 3.250 0.540 ;
        RECT  3.160 0.610 3.230 0.935 ;
        RECT  2.935 0.470 3.180 0.540 ;
        RECT  2.610 0.865 3.160 0.935 ;
        RECT  3.040 0.200 3.110 0.390 ;
        RECT  2.750 0.320 3.040 0.390 ;
        RECT  2.865 0.470 2.935 0.645 ;
        RECT  2.750 0.710 2.825 0.785 ;
        RECT  2.680 0.195 2.750 0.785 ;
        RECT  2.460 0.195 2.680 0.265 ;
        RECT  2.535 0.345 2.610 0.935 ;
        RECT  2.385 1.005 2.550 1.075 ;
        RECT  2.390 0.195 2.460 0.365 ;
        RECT  2.125 0.295 2.390 0.365 ;
        RECT  2.315 0.990 2.385 1.075 ;
        RECT  0.555 0.990 2.315 1.060 ;
        RECT  2.220 0.490 2.290 0.920 ;
        RECT  1.305 0.850 2.220 0.920 ;
        RECT  2.055 0.195 2.125 0.365 ;
        RECT  0.985 0.195 2.055 0.265 ;
        RECT  1.900 0.350 1.970 0.775 ;
        RECT  1.890 0.520 1.900 0.775 ;
        RECT  1.835 0.520 1.890 0.640 ;
        RECT  1.495 0.345 1.745 0.415 ;
        RECT  1.425 0.345 1.495 0.780 ;
        RECT  1.165 0.345 1.425 0.415 ;
        RECT  1.305 0.520 1.355 0.640 ;
        RECT  1.235 0.520 1.305 0.920 ;
        RECT  0.865 0.850 1.235 0.920 ;
        RECT  1.095 0.345 1.165 0.625 ;
        RECT  1.075 0.535 1.095 0.625 ;
        RECT  1.005 0.695 1.085 0.765 ;
        RECT  1.005 0.350 1.025 0.470 ;
        RECT  0.935 0.350 1.005 0.765 ;
        RECT  0.855 0.185 0.985 0.265 ;
        RECT  0.785 0.350 0.865 0.920 ;
        RECT  0.290 0.195 0.855 0.265 ;
        RECT  0.675 0.350 0.785 0.420 ;
        RECT  0.655 0.850 0.785 0.920 ;
        RECT  0.465 0.865 0.555 1.060 ;
        RECT  0.375 0.390 0.465 0.935 ;
        RECT  0.150 0.865 0.375 0.935 ;
        RECT  0.220 0.195 0.290 0.705 ;
        RECT  0.080 0.205 0.150 0.935 ;
        RECT  0.055 0.205 0.080 0.325 ;
    END
END DFNSNQD4BWP40

MACRO DFQD0BWP40
    CLASS CORE ;
    FOREIGN DFQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.195 3.185 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.970 0.315 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.735 -0.115 2.530 0.115 ;
        RECT  1.615 -0.115 1.735 0.125 ;
        RECT  1.155 -0.115 1.615 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.145 3.220 1.375 ;
        RECT  2.900 0.940 2.970 1.375 ;
        RECT  2.595 1.145 2.900 1.375 ;
        RECT  2.465 1.135 2.595 1.375 ;
        RECT  1.795 1.145 2.465 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.395 3.015 0.765 ;
        RECT  2.790 0.395 2.945 0.465 ;
        RECT  2.790 0.695 2.945 0.765 ;
        RECT  2.720 0.220 2.790 0.465 ;
        RECT  2.720 0.695 2.790 1.050 ;
        RECT  2.640 0.545 2.735 0.615 ;
        RECT  2.470 0.395 2.720 0.465 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.395 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  2.000 0.195 2.230 0.265 ;
        RECT  2.080 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.930 0.195 2.000 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  1.550 0.195 1.930 0.265 ;
        RECT  1.460 0.820 1.930 0.890 ;
        RECT  1.765 0.345 1.835 0.615 ;
        RECT  1.275 0.545 1.765 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.480 0.195 1.550 0.450 ;
        RECT  0.925 0.195 1.480 0.265 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.765 0.385 1.835 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.885 0.455 ;
    END
END DFQD0BWP40

MACRO DFQD1BWP40
    CLASS CORE ;
    FOREIGN DFQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.195 3.185 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.970 0.315 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.785 -0.115 2.530 0.115 ;
        RECT  1.665 -0.115 1.785 0.125 ;
        RECT  1.155 -0.115 1.665 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.145 3.220 1.375 ;
        RECT  2.900 0.845 2.970 1.375 ;
        RECT  2.630 1.145 2.900 1.375 ;
        RECT  2.500 1.025 2.630 1.375 ;
        RECT  1.795 1.145 2.500 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.395 3.015 0.765 ;
        RECT  2.790 0.395 2.945 0.465 ;
        RECT  2.790 0.695 2.945 0.765 ;
        RECT  2.720 0.195 2.790 0.465 ;
        RECT  2.720 0.695 2.790 1.050 ;
        RECT  2.640 0.545 2.735 0.615 ;
        RECT  2.470 0.395 2.720 0.465 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.395 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  1.995 0.195 2.230 0.265 ;
        RECT  2.075 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.925 0.195 1.995 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  0.925 0.195 1.925 0.265 ;
        RECT  1.460 0.820 1.925 0.890 ;
        RECT  1.595 0.545 1.835 0.615 ;
        RECT  1.525 0.345 1.595 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.275 0.545 1.525 0.615 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.525 0.385 1.595 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.645 0.455 ;
    END
END DFQD1BWP40

MACRO DFQD2BWP40
    CLASS CORE ;
    FOREIGN DFQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.100 0.195 3.205 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.430 -0.115 3.500 0.115 ;
        RECT  3.355 -0.115 3.430 0.460 ;
        RECT  2.970 -0.115 3.355 0.115 ;
        RECT  2.900 -0.115 2.970 0.315 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.785 -0.115 2.530 0.115 ;
        RECT  1.665 -0.115 1.785 0.125 ;
        RECT  1.155 -0.115 1.665 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.425 1.145 3.500 1.375 ;
        RECT  3.355 0.705 3.425 1.375 ;
        RECT  2.970 1.145 3.355 1.375 ;
        RECT  2.900 0.845 2.970 1.375 ;
        RECT  2.630 1.145 2.900 1.375 ;
        RECT  2.505 1.025 2.630 1.375 ;
        RECT  1.795 1.145 2.505 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.395 3.015 0.765 ;
        RECT  2.790 0.395 2.945 0.465 ;
        RECT  2.790 0.695 2.945 0.765 ;
        RECT  2.720 0.195 2.790 0.465 ;
        RECT  2.720 0.695 2.790 1.065 ;
        RECT  2.640 0.545 2.745 0.615 ;
        RECT  2.470 0.395 2.720 0.465 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.395 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  1.995 0.195 2.230 0.265 ;
        RECT  2.075 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.925 0.195 1.995 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  0.925 0.195 1.925 0.265 ;
        RECT  1.460 0.820 1.925 0.890 ;
        RECT  1.595 0.545 1.835 0.615 ;
        RECT  1.525 0.345 1.595 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.275 0.545 1.525 0.615 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.525 0.385 1.595 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.645 0.455 ;
    END
END DFQD2BWP40

MACRO DFQD4BWP40
    CLASS CORE ;
    FOREIGN DFQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.195 3.840 0.475 ;
        RECT  3.745 0.660 3.840 1.065 ;
        RECT  3.675 0.355 3.745 0.475 ;
        RECT  3.675 0.660 3.745 0.790 ;
        RECT  3.465 0.355 3.675 0.790 ;
        RECT  3.435 0.355 3.465 0.480 ;
        RECT  3.435 0.665 3.465 0.790 ;
        RECT  3.365 0.215 3.435 0.480 ;
        RECT  3.365 0.665 3.435 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.010 0.420 ;
        RECT  3.630 -0.115 3.935 0.115 ;
        RECT  3.550 -0.115 3.630 0.275 ;
        RECT  3.240 -0.115 3.550 0.115 ;
        RECT  3.170 -0.115 3.240 0.325 ;
        RECT  3.035 -0.115 3.170 0.115 ;
        RECT  2.965 -0.115 3.035 0.325 ;
        RECT  2.590 -0.115 2.965 0.115 ;
        RECT  2.520 -0.115 2.590 0.325 ;
        RECT  1.785 -0.115 2.520 0.115 ;
        RECT  1.665 -0.115 1.785 0.125 ;
        RECT  1.155 -0.115 1.665 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.935 0.685 4.010 1.375 ;
        RECT  3.645 1.145 3.935 1.375 ;
        RECT  3.535 0.905 3.645 1.375 ;
        RECT  3.240 1.145 3.535 1.375 ;
        RECT  3.170 0.845 3.240 1.375 ;
        RECT  3.035 1.145 3.170 1.375 ;
        RECT  2.965 0.845 3.035 1.375 ;
        RECT  2.595 1.145 2.965 1.375 ;
        RECT  2.465 1.130 2.595 1.375 ;
        RECT  1.745 1.145 2.465 1.375 ;
        RECT  1.675 0.980 1.745 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.745 0.195 3.840 0.475 ;
        RECT  3.745 0.660 3.840 1.065 ;
        RECT  3.365 0.215 3.395 0.480 ;
        RECT  3.365 0.665 3.395 1.065 ;
        RECT  3.195 0.405 3.265 0.765 ;
        RECT  2.780 0.405 3.195 0.475 ;
        RECT  2.780 0.695 3.195 0.765 ;
        RECT  2.630 0.545 2.915 0.615 ;
        RECT  2.710 0.195 2.780 0.475 ;
        RECT  2.710 0.695 2.780 1.030 ;
        RECT  2.470 0.405 2.710 0.475 ;
        RECT  2.560 0.545 2.630 0.910 ;
        RECT  2.115 0.840 2.560 0.910 ;
        RECT  2.400 0.405 2.470 0.580 ;
        RECT  2.255 0.690 2.365 0.760 ;
        RECT  2.185 0.195 2.255 0.760 ;
        RECT  2.085 0.195 2.185 0.265 ;
        RECT  2.045 0.345 2.115 0.910 ;
        RECT  1.975 0.185 2.085 0.265 ;
        RECT  1.935 0.185 1.975 0.890 ;
        RECT  1.905 0.195 1.935 0.890 ;
        RECT  0.925 0.195 1.905 0.265 ;
        RECT  1.460 0.820 1.905 0.890 ;
        RECT  1.755 0.345 1.825 0.635 ;
        RECT  1.275 0.545 1.755 0.615 ;
        RECT  1.405 0.985 1.525 1.075 ;
        RECT  0.340 0.985 1.405 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.755 0.385 1.825 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.875 0.455 ;
    END
END DFQD4BWP40

MACRO DFQND0BWP40
    CLASS CORE ;
    FOREIGN DFQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.195 3.185 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.970 0.315 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.735 -0.115 2.530 0.115 ;
        RECT  1.615 -0.115 1.735 0.125 ;
        RECT  1.155 -0.115 1.615 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.145 3.220 1.375 ;
        RECT  2.900 0.940 2.970 1.375 ;
        RECT  2.595 1.145 2.900 1.375 ;
        RECT  2.465 1.135 2.595 1.375 ;
        RECT  1.795 1.145 2.465 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.395 3.015 0.765 ;
        RECT  2.790 0.395 2.945 0.465 ;
        RECT  2.790 0.695 2.945 0.765 ;
        RECT  2.640 0.545 2.830 0.615 ;
        RECT  2.720 0.220 2.790 0.465 ;
        RECT  2.720 0.695 2.790 1.050 ;
        RECT  2.470 0.395 2.720 0.465 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.395 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  2.000 0.195 2.230 0.265 ;
        RECT  2.080 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.930 0.195 2.000 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  1.550 0.195 1.930 0.265 ;
        RECT  1.460 0.820 1.930 0.890 ;
        RECT  1.765 0.345 1.835 0.615 ;
        RECT  1.275 0.545 1.765 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.480 0.195 1.550 0.450 ;
        RECT  0.925 0.195 1.480 0.265 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.765 0.385 1.835 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.885 0.455 ;
    END
END DFQND0BWP40

MACRO DFQND1BWP40
    CLASS CORE ;
    FOREIGN DFQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.195 3.185 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.115 3.220 0.115 ;
        RECT  2.900 -0.115 2.970 0.315 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.785 -0.115 2.530 0.115 ;
        RECT  1.665 -0.115 1.785 0.125 ;
        RECT  1.155 -0.115 1.665 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.145 3.220 1.375 ;
        RECT  2.900 0.845 2.970 1.375 ;
        RECT  2.630 1.145 2.900 1.375 ;
        RECT  2.500 1.025 2.630 1.375 ;
        RECT  1.795 1.145 2.500 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.395 3.015 0.765 ;
        RECT  2.790 0.395 2.945 0.465 ;
        RECT  2.790 0.695 2.945 0.765 ;
        RECT  2.640 0.545 2.840 0.615 ;
        RECT  2.720 0.195 2.790 0.465 ;
        RECT  2.720 0.695 2.790 1.050 ;
        RECT  2.470 0.395 2.720 0.465 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.395 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  1.995 0.195 2.230 0.265 ;
        RECT  2.075 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.925 0.195 1.995 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  0.925 0.195 1.925 0.265 ;
        RECT  1.460 0.820 1.925 0.890 ;
        RECT  1.595 0.545 1.835 0.615 ;
        RECT  1.525 0.345 1.595 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.275 0.545 1.525 0.615 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.525 0.385 1.595 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.645 0.455 ;
    END
END DFQND1BWP40

MACRO DFQND2BWP40
    CLASS CORE ;
    FOREIGN DFQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.195 3.215 1.065 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.028000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.115 3.500 0.115 ;
        RECT  3.360 -0.115 3.445 0.485 ;
        RECT  2.970 -0.115 3.360 0.115 ;
        RECT  2.900 -0.115 2.970 0.325 ;
        RECT  2.600 -0.115 2.900 0.115 ;
        RECT  2.530 -0.115 2.600 0.315 ;
        RECT  1.785 -0.115 2.530 0.115 ;
        RECT  1.665 -0.115 1.785 0.125 ;
        RECT  1.155 -0.115 1.665 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.435 1.145 3.500 1.375 ;
        RECT  3.360 0.695 3.435 1.375 ;
        RECT  2.970 1.145 3.360 1.375 ;
        RECT  2.900 0.845 2.970 1.375 ;
        RECT  2.630 1.145 2.900 1.375 ;
        RECT  2.500 1.025 2.630 1.375 ;
        RECT  1.795 1.145 2.500 1.375 ;
        RECT  1.675 1.135 1.795 1.375 ;
        RECT  1.145 1.145 1.675 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.915 0.405 2.985 0.765 ;
        RECT  2.790 0.405 2.915 0.475 ;
        RECT  2.790 0.695 2.915 0.765 ;
        RECT  2.640 0.545 2.805 0.615 ;
        RECT  2.720 0.195 2.790 0.475 ;
        RECT  2.720 0.695 2.790 1.030 ;
        RECT  2.470 0.405 2.720 0.475 ;
        RECT  2.570 0.545 2.640 0.910 ;
        RECT  2.150 0.840 2.570 0.910 ;
        RECT  2.400 0.405 2.470 0.580 ;
        RECT  2.300 0.685 2.365 0.755 ;
        RECT  2.230 0.195 2.300 0.755 ;
        RECT  1.995 0.195 2.230 0.265 ;
        RECT  2.075 0.335 2.150 0.910 ;
        RECT  1.965 0.985 2.095 1.075 ;
        RECT  1.925 0.195 1.995 0.890 ;
        RECT  1.575 0.985 1.965 1.055 ;
        RECT  0.925 0.195 1.925 0.265 ;
        RECT  1.460 0.820 1.925 0.890 ;
        RECT  1.595 0.545 1.835 0.615 ;
        RECT  1.525 0.345 1.595 0.615 ;
        RECT  1.455 0.985 1.575 1.075 ;
        RECT  1.275 0.545 1.525 0.615 ;
        RECT  0.340 0.985 1.455 1.055 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.265 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.195 0.795 0.265 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.195 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.525 0.385 1.595 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.645 0.455 ;
    END
END DFQND2BWP40

MACRO DFQND4BWP40
    CLASS CORE ;
    FOREIGN DFQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.885 0.195 3.980 0.480 ;
        RECT  3.885 0.665 3.980 1.065 ;
        RECT  3.815 0.355 3.885 0.480 ;
        RECT  3.815 0.665 3.885 0.795 ;
        RECT  3.605 0.355 3.815 0.795 ;
        RECT  3.580 0.355 3.605 0.485 ;
        RECT  3.575 0.665 3.605 0.795 ;
        RECT  3.505 0.215 3.580 0.485 ;
        RECT  3.505 0.665 3.575 1.065 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.028800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.695 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.590 0.190 0.715 ;
        RECT  0.035 0.590 0.105 0.905 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 -0.115 4.200 0.115 ;
        RECT  4.070 -0.115 4.150 0.415 ;
        RECT  3.770 -0.115 4.070 0.115 ;
        RECT  3.695 -0.115 3.770 0.260 ;
        RECT  3.380 -0.115 3.695 0.115 ;
        RECT  3.310 -0.115 3.380 0.315 ;
        RECT  3.010 -0.115 3.310 0.115 ;
        RECT  2.940 -0.115 3.010 0.315 ;
        RECT  1.970 -0.115 2.940 0.115 ;
        RECT  1.840 -0.115 1.970 0.130 ;
        RECT  1.575 -0.115 1.840 0.115 ;
        RECT  1.455 -0.115 1.575 0.130 ;
        RECT  1.155 -0.115 1.455 0.115 ;
        RECT  1.025 -0.115 1.155 0.125 ;
        RECT  0.370 -0.115 1.025 0.115 ;
        RECT  0.250 -0.115 0.370 0.250 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.150 1.145 4.200 1.375 ;
        RECT  4.075 0.710 4.150 1.375 ;
        RECT  3.790 1.145 4.075 1.375 ;
        RECT  3.670 0.905 3.790 1.375 ;
        RECT  3.380 1.145 3.670 1.375 ;
        RECT  3.310 0.845 3.380 1.375 ;
        RECT  3.005 1.145 3.310 1.375 ;
        RECT  2.885 1.130 3.005 1.375 ;
        RECT  1.965 1.145 2.885 1.375 ;
        RECT  1.845 0.980 1.965 1.375 ;
        RECT  1.615 1.145 1.845 1.375 ;
        RECT  1.545 0.820 1.615 1.375 ;
        RECT  1.460 0.820 1.545 0.890 ;
        RECT  1.145 1.145 1.545 1.375 ;
        RECT  1.025 1.135 1.145 1.375 ;
        RECT  0.395 1.145 1.025 1.375 ;
        RECT  0.275 1.135 0.395 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.195 3.980 0.480 ;
        RECT  3.885 0.665 3.980 1.065 ;
        RECT  3.505 0.215 3.535 0.485 ;
        RECT  3.505 0.665 3.535 1.065 ;
        RECT  3.365 0.395 3.435 0.765 ;
        RECT  3.200 0.395 3.365 0.465 ;
        RECT  3.200 0.695 3.365 0.765 ;
        RECT  3.050 0.545 3.235 0.615 ;
        RECT  3.130 0.195 3.200 0.465 ;
        RECT  3.130 0.695 3.200 0.995 ;
        RECT  2.890 0.395 3.130 0.465 ;
        RECT  2.980 0.545 3.050 0.910 ;
        RECT  2.585 0.840 2.980 0.910 ;
        RECT  2.820 0.395 2.890 0.580 ;
        RECT  2.725 0.685 2.785 0.755 ;
        RECT  2.655 0.200 2.725 0.755 ;
        RECT  2.445 0.200 2.655 0.270 ;
        RECT  2.515 0.350 2.585 0.910 ;
        RECT  2.375 0.200 2.445 0.615 ;
        RECT  1.770 0.840 2.415 0.910 ;
        RECT  0.925 0.200 2.375 0.270 ;
        RECT  2.175 0.545 2.375 0.615 ;
        RECT  2.225 0.345 2.305 0.465 ;
        RECT  1.655 0.345 2.225 0.415 ;
        RECT  2.055 0.545 2.175 0.770 ;
        RECT  1.685 0.750 1.770 0.910 ;
        RECT  1.500 0.355 1.570 0.605 ;
        RECT  1.275 0.535 1.500 0.605 ;
        RECT  1.345 0.985 1.465 1.075 ;
        RECT  1.115 0.355 1.400 0.425 ;
        RECT  1.115 0.825 1.390 0.895 ;
        RECT  0.340 0.985 1.345 1.055 ;
        RECT  1.045 0.355 1.115 0.895 ;
        RECT  0.905 0.350 0.975 0.900 ;
        RECT  0.795 0.185 0.925 0.270 ;
        RECT  0.765 0.350 0.835 0.905 ;
        RECT  0.525 0.200 0.795 0.270 ;
        RECT  0.685 0.350 0.765 0.420 ;
        RECT  0.685 0.835 0.765 0.905 ;
        RECT  0.455 0.200 0.525 0.690 ;
        RECT  0.425 0.590 0.455 0.690 ;
        RECT  0.340 0.390 0.385 0.510 ;
        RECT  0.270 0.390 0.340 1.055 ;
        RECT  0.140 0.390 0.270 0.470 ;
        RECT  0.035 0.985 0.270 1.055 ;
        RECT  0.055 0.195 0.140 0.470 ;
        LAYER VIA1 ;
        RECT  1.500 0.385 1.570 0.455 ;
        RECT  0.765 0.385 0.835 0.455 ;
        LAYER M2 ;
        RECT  0.715 0.385 1.620 0.455 ;
    END
END DFQND4BWP40

MACRO DFSNQD0BWP40
    CLASS CORE ;
    FOREIGN DFSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 1.075 ;
        RECT  3.795 0.185 3.815 0.305 ;
        RECT  3.795 0.960 3.815 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.685 -0.115 3.920 0.115 ;
        RECT  3.595 -0.115 3.685 0.265 ;
        RECT  3.235 -0.115 3.595 0.115 ;
        RECT  3.135 -0.115 3.235 0.255 ;
        RECT  2.780 -0.115 3.135 0.115 ;
        RECT  2.710 -0.115 2.780 0.425 ;
        RECT  2.000 -0.115 2.710 0.115 ;
        RECT  1.930 -0.115 2.000 0.255 ;
        RECT  0.315 -0.115 1.930 0.115 ;
        RECT  0.245 -0.115 0.315 0.255 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 1.145 3.920 1.375 ;
        RECT  3.580 1.050 3.700 1.375 ;
        RECT  0.355 1.145 3.580 1.375 ;
        RECT  0.240 1.045 0.355 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.725 0.525 3.745 0.635 ;
        RECT  3.645 0.525 3.725 0.980 ;
        RECT  3.225 0.910 3.645 0.980 ;
        RECT  3.375 0.240 3.480 0.310 ;
        RECT  3.375 0.770 3.475 0.840 ;
        RECT  3.305 0.240 3.375 0.840 ;
        RECT  3.155 0.335 3.225 1.035 ;
        RECT  2.920 0.335 3.155 0.405 ;
        RECT  2.780 0.965 3.155 1.035 ;
        RECT  3.015 0.485 3.085 0.895 ;
        RECT  2.390 0.825 3.015 0.895 ;
        RECT  2.655 0.965 2.780 1.075 ;
        RECT  2.570 0.685 2.635 0.755 ;
        RECT  2.500 0.195 2.570 0.755 ;
        RECT  2.225 0.195 2.500 0.265 ;
        RECT  2.390 0.345 2.420 0.445 ;
        RECT  2.310 0.345 2.390 0.895 ;
        RECT  1.915 0.995 2.350 1.065 ;
        RECT  2.155 0.195 2.225 0.425 ;
        RECT  1.835 0.350 2.155 0.425 ;
        RECT  2.040 0.520 2.115 0.915 ;
        RECT  1.310 0.845 2.040 0.915 ;
        RECT  1.795 0.995 1.915 1.075 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.525 0.995 1.795 1.065 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.345 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.455 0.895 0.525 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.895 0.455 0.965 ;
        RECT  0.330 0.325 0.385 0.500 ;
        RECT  0.260 0.325 0.330 0.965 ;
        RECT  0.125 0.325 0.260 0.395 ;
        RECT  0.125 0.895 0.260 0.965 ;
        RECT  0.055 0.200 0.125 0.395 ;
        RECT  0.055 0.895 0.125 1.045 ;
    END
END DFSNQD0BWP40

MACRO DFSNQD1BWP40
    CLASS CORE ;
    FOREIGN DFSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.185 3.885 1.075 ;
        RECT  3.795 0.185 3.815 0.465 ;
        RECT  3.795 0.685 3.815 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.675 -0.115 3.920 0.115 ;
        RECT  3.605 -0.115 3.675 0.375 ;
        RECT  3.235 -0.115 3.605 0.115 ;
        RECT  3.135 -0.115 3.235 0.255 ;
        RECT  2.780 -0.115 3.135 0.115 ;
        RECT  2.710 -0.115 2.780 0.425 ;
        RECT  2.000 -0.115 2.710 0.115 ;
        RECT  1.930 -0.115 2.000 0.255 ;
        RECT  0.315 -0.115 1.930 0.115 ;
        RECT  0.245 -0.115 0.315 0.255 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 1.145 3.920 1.375 ;
        RECT  3.580 1.050 3.700 1.375 ;
        RECT  0.335 1.145 3.580 1.375 ;
        RECT  0.265 1.020 0.335 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.725 0.525 3.745 0.635 ;
        RECT  3.645 0.525 3.725 0.980 ;
        RECT  3.225 0.910 3.645 0.980 ;
        RECT  3.375 0.270 3.480 0.340 ;
        RECT  3.375 0.770 3.465 0.840 ;
        RECT  3.305 0.270 3.375 0.840 ;
        RECT  3.155 0.340 3.225 1.035 ;
        RECT  2.900 0.340 3.155 0.410 ;
        RECT  2.780 0.965 3.155 1.035 ;
        RECT  3.015 0.490 3.085 0.895 ;
        RECT  2.390 0.825 3.015 0.895 ;
        RECT  2.655 0.965 2.780 1.075 ;
        RECT  2.570 0.685 2.635 0.755 ;
        RECT  2.500 0.195 2.570 0.755 ;
        RECT  2.225 0.195 2.500 0.265 ;
        RECT  2.390 0.345 2.420 0.445 ;
        RECT  2.310 0.345 2.390 0.895 ;
        RECT  1.915 0.995 2.350 1.065 ;
        RECT  2.155 0.195 2.225 0.425 ;
        RECT  1.835 0.350 2.155 0.425 ;
        RECT  2.040 0.520 2.115 0.915 ;
        RECT  1.310 0.845 2.040 0.915 ;
        RECT  1.795 0.995 1.915 1.075 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.525 0.995 1.795 1.065 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.345 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.455 0.860 0.525 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.860 0.455 0.930 ;
        RECT  0.330 0.325 0.385 0.500 ;
        RECT  0.260 0.325 0.330 0.930 ;
        RECT  0.125 0.325 0.260 0.395 ;
        RECT  0.145 0.860 0.260 0.930 ;
        RECT  0.035 0.860 0.145 1.035 ;
        RECT  0.055 0.225 0.125 0.395 ;
    END
END DFSNQD1BWP40

MACRO DFSNQD2BWP40
    CLASS CORE ;
    FOREIGN DFSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.820 0.370 3.885 0.880 ;
        RECT  3.815 0.195 3.820 1.075 ;
        RECT  3.745 0.195 3.815 0.445 ;
        RECT  3.745 0.805 3.815 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.255 ;
        RECT  3.625 -0.115 3.935 0.115 ;
        RECT  3.555 -0.115 3.625 0.425 ;
        RECT  3.225 -0.115 3.555 0.115 ;
        RECT  3.135 -0.115 3.225 0.270 ;
        RECT  2.780 -0.115 3.135 0.115 ;
        RECT  2.710 -0.115 2.780 0.425 ;
        RECT  2.000 -0.115 2.710 0.115 ;
        RECT  1.930 -0.115 2.000 0.255 ;
        RECT  0.315 -0.115 1.930 0.115 ;
        RECT  0.245 -0.115 0.315 0.255 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.145 4.060 1.375 ;
        RECT  3.935 0.950 4.005 1.375 ;
        RECT  3.650 1.145 3.935 1.375 ;
        RECT  3.530 1.030 3.650 1.375 ;
        RECT  0.335 1.145 3.530 1.375 ;
        RECT  0.265 1.020 0.335 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.615 0.525 3.745 0.635 ;
        RECT  3.535 0.525 3.615 0.960 ;
        RECT  3.225 0.890 3.535 0.960 ;
        RECT  3.365 0.265 3.455 0.335 ;
        RECT  3.365 0.750 3.440 0.820 ;
        RECT  3.295 0.265 3.365 0.820 ;
        RECT  3.155 0.340 3.225 0.960 ;
        RECT  2.930 0.340 3.155 0.410 ;
        RECT  3.015 0.490 3.085 0.895 ;
        RECT  2.390 0.825 3.015 0.895 ;
        RECT  2.860 0.340 2.930 0.565 ;
        RECT  2.640 0.495 2.860 0.565 ;
        RECT  2.570 0.685 2.635 0.755 ;
        RECT  2.500 0.195 2.570 0.755 ;
        RECT  2.225 0.195 2.500 0.265 ;
        RECT  2.390 0.345 2.420 0.445 ;
        RECT  2.310 0.345 2.390 0.895 ;
        RECT  1.915 0.995 2.350 1.065 ;
        RECT  2.155 0.195 2.225 0.425 ;
        RECT  1.835 0.350 2.155 0.425 ;
        RECT  2.040 0.520 2.115 0.915 ;
        RECT  1.310 0.845 2.040 0.915 ;
        RECT  1.795 0.995 1.915 1.075 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.525 0.995 1.795 1.065 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.345 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.455 0.860 0.525 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.860 0.455 0.930 ;
        RECT  0.330 0.325 0.385 0.500 ;
        RECT  0.260 0.325 0.330 0.930 ;
        RECT  0.125 0.325 0.260 0.395 ;
        RECT  0.145 0.860 0.260 0.930 ;
        RECT  0.035 0.860 0.145 1.035 ;
        RECT  0.055 0.225 0.125 0.395 ;
    END
END DFSNQD2BWP40

MACRO DFSNQD4BWP40
    CLASS CORE ;
    FOREIGN DFSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.585 0.185 4.680 0.460 ;
        RECT  4.585 0.785 4.670 1.075 ;
        RECT  4.515 0.330 4.585 0.460 ;
        RECT  4.515 0.785 4.585 0.905 ;
        RECT  4.305 0.330 4.515 0.905 ;
        RECT  4.295 0.330 4.305 0.460 ;
        RECT  4.295 0.785 4.305 0.905 ;
        RECT  4.205 0.185 4.295 0.460 ;
        RECT  4.205 0.785 4.295 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.410 ;
        RECT  4.465 -0.115 4.775 0.115 ;
        RECT  4.395 -0.115 4.465 0.255 ;
        RECT  4.090 -0.115 4.395 0.115 ;
        RECT  4.015 -0.115 4.090 0.420 ;
        RECT  3.355 -0.115 4.015 0.115 ;
        RECT  3.225 -0.115 3.355 0.250 ;
        RECT  2.885 -0.115 3.225 0.115 ;
        RECT  2.815 -0.115 2.885 0.425 ;
        RECT  2.000 -0.115 2.815 0.115 ;
        RECT  1.930 -0.115 2.000 0.255 ;
        RECT  0.315 -0.115 1.930 0.115 ;
        RECT  0.245 -0.115 0.315 0.255 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.725 4.845 1.375 ;
        RECT  4.465 1.145 4.775 1.375 ;
        RECT  4.395 0.995 4.465 1.375 ;
        RECT  4.120 1.145 4.395 1.375 ;
        RECT  3.990 1.030 4.120 1.375 ;
        RECT  3.745 1.145 3.990 1.375 ;
        RECT  3.610 1.030 3.745 1.375 ;
        RECT  0.335 1.145 3.610 1.375 ;
        RECT  0.265 1.020 0.335 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.585 0.185 4.680 0.460 ;
        RECT  4.585 0.785 4.670 1.075 ;
        RECT  4.205 0.185 4.235 0.460 ;
        RECT  4.205 0.785 4.235 1.075 ;
        RECT  4.135 0.545 4.235 0.615 ;
        RECT  4.050 0.545 4.135 0.960 ;
        RECT  3.575 0.890 4.050 0.960 ;
        RECT  3.785 0.750 3.920 0.820 ;
        RECT  3.785 0.245 3.915 0.315 ;
        RECT  3.715 0.245 3.785 0.820 ;
        RECT  3.505 0.340 3.575 0.960 ;
        RECT  3.025 0.340 3.505 0.410 ;
        RECT  3.235 0.890 3.505 0.960 ;
        RECT  3.165 0.550 3.375 0.620 ;
        RECT  3.095 0.550 3.165 0.895 ;
        RECT  2.500 0.825 3.095 0.895 ;
        RECT  2.955 0.340 3.025 0.575 ;
        RECT  2.750 0.505 2.955 0.575 ;
        RECT  2.680 0.685 2.740 0.755 ;
        RECT  2.610 0.195 2.680 0.755 ;
        RECT  2.295 0.195 2.610 0.265 ;
        RECT  2.415 0.345 2.500 0.895 ;
        RECT  1.915 0.995 2.455 1.065 ;
        RECT  2.225 0.195 2.295 0.425 ;
        RECT  1.835 0.350 2.225 0.425 ;
        RECT  2.090 0.520 2.165 0.915 ;
        RECT  1.310 0.845 2.090 0.915 ;
        RECT  1.795 0.995 1.915 1.075 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.525 0.995 1.795 1.065 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.340 0.345 1.380 0.415 ;
        RECT  1.150 0.335 1.340 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.335 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.455 0.860 0.525 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.860 0.455 0.930 ;
        RECT  0.330 0.325 0.385 0.500 ;
        RECT  0.260 0.325 0.330 0.930 ;
        RECT  0.125 0.325 0.260 0.395 ;
        RECT  0.140 0.860 0.260 0.930 ;
        RECT  0.035 0.860 0.140 1.030 ;
        RECT  0.055 0.225 0.125 0.395 ;
    END
END DFSNQD4BWP40

MACRO DFSNQND0BWP40
    CLASS CORE ;
    FOREIGN DFSNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.075 ;
        RECT  3.935 0.185 3.955 0.310 ;
        RECT  3.935 0.950 3.955 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.840 -0.115 4.060 0.115 ;
        RECT  3.720 -0.115 3.840 0.180 ;
        RECT  3.425 -0.115 3.720 0.115 ;
        RECT  3.305 -0.115 3.425 0.210 ;
        RECT  3.005 -0.115 3.305 0.115 ;
        RECT  2.865 -0.115 3.005 0.210 ;
        RECT  2.060 -0.115 2.865 0.115 ;
        RECT  1.990 -0.115 2.060 0.255 ;
        RECT  0.320 -0.115 1.990 0.115 ;
        RECT  0.240 -0.115 0.320 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.825 1.145 4.060 1.375 ;
        RECT  3.735 0.860 3.825 1.375 ;
        RECT  3.045 1.145 3.735 1.375 ;
        RECT  2.905 1.060 3.045 1.375 ;
        RECT  0.340 1.145 2.905 1.375 ;
        RECT  0.260 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.795 0.525 3.885 0.635 ;
        RECT  3.720 0.280 3.795 0.635 ;
        RECT  2.905 0.280 3.720 0.350 ;
        RECT  3.410 0.420 3.630 0.495 ;
        RECT  3.535 0.795 3.625 0.865 ;
        RECT  3.395 0.970 3.570 1.040 ;
        RECT  3.465 0.650 3.535 0.865 ;
        RECT  3.410 0.650 3.465 0.720 ;
        RECT  3.340 0.420 3.410 0.720 ;
        RECT  3.325 0.800 3.395 1.040 ;
        RECT  3.270 0.800 3.325 0.870 ;
        RECT  3.200 0.430 3.270 0.870 ;
        RECT  3.075 0.430 3.200 0.500 ;
        RECT  3.050 0.645 3.120 0.990 ;
        RECT  2.635 0.920 3.050 0.990 ;
        RECT  2.835 0.280 2.905 0.850 ;
        RECT  2.725 0.280 2.835 0.415 ;
        RECT  2.720 0.780 2.835 0.850 ;
        RECT  2.655 0.625 2.735 0.695 ;
        RECT  2.585 0.195 2.655 0.695 ;
        RECT  2.565 0.855 2.635 0.990 ;
        RECT  2.230 0.195 2.585 0.265 ;
        RECT  2.475 0.855 2.565 0.925 ;
        RECT  2.475 0.335 2.515 0.450 ;
        RECT  1.960 0.995 2.485 1.065 ;
        RECT  2.385 0.335 2.475 0.925 ;
        RECT  2.160 0.195 2.230 0.425 ;
        RECT  2.125 0.520 2.215 0.915 ;
        RECT  1.835 0.350 2.160 0.425 ;
        RECT  1.310 0.845 2.125 0.915 ;
        RECT  1.840 0.995 1.960 1.075 ;
        RECT  0.520 0.995 1.840 1.065 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.345 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.450 0.845 0.520 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.845 0.450 0.915 ;
        RECT  0.330 0.340 0.385 0.500 ;
        RECT  0.260 0.340 0.330 0.915 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.130 0.845 0.260 0.915 ;
        RECT  0.055 0.845 0.130 1.045 ;
        RECT  0.055 0.200 0.125 0.410 ;
    END
END DFSNQND0BWP40

MACRO DFSNQND1BWP40
    CLASS CORE ;
    FOREIGN DFSNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.185 4.025 1.075 ;
        RECT  3.935 0.185 3.955 0.465 ;
        RECT  3.935 0.685 3.955 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.825 -0.115 4.060 0.115 ;
        RECT  3.705 -0.115 3.825 0.210 ;
        RECT  3.425 -0.115 3.705 0.115 ;
        RECT  3.305 -0.115 3.425 0.210 ;
        RECT  3.005 -0.115 3.305 0.115 ;
        RECT  2.865 -0.115 3.005 0.210 ;
        RECT  2.060 -0.115 2.865 0.115 ;
        RECT  1.990 -0.115 2.060 0.255 ;
        RECT  0.320 -0.115 1.990 0.115 ;
        RECT  0.240 -0.115 0.320 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.745 3.815 1.375 ;
        RECT  3.045 1.145 3.745 1.375 ;
        RECT  2.905 1.060 3.045 1.375 ;
        RECT  0.340 1.145 2.905 1.375 ;
        RECT  0.260 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.795 0.525 3.885 0.635 ;
        RECT  3.720 0.280 3.795 0.635 ;
        RECT  2.905 0.280 3.720 0.350 ;
        RECT  3.410 0.420 3.625 0.495 ;
        RECT  3.535 0.795 3.625 0.865 ;
        RECT  3.395 0.970 3.570 1.040 ;
        RECT  3.465 0.650 3.535 0.865 ;
        RECT  3.410 0.650 3.465 0.720 ;
        RECT  3.340 0.420 3.410 0.720 ;
        RECT  3.325 0.800 3.395 1.040 ;
        RECT  3.270 0.800 3.325 0.870 ;
        RECT  3.200 0.430 3.270 0.870 ;
        RECT  3.075 0.430 3.200 0.500 ;
        RECT  3.050 0.645 3.120 0.990 ;
        RECT  2.635 0.920 3.050 0.990 ;
        RECT  2.835 0.280 2.905 0.850 ;
        RECT  2.725 0.280 2.835 0.415 ;
        RECT  2.720 0.780 2.835 0.850 ;
        RECT  2.655 0.625 2.740 0.695 ;
        RECT  2.585 0.195 2.655 0.695 ;
        RECT  2.565 0.855 2.635 0.990 ;
        RECT  2.230 0.195 2.585 0.265 ;
        RECT  2.475 0.855 2.565 0.925 ;
        RECT  2.475 0.335 2.515 0.450 ;
        RECT  1.960 0.995 2.485 1.065 ;
        RECT  2.395 0.335 2.475 0.925 ;
        RECT  2.160 0.195 2.230 0.425 ;
        RECT  2.125 0.520 2.215 0.915 ;
        RECT  1.835 0.350 2.160 0.425 ;
        RECT  1.310 0.845 2.125 0.915 ;
        RECT  1.840 0.995 1.960 1.075 ;
        RECT  0.520 0.995 1.840 1.065 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.150 0.345 1.380 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.345 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.525 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.455 0.195 0.525 0.700 ;
        RECT  0.450 0.845 0.520 1.065 ;
        RECT  0.400 0.580 0.455 0.700 ;
        RECT  0.330 0.845 0.450 0.915 ;
        RECT  0.330 0.340 0.385 0.500 ;
        RECT  0.260 0.340 0.330 0.915 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.140 0.845 0.260 0.915 ;
        RECT  0.035 0.845 0.140 1.030 ;
        RECT  0.055 0.210 0.125 0.410 ;
    END
END DFSNQND1BWP40

MACRO DFSNQND2BWP40
    CLASS CORE ;
    FOREIGN DFSNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 0.370 4.025 0.880 ;
        RECT  3.955 0.195 3.960 1.075 ;
        RECT  3.885 0.195 3.955 0.445 ;
        RECT  3.885 0.805 3.955 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 -0.115 4.200 0.115 ;
        RECT  4.075 -0.115 4.145 0.275 ;
        RECT  3.790 -0.115 4.075 0.115 ;
        RECT  3.670 -0.115 3.790 0.180 ;
        RECT  3.395 -0.115 3.670 0.115 ;
        RECT  3.275 -0.115 3.395 0.210 ;
        RECT  3.005 -0.115 3.275 0.115 ;
        RECT  2.865 -0.115 3.005 0.210 ;
        RECT  2.060 -0.115 2.865 0.115 ;
        RECT  1.990 -0.115 2.060 0.255 ;
        RECT  0.320 -0.115 1.990 0.115 ;
        RECT  0.240 -0.115 0.320 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.145 1.145 4.200 1.375 ;
        RECT  4.075 0.950 4.145 1.375 ;
        RECT  3.765 1.145 4.075 1.375 ;
        RECT  3.695 0.725 3.765 1.375 ;
        RECT  3.040 1.145 3.695 1.375 ;
        RECT  2.905 1.060 3.040 1.375 ;
        RECT  0.340 1.145 2.905 1.375 ;
        RECT  0.260 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.795 0.525 3.885 0.635 ;
        RECT  3.720 0.280 3.795 0.635 ;
        RECT  2.905 0.280 3.720 0.350 ;
        RECT  3.530 0.795 3.625 0.865 ;
        RECT  3.380 0.420 3.595 0.495 ;
        RECT  3.390 0.990 3.540 1.060 ;
        RECT  3.460 0.620 3.530 0.865 ;
        RECT  3.380 0.620 3.460 0.700 ;
        RECT  3.320 0.800 3.390 1.060 ;
        RECT  3.310 0.420 3.380 0.700 ;
        RECT  3.240 0.800 3.320 0.870 ;
        RECT  3.170 0.430 3.240 0.870 ;
        RECT  3.075 0.430 3.170 0.500 ;
        RECT  3.020 0.645 3.090 0.990 ;
        RECT  2.635 0.920 3.020 0.990 ;
        RECT  2.835 0.280 2.905 0.850 ;
        RECT  2.725 0.280 2.835 0.415 ;
        RECT  2.715 0.780 2.835 0.850 ;
        RECT  2.655 0.625 2.740 0.695 ;
        RECT  2.585 0.195 2.655 0.695 ;
        RECT  2.565 0.855 2.635 0.990 ;
        RECT  2.230 0.195 2.585 0.265 ;
        RECT  2.475 0.855 2.565 0.925 ;
        RECT  2.475 0.335 2.515 0.450 ;
        RECT  1.960 0.995 2.485 1.065 ;
        RECT  2.385 0.335 2.475 0.925 ;
        RECT  2.160 0.195 2.230 0.425 ;
        RECT  2.120 0.520 2.210 0.915 ;
        RECT  1.835 0.350 2.160 0.425 ;
        RECT  1.310 0.845 2.120 0.915 ;
        RECT  1.840 0.995 1.960 1.075 ;
        RECT  0.520 0.995 1.840 1.065 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.340 0.345 1.380 0.415 ;
        RECT  1.150 0.335 1.340 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.335 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.520 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.450 0.195 0.520 0.700 ;
        RECT  0.450 0.845 0.520 1.065 ;
        RECT  0.400 0.580 0.450 0.700 ;
        RECT  0.330 0.845 0.450 0.915 ;
        RECT  0.330 0.340 0.380 0.500 ;
        RECT  0.260 0.340 0.330 0.915 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.140 0.845 0.260 0.915 ;
        RECT  0.035 0.845 0.140 1.030 ;
        RECT  0.055 0.210 0.125 0.410 ;
    END
END DFSNQND2BWP40

MACRO DFSNQND4BWP40
    CLASS CORE ;
    FOREIGN DFSNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.525 1.675 0.765 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.190 4.820 0.440 ;
        RECT  4.725 0.745 4.820 1.005 ;
        RECT  4.655 0.355 4.725 0.440 ;
        RECT  4.655 0.745 4.725 0.830 ;
        RECT  4.445 0.355 4.655 0.830 ;
        RECT  4.420 0.355 4.445 0.475 ;
        RECT  4.420 0.710 4.445 0.830 ;
        RECT  4.350 0.205 4.420 0.475 ;
        RECT  4.350 0.710 4.420 1.020 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.029600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.495 0.685 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.430 ;
        RECT  4.610 -0.115 4.910 0.115 ;
        RECT  4.535 -0.115 4.610 0.270 ;
        RECT  4.250 -0.115 4.535 0.115 ;
        RECT  4.130 -0.115 4.250 0.210 ;
        RECT  3.860 -0.115 4.130 0.115 ;
        RECT  3.740 -0.115 3.860 0.210 ;
        RECT  3.445 -0.115 3.740 0.115 ;
        RECT  3.320 -0.115 3.445 0.210 ;
        RECT  3.075 -0.115 3.320 0.115 ;
        RECT  2.950 -0.115 3.075 0.210 ;
        RECT  2.060 -0.115 2.950 0.115 ;
        RECT  1.990 -0.115 2.060 0.255 ;
        RECT  0.320 -0.115 1.990 0.115 ;
        RECT  0.240 -0.115 0.320 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.900 0.705 4.990 1.375 ;
        RECT  4.625 1.145 4.900 1.375 ;
        RECT  4.515 0.905 4.625 1.375 ;
        RECT  4.230 1.145 4.515 1.375 ;
        RECT  4.155 0.720 4.230 1.375 ;
        RECT  3.485 1.145 4.155 1.375 ;
        RECT  3.355 1.050 3.485 1.375 ;
        RECT  3.090 1.145 3.355 1.375 ;
        RECT  2.950 1.050 3.090 1.375 ;
        RECT  0.340 1.145 2.950 1.375 ;
        RECT  0.260 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.190 4.820 0.440 ;
        RECT  4.725 0.745 4.820 1.005 ;
        RECT  4.350 0.205 4.375 0.475 ;
        RECT  4.350 0.710 4.375 1.020 ;
        RECT  4.215 0.545 4.365 0.620 ;
        RECT  4.140 0.280 4.215 0.620 ;
        RECT  3.265 0.280 4.140 0.350 ;
        RECT  3.830 0.420 4.060 0.495 ;
        RECT  4.010 1.005 4.055 1.075 ;
        RECT  3.940 0.720 4.010 1.075 ;
        RECT  3.830 0.720 3.940 0.790 ;
        RECT  3.690 0.970 3.860 1.040 ;
        RECT  3.760 0.420 3.830 0.790 ;
        RECT  3.620 0.430 3.690 1.040 ;
        RECT  3.405 0.430 3.620 0.500 ;
        RECT  3.470 0.645 3.540 0.980 ;
        RECT  2.665 0.910 3.470 0.980 ;
        RECT  3.335 0.430 3.405 0.565 ;
        RECT  3.070 0.495 3.335 0.565 ;
        RECT  2.920 0.770 3.280 0.840 ;
        RECT  3.145 0.280 3.265 0.400 ;
        RECT  2.920 0.280 3.145 0.350 ;
        RECT  3.000 0.495 3.070 0.645 ;
        RECT  2.850 0.280 2.920 0.840 ;
        RECT  2.780 0.280 2.850 0.415 ;
        RECT  2.765 0.770 2.850 0.840 ;
        RECT  2.680 0.625 2.770 0.695 ;
        RECT  2.610 0.195 2.680 0.695 ;
        RECT  2.595 0.855 2.665 0.980 ;
        RECT  2.230 0.195 2.610 0.265 ;
        RECT  2.530 0.855 2.595 0.925 ;
        RECT  2.460 0.335 2.530 0.925 ;
        RECT  1.960 0.995 2.480 1.065 ;
        RECT  2.160 0.195 2.230 0.425 ;
        RECT  2.125 0.520 2.215 0.915 ;
        RECT  1.835 0.350 2.160 0.425 ;
        RECT  1.310 0.845 2.125 0.915 ;
        RECT  1.840 0.995 1.960 1.075 ;
        RECT  0.520 0.995 1.840 1.065 ;
        RECT  1.815 0.350 1.835 0.775 ;
        RECT  1.745 0.195 1.815 0.775 ;
        RECT  0.935 0.195 1.745 0.265 ;
        RECT  1.470 0.345 1.610 0.455 ;
        RECT  1.380 0.345 1.470 0.775 ;
        RECT  1.340 0.345 1.380 0.415 ;
        RECT  1.150 0.335 1.340 0.415 ;
        RECT  1.240 0.510 1.310 0.915 ;
        RECT  0.825 0.845 1.240 0.915 ;
        RECT  1.070 0.335 1.150 0.625 ;
        RECT  1.035 0.535 1.070 0.625 ;
        RECT  0.965 0.700 1.040 0.770 ;
        RECT  0.965 0.350 0.985 0.470 ;
        RECT  0.895 0.350 0.965 0.770 ;
        RECT  0.810 0.185 0.935 0.265 ;
        RECT  0.755 0.335 0.825 0.915 ;
        RECT  0.520 0.195 0.810 0.265 ;
        RECT  0.630 0.335 0.755 0.405 ;
        RECT  0.610 0.845 0.755 0.915 ;
        RECT  0.450 0.195 0.520 0.700 ;
        RECT  0.450 0.845 0.520 1.065 ;
        RECT  0.400 0.580 0.450 0.700 ;
        RECT  0.330 0.845 0.450 0.915 ;
        RECT  0.330 0.340 0.380 0.500 ;
        RECT  0.260 0.340 0.330 0.915 ;
        RECT  0.125 0.340 0.260 0.410 ;
        RECT  0.140 0.845 0.260 0.915 ;
        RECT  0.035 0.845 0.140 1.040 ;
        RECT  0.055 0.210 0.125 0.410 ;
    END
END DFSNQND4BWP40

MACRO EDFCNQD0BWP40
    CLASS CORE ;
    FOREIGN EDFCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.075 ;
        RECT  4.635 0.185 4.655 0.295 ;
        RECT  4.635 0.905 4.655 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.021400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.410 0.625 ;
        RECT  0.940 0.355 1.135 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.385 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.510 -0.115 4.760 0.115 ;
        RECT  4.390 -0.115 4.510 0.255 ;
        RECT  3.940 -0.115 4.390 0.115 ;
        RECT  3.815 -0.115 3.940 0.245 ;
        RECT  3.100 -0.115 3.815 0.115 ;
        RECT  2.980 -0.115 3.100 0.195 ;
        RECT  1.520 -0.115 2.980 0.115 ;
        RECT  1.400 -0.115 1.520 0.125 ;
        RECT  1.190 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.315 -0.115 1.070 0.115 ;
        RECT  0.245 -0.115 0.315 0.330 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.145 4.760 1.375 ;
        RECT  4.410 1.025 4.530 1.375 ;
        RECT  4.060 1.145 4.410 1.375 ;
        RECT  3.940 1.040 4.060 1.375 ;
        RECT  3.100 1.145 3.940 1.375 ;
        RECT  2.980 1.070 3.100 1.375 ;
        RECT  2.490 1.145 2.980 1.375 ;
        RECT  2.365 1.070 2.490 1.375 ;
        RECT  1.540 1.145 2.365 1.375 ;
        RECT  1.420 1.135 1.540 1.375 ;
        RECT  1.170 1.145 1.420 1.375 ;
        RECT  1.050 1.135 1.170 1.375 ;
        RECT  0.340 1.145 1.050 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.480 0.325 4.550 0.920 ;
        RECT  3.870 0.325 4.480 0.395 ;
        RECT  4.310 0.850 4.480 0.920 ;
        RECT  4.190 0.850 4.310 0.995 ;
        RECT  4.070 0.510 4.165 0.630 ;
        RECT  4.000 0.510 4.070 0.910 ;
        RECT  3.460 0.840 4.000 0.910 ;
        RECT  3.800 0.325 3.870 0.595 ;
        RECT  3.685 0.685 3.755 0.765 ;
        RECT  3.615 0.195 3.685 0.765 ;
        RECT  3.260 0.195 3.615 0.265 ;
        RECT  3.390 0.345 3.460 1.000 ;
        RECT  2.090 0.930 3.390 1.000 ;
        RECT  3.190 0.195 3.260 0.335 ;
        RECT  3.155 0.405 3.230 0.860 ;
        RECT  2.900 0.265 3.190 0.335 ;
        RECT  2.750 0.405 3.155 0.475 ;
        RECT  2.775 0.780 3.155 0.860 ;
        RECT  2.595 0.610 3.055 0.690 ;
        RECT  2.830 0.195 2.900 0.335 ;
        RECT  2.095 0.195 2.830 0.265 ;
        RECT  2.680 0.335 2.750 0.475 ;
        RECT  2.280 0.780 2.695 0.850 ;
        RECT  2.420 0.335 2.680 0.405 ;
        RECT  2.515 0.495 2.595 0.690 ;
        RECT  2.350 0.335 2.420 0.625 ;
        RECT  2.210 0.345 2.280 0.850 ;
        RECT  2.065 0.345 2.135 0.780 ;
        RECT  2.020 0.850 2.090 1.000 ;
        RECT  1.995 0.345 2.065 0.425 ;
        RECT  2.010 0.710 2.065 0.780 ;
        RECT  1.070 0.850 2.020 0.920 ;
        RECT  1.855 0.530 1.990 0.640 ;
        RECT  0.650 0.195 1.950 0.265 ;
        RECT  1.810 0.995 1.940 1.075 ;
        RECT  1.785 0.345 1.855 0.770 ;
        RECT  0.640 0.995 1.810 1.065 ;
        RECT  1.645 0.345 1.785 0.465 ;
        RECT  1.640 0.700 1.785 0.770 ;
        RECT  1.550 0.545 1.660 0.615 ;
        RECT  1.480 0.335 1.550 0.780 ;
        RECT  1.220 0.335 1.480 0.405 ;
        RECT  1.200 0.710 1.480 0.780 ;
        RECT  0.940 0.700 1.070 0.920 ;
        RECT  0.765 0.490 0.850 0.920 ;
        RECT  0.140 0.850 0.765 0.920 ;
        RECT  0.625 0.345 0.695 0.780 ;
        RECT  0.415 0.345 0.625 0.415 ;
        RECT  0.430 0.710 0.625 0.780 ;
        RECT  0.105 0.850 0.140 1.070 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.035 0.210 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.520 0.525 2.590 0.595 ;
        RECT  2.065 0.525 2.135 0.595 ;
        LAYER M2 ;
        RECT  2.015 0.525 2.640 0.595 ;
    END
END EDFCNQD0BWP40

MACRO EDFCNQD1BWP40
    CLASS CORE ;
    FOREIGN EDFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.088550 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.185 4.725 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.022000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.410 0.625 ;
        RECT  0.940 0.355 1.135 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.040400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.385 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.510 -0.115 4.760 0.115 ;
        RECT  4.390 -0.115 4.510 0.240 ;
        RECT  3.940 -0.115 4.390 0.115 ;
        RECT  3.815 -0.115 3.940 0.245 ;
        RECT  3.100 -0.115 3.815 0.115 ;
        RECT  2.980 -0.115 3.100 0.195 ;
        RECT  1.520 -0.115 2.980 0.115 ;
        RECT  1.400 -0.115 1.520 0.125 ;
        RECT  1.190 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.315 -0.115 1.070 0.115 ;
        RECT  0.245 -0.115 0.315 0.330 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.145 4.760 1.375 ;
        RECT  4.410 1.025 4.530 1.375 ;
        RECT  4.060 1.145 4.410 1.375 ;
        RECT  3.940 1.040 4.060 1.375 ;
        RECT  3.100 1.145 3.940 1.375 ;
        RECT  2.980 1.070 3.100 1.375 ;
        RECT  2.490 1.145 2.980 1.375 ;
        RECT  2.365 1.070 2.490 1.375 ;
        RECT  1.540 1.145 2.365 1.375 ;
        RECT  1.420 1.135 1.540 1.375 ;
        RECT  1.170 1.145 1.420 1.375 ;
        RECT  1.050 1.135 1.170 1.375 ;
        RECT  0.340 1.145 1.050 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.480 0.320 4.550 0.920 ;
        RECT  3.870 0.320 4.480 0.390 ;
        RECT  4.190 0.850 4.480 0.920 ;
        RECT  4.070 0.510 4.165 0.630 ;
        RECT  4.000 0.510 4.070 0.910 ;
        RECT  3.460 0.840 4.000 0.910 ;
        RECT  3.800 0.320 3.870 0.595 ;
        RECT  3.685 0.685 3.755 0.765 ;
        RECT  3.615 0.195 3.685 0.765 ;
        RECT  3.260 0.195 3.615 0.265 ;
        RECT  3.390 0.345 3.460 1.000 ;
        RECT  2.090 0.930 3.390 1.000 ;
        RECT  3.190 0.195 3.260 0.335 ;
        RECT  3.155 0.405 3.230 0.860 ;
        RECT  2.900 0.265 3.190 0.335 ;
        RECT  2.750 0.405 3.155 0.475 ;
        RECT  2.775 0.780 3.155 0.860 ;
        RECT  2.595 0.610 3.055 0.690 ;
        RECT  2.830 0.195 2.900 0.335 ;
        RECT  2.095 0.195 2.830 0.265 ;
        RECT  2.680 0.335 2.750 0.475 ;
        RECT  2.280 0.780 2.695 0.850 ;
        RECT  2.420 0.335 2.680 0.405 ;
        RECT  2.515 0.495 2.595 0.690 ;
        RECT  2.350 0.335 2.420 0.625 ;
        RECT  2.210 0.345 2.280 0.850 ;
        RECT  2.065 0.345 2.135 0.780 ;
        RECT  2.020 0.850 2.090 1.000 ;
        RECT  1.995 0.345 2.065 0.425 ;
        RECT  2.010 0.710 2.065 0.780 ;
        RECT  1.070 0.850 2.020 0.920 ;
        RECT  1.855 0.530 1.990 0.640 ;
        RECT  0.650 0.195 1.950 0.265 ;
        RECT  1.810 0.995 1.940 1.075 ;
        RECT  1.785 0.345 1.855 0.770 ;
        RECT  0.640 0.995 1.810 1.065 ;
        RECT  1.645 0.345 1.785 0.465 ;
        RECT  1.640 0.700 1.785 0.770 ;
        RECT  1.550 0.545 1.660 0.615 ;
        RECT  1.480 0.335 1.550 0.780 ;
        RECT  1.220 0.335 1.480 0.405 ;
        RECT  1.200 0.710 1.480 0.780 ;
        RECT  0.940 0.700 1.070 0.920 ;
        RECT  0.765 0.490 0.850 0.920 ;
        RECT  0.140 0.850 0.765 0.920 ;
        RECT  0.625 0.345 0.695 0.780 ;
        RECT  0.415 0.345 0.625 0.415 ;
        RECT  0.430 0.710 0.625 0.780 ;
        RECT  0.105 0.850 0.140 1.070 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.035 0.210 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.520 0.525 2.590 0.595 ;
        RECT  2.065 0.525 2.135 0.595 ;
        LAYER M2 ;
        RECT  2.015 0.525 2.640 0.595 ;
    END
END EDFCNQD1BWP40

MACRO EDFCNQD2BWP40
    CLASS CORE ;
    FOREIGN EDFCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.150150 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.185 4.725 1.075 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.022000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.410 0.625 ;
        RECT  0.940 0.355 1.135 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.040400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.385 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.965 -0.115 5.040 0.115 ;
        RECT  4.885 -0.115 4.965 0.500 ;
        RECT  4.510 -0.115 4.885 0.115 ;
        RECT  4.390 -0.115 4.510 0.240 ;
        RECT  3.940 -0.115 4.390 0.115 ;
        RECT  3.815 -0.115 3.940 0.245 ;
        RECT  3.100 -0.115 3.815 0.115 ;
        RECT  2.980 -0.115 3.100 0.195 ;
        RECT  1.520 -0.115 2.980 0.115 ;
        RECT  1.400 -0.115 1.520 0.125 ;
        RECT  1.190 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.315 -0.115 1.070 0.115 ;
        RECT  0.245 -0.115 0.315 0.330 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.965 1.145 5.040 1.375 ;
        RECT  4.885 0.665 4.965 1.375 ;
        RECT  4.530 1.145 4.885 1.375 ;
        RECT  4.410 1.025 4.530 1.375 ;
        RECT  4.060 1.145 4.410 1.375 ;
        RECT  3.940 1.040 4.060 1.375 ;
        RECT  3.100 1.145 3.940 1.375 ;
        RECT  2.980 1.070 3.100 1.375 ;
        RECT  2.490 1.145 2.980 1.375 ;
        RECT  2.365 1.070 2.490 1.375 ;
        RECT  1.540 1.145 2.365 1.375 ;
        RECT  1.420 1.135 1.540 1.375 ;
        RECT  1.170 1.145 1.420 1.375 ;
        RECT  1.050 1.135 1.170 1.375 ;
        RECT  0.340 1.145 1.050 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.480 0.320 4.550 0.920 ;
        RECT  3.870 0.320 4.480 0.390 ;
        RECT  4.190 0.850 4.480 0.920 ;
        RECT  4.070 0.510 4.165 0.630 ;
        RECT  4.000 0.510 4.070 0.910 ;
        RECT  3.460 0.840 4.000 0.910 ;
        RECT  3.800 0.320 3.870 0.595 ;
        RECT  3.685 0.685 3.755 0.765 ;
        RECT  3.615 0.195 3.685 0.765 ;
        RECT  3.260 0.195 3.615 0.265 ;
        RECT  3.390 0.345 3.460 1.000 ;
        RECT  2.090 0.930 3.390 1.000 ;
        RECT  3.190 0.195 3.260 0.335 ;
        RECT  3.155 0.405 3.230 0.860 ;
        RECT  2.900 0.265 3.190 0.335 ;
        RECT  2.750 0.405 3.155 0.475 ;
        RECT  2.775 0.780 3.155 0.860 ;
        RECT  2.595 0.610 3.055 0.690 ;
        RECT  2.830 0.195 2.900 0.335 ;
        RECT  2.095 0.195 2.830 0.265 ;
        RECT  2.680 0.335 2.750 0.475 ;
        RECT  2.280 0.780 2.695 0.850 ;
        RECT  2.420 0.335 2.680 0.405 ;
        RECT  2.515 0.495 2.595 0.690 ;
        RECT  2.350 0.335 2.420 0.625 ;
        RECT  2.210 0.345 2.280 0.850 ;
        RECT  2.065 0.345 2.135 0.780 ;
        RECT  2.020 0.850 2.090 1.000 ;
        RECT  1.995 0.345 2.065 0.425 ;
        RECT  2.010 0.710 2.065 0.780 ;
        RECT  1.070 0.850 2.020 0.920 ;
        RECT  1.855 0.530 1.990 0.640 ;
        RECT  0.650 0.195 1.950 0.265 ;
        RECT  1.810 0.995 1.940 1.075 ;
        RECT  1.785 0.345 1.855 0.770 ;
        RECT  0.640 0.995 1.810 1.065 ;
        RECT  1.645 0.345 1.785 0.465 ;
        RECT  1.640 0.700 1.785 0.770 ;
        RECT  1.550 0.545 1.660 0.615 ;
        RECT  1.480 0.335 1.550 0.780 ;
        RECT  1.220 0.335 1.480 0.405 ;
        RECT  1.200 0.710 1.480 0.780 ;
        RECT  0.940 0.700 1.070 0.920 ;
        RECT  0.765 0.490 0.850 0.920 ;
        RECT  0.140 0.850 0.765 0.920 ;
        RECT  0.625 0.345 0.695 0.780 ;
        RECT  0.415 0.345 0.625 0.415 ;
        RECT  0.430 0.710 0.625 0.780 ;
        RECT  0.105 0.850 0.140 1.070 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.035 0.210 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.520 0.525 2.590 0.595 ;
        RECT  2.065 0.525 2.135 0.595 ;
        LAYER M2 ;
        RECT  2.015 0.525 2.640 0.595 ;
    END
END EDFCNQD2BWP40

MACRO EDFCNQD4BWP40
    CLASS CORE ;
    FOREIGN EDFCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.237000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.195 5.380 0.475 ;
        RECT  5.285 0.710 5.380 1.010 ;
        RECT  5.215 0.355 5.285 0.475 ;
        RECT  5.215 0.710 5.285 0.830 ;
        RECT  5.005 0.355 5.215 0.830 ;
        RECT  4.980 0.355 5.005 0.475 ;
        RECT  4.980 0.710 5.005 0.830 ;
        RECT  4.910 0.195 4.980 0.475 ;
        RECT  4.910 0.710 4.980 1.010 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.022000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.410 0.625 ;
        RECT  0.940 0.355 1.135 0.625 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.047600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.505 0.495 4.655 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.545 0.450 ;
        RECT  5.190 -0.115 5.470 0.115 ;
        RECT  5.065 -0.115 5.190 0.235 ;
        RECT  4.810 -0.115 5.065 0.115 ;
        RECT  4.690 -0.115 4.810 0.145 ;
        RECT  3.995 -0.115 4.690 0.115 ;
        RECT  3.870 -0.115 3.995 0.245 ;
        RECT  3.100 -0.115 3.870 0.115 ;
        RECT  2.980 -0.115 3.100 0.195 ;
        RECT  1.520 -0.115 2.980 0.115 ;
        RECT  1.400 -0.115 1.520 0.125 ;
        RECT  1.190 -0.115 1.400 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.315 -0.115 1.070 0.115 ;
        RECT  0.245 -0.115 0.315 0.330 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 1.145 5.600 1.375 ;
        RECT  5.475 0.700 5.550 1.375 ;
        RECT  5.190 1.145 5.475 1.375 ;
        RECT  5.065 0.905 5.190 1.375 ;
        RECT  4.810 1.145 5.065 1.375 ;
        RECT  4.690 1.025 4.810 1.375 ;
        RECT  4.425 1.145 4.690 1.375 ;
        RECT  4.305 1.040 4.425 1.375 ;
        RECT  4.050 1.145 4.305 1.375 ;
        RECT  3.930 1.025 4.050 1.375 ;
        RECT  3.100 1.145 3.930 1.375 ;
        RECT  2.980 1.070 3.100 1.375 ;
        RECT  2.490 1.145 2.980 1.375 ;
        RECT  2.365 1.070 2.490 1.375 ;
        RECT  1.540 1.145 2.365 1.375 ;
        RECT  1.420 1.135 1.540 1.375 ;
        RECT  1.170 1.145 1.420 1.375 ;
        RECT  1.050 1.135 1.170 1.375 ;
        RECT  0.340 1.145 1.050 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.195 5.380 0.475 ;
        RECT  5.285 0.710 5.380 1.010 ;
        RECT  4.910 0.195 4.935 0.475 ;
        RECT  4.910 0.710 4.935 1.010 ;
        RECT  4.820 0.545 4.925 0.620 ;
        RECT  4.750 0.340 4.820 0.920 ;
        RECT  3.855 0.340 4.750 0.410 ;
        RECT  4.120 0.850 4.750 0.920 ;
        RECT  4.115 0.195 4.620 0.265 ;
        RECT  4.040 0.530 4.380 0.610 ;
        RECT  3.970 0.530 4.040 0.910 ;
        RECT  3.460 0.840 3.970 0.910 ;
        RECT  3.785 0.340 3.855 0.595 ;
        RECT  3.620 0.685 3.755 0.765 ;
        RECT  3.550 0.195 3.620 0.765 ;
        RECT  3.260 0.195 3.550 0.265 ;
        RECT  3.390 0.345 3.460 1.000 ;
        RECT  2.090 0.930 3.390 1.000 ;
        RECT  3.190 0.195 3.260 0.335 ;
        RECT  3.155 0.405 3.230 0.860 ;
        RECT  2.900 0.265 3.190 0.335 ;
        RECT  2.750 0.405 3.155 0.475 ;
        RECT  2.775 0.780 3.155 0.860 ;
        RECT  2.595 0.610 3.055 0.690 ;
        RECT  2.830 0.195 2.900 0.335 ;
        RECT  2.095 0.195 2.830 0.265 ;
        RECT  2.680 0.335 2.750 0.475 ;
        RECT  2.280 0.780 2.695 0.850 ;
        RECT  2.420 0.335 2.680 0.405 ;
        RECT  2.515 0.495 2.595 0.690 ;
        RECT  2.350 0.335 2.420 0.625 ;
        RECT  2.210 0.345 2.280 0.850 ;
        RECT  2.065 0.345 2.135 0.780 ;
        RECT  2.020 0.850 2.090 1.000 ;
        RECT  1.995 0.345 2.065 0.425 ;
        RECT  2.010 0.710 2.065 0.780 ;
        RECT  1.070 0.850 2.020 0.920 ;
        RECT  1.855 0.530 1.990 0.640 ;
        RECT  0.650 0.195 1.950 0.265 ;
        RECT  1.810 0.995 1.940 1.075 ;
        RECT  1.785 0.345 1.855 0.770 ;
        RECT  0.640 0.995 1.810 1.065 ;
        RECT  1.645 0.345 1.785 0.465 ;
        RECT  1.640 0.700 1.785 0.770 ;
        RECT  1.550 0.545 1.660 0.615 ;
        RECT  1.480 0.335 1.550 0.780 ;
        RECT  1.220 0.335 1.480 0.405 ;
        RECT  1.200 0.710 1.480 0.780 ;
        RECT  0.940 0.700 1.070 0.920 ;
        RECT  0.765 0.490 0.850 0.920 ;
        RECT  0.140 0.850 0.765 0.920 ;
        RECT  0.625 0.345 0.695 0.780 ;
        RECT  0.415 0.345 0.625 0.415 ;
        RECT  0.430 0.710 0.625 0.780 ;
        RECT  0.105 0.850 0.140 1.070 ;
        RECT  0.105 0.210 0.125 0.330 ;
        RECT  0.035 0.210 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.520 0.525 2.590 0.595 ;
        RECT  2.065 0.525 2.135 0.595 ;
        LAYER M2 ;
        RECT  2.015 0.525 2.640 0.595 ;
    END
END EDFCNQD4BWP40

MACRO EDFQD0BWP40
    CLASS CORE ;
    FOREIGN EDFQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.021400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.285 0.775 ;
        RECT  0.175 0.470 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.635 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.155 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.270 ;
        RECT  2.595 -0.115 3.375 0.115 ;
        RECT  2.525 -0.115 2.595 0.260 ;
        RECT  2.010 -0.115 2.525 0.115 ;
        RECT  1.890 -0.115 2.010 0.125 ;
        RECT  1.120 -0.115 1.890 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.390 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.950 3.815 1.375 ;
        RECT  3.470 1.145 3.745 1.375 ;
        RECT  3.350 1.010 3.470 1.375 ;
        RECT  2.630 1.145 3.350 1.375 ;
        RECT  2.510 1.050 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 1.050 2.060 1.375 ;
        RECT  1.050 1.145 1.940 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.340 1.145 0.930 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.705 0.395 3.775 0.810 ;
        RECT  3.635 0.395 3.705 0.465 ;
        RECT  3.635 0.740 3.705 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 1.055 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.920 ;
        RECT  3.015 0.850 3.415 0.920 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.110 0.195 3.185 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.945 0.345 3.015 0.980 ;
        RECT  1.615 0.910 2.945 0.980 ;
        RECT  2.790 0.195 2.860 0.840 ;
        RECT  2.405 0.340 2.790 0.410 ;
        RECT  2.420 0.750 2.790 0.840 ;
        RECT  2.270 0.520 2.710 0.650 ;
        RECT  2.340 0.730 2.420 0.840 ;
        RECT  2.335 0.195 2.405 0.410 ;
        RECT  1.630 0.195 2.335 0.265 ;
        RECT  2.200 0.730 2.255 0.800 ;
        RECT  2.200 0.350 2.220 0.470 ;
        RECT  2.130 0.350 2.200 0.800 ;
        RECT  1.885 0.535 2.130 0.655 ;
        RECT  1.815 0.770 1.870 0.840 ;
        RECT  1.745 0.370 1.815 0.840 ;
        RECT  1.615 0.690 1.640 0.760 ;
        RECT  1.545 0.350 1.615 0.760 ;
        RECT  1.545 0.845 1.615 0.980 ;
        RECT  1.520 0.690 1.545 0.760 ;
        RECT  1.025 0.845 1.545 0.915 ;
        RECT  0.595 0.195 1.470 0.265 ;
        RECT  0.605 0.985 1.450 1.055 ;
        RECT  1.250 0.345 1.320 0.775 ;
        RECT  1.150 0.345 1.250 0.425 ;
        RECT  1.145 0.705 1.250 0.775 ;
        RECT  0.955 0.700 1.025 0.915 ;
        RECT  0.880 0.700 0.955 0.820 ;
        RECT  0.735 0.505 0.805 0.915 ;
        RECT  0.140 0.845 0.735 0.915 ;
        RECT  0.595 0.335 0.665 0.775 ;
        RECT  0.535 0.335 0.595 0.405 ;
        RECT  0.365 0.705 0.595 0.775 ;
        RECT  0.415 0.305 0.535 0.405 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.315 0.525 2.385 0.595 ;
        RECT  1.545 0.525 1.615 0.595 ;
        LAYER M2 ;
        RECT  1.495 0.525 2.435 0.595 ;
    END
END EDFQD0BWP40

MACRO EDFQD1BWP40
    CLASS CORE ;
    FOREIGN EDFQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.285 0.775 ;
        RECT  0.175 0.470 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.635 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.150 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.595 -0.115 3.375 0.115 ;
        RECT  2.525 -0.115 2.595 0.260 ;
        RECT  2.010 -0.115 2.525 0.115 ;
        RECT  1.890 -0.115 2.010 0.125 ;
        RECT  1.120 -0.115 1.890 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.390 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.470 1.145 3.745 1.375 ;
        RECT  3.350 1.010 3.470 1.375 ;
        RECT  2.630 1.145 3.350 1.375 ;
        RECT  2.510 1.050 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 1.050 2.060 1.375 ;
        RECT  1.050 1.145 1.940 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.340 1.145 0.930 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.705 0.395 3.775 0.810 ;
        RECT  3.635 0.395 3.705 0.465 ;
        RECT  3.635 0.740 3.705 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 1.065 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.920 ;
        RECT  3.015 0.850 3.415 0.920 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.110 0.195 3.185 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.945 0.350 3.015 0.980 ;
        RECT  1.615 0.910 2.945 0.980 ;
        RECT  2.790 0.195 2.860 0.840 ;
        RECT  2.440 0.340 2.790 0.410 ;
        RECT  2.420 0.750 2.790 0.840 ;
        RECT  2.270 0.520 2.710 0.650 ;
        RECT  2.370 0.195 2.440 0.410 ;
        RECT  2.340 0.730 2.420 0.840 ;
        RECT  1.630 0.195 2.370 0.265 ;
        RECT  2.200 0.730 2.255 0.800 ;
        RECT  2.200 0.350 2.220 0.470 ;
        RECT  2.130 0.350 2.200 0.800 ;
        RECT  1.885 0.535 2.130 0.655 ;
        RECT  1.815 0.770 1.870 0.840 ;
        RECT  1.745 0.370 1.815 0.840 ;
        RECT  1.615 0.690 1.640 0.760 ;
        RECT  1.545 0.350 1.615 0.760 ;
        RECT  1.545 0.845 1.615 0.980 ;
        RECT  1.520 0.690 1.545 0.760 ;
        RECT  1.025 0.845 1.545 0.915 ;
        RECT  0.595 0.195 1.470 0.265 ;
        RECT  0.605 0.985 1.450 1.055 ;
        RECT  1.250 0.345 1.320 0.775 ;
        RECT  1.150 0.345 1.250 0.425 ;
        RECT  1.145 0.705 1.250 0.775 ;
        RECT  0.955 0.700 1.025 0.915 ;
        RECT  0.880 0.700 0.955 0.820 ;
        RECT  0.735 0.505 0.805 0.915 ;
        RECT  0.140 0.845 0.735 0.915 ;
        RECT  0.595 0.335 0.665 0.775 ;
        RECT  0.535 0.335 0.595 0.405 ;
        RECT  0.365 0.705 0.595 0.775 ;
        RECT  0.415 0.305 0.535 0.405 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.315 0.525 2.385 0.595 ;
        RECT  1.545 0.525 1.615 0.595 ;
        LAYER M2 ;
        RECT  1.495 0.525 2.435 0.595 ;
    END
END EDFQD1BWP40

MACRO EDFQD2BWP40
    CLASS CORE ;
    FOREIGN EDFQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.285 0.775 ;
        RECT  0.175 0.470 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.635 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.150 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.260 -0.115 4.340 0.115 ;
        RECT  4.185 -0.115 4.260 0.450 ;
        RECT  3.815 -0.115 4.185 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.595 -0.115 3.375 0.115 ;
        RECT  2.525 -0.115 2.595 0.260 ;
        RECT  2.010 -0.115 2.525 0.115 ;
        RECT  1.890 -0.115 2.010 0.125 ;
        RECT  1.120 -0.115 1.890 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.390 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 1.145 4.340 1.375 ;
        RECT  4.195 0.675 4.270 1.375 ;
        RECT  3.815 1.145 4.195 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.470 1.145 3.745 1.375 ;
        RECT  3.350 1.010 3.470 1.375 ;
        RECT  2.630 1.145 3.350 1.375 ;
        RECT  2.510 1.050 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 1.050 2.060 1.375 ;
        RECT  1.050 1.145 1.940 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.340 1.145 0.930 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.705 0.395 3.775 0.810 ;
        RECT  3.635 0.395 3.705 0.465 ;
        RECT  3.635 0.740 3.705 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 1.045 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.920 ;
        RECT  3.015 0.850 3.415 0.920 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.110 0.195 3.185 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.945 0.350 3.015 0.980 ;
        RECT  1.615 0.910 2.945 0.980 ;
        RECT  2.790 0.195 2.860 0.840 ;
        RECT  2.440 0.340 2.790 0.410 ;
        RECT  2.420 0.750 2.790 0.840 ;
        RECT  2.270 0.520 2.710 0.650 ;
        RECT  2.370 0.195 2.440 0.410 ;
        RECT  2.340 0.730 2.420 0.840 ;
        RECT  1.630 0.195 2.370 0.265 ;
        RECT  2.200 0.730 2.255 0.800 ;
        RECT  2.200 0.350 2.220 0.470 ;
        RECT  2.130 0.350 2.200 0.800 ;
        RECT  1.885 0.535 2.130 0.655 ;
        RECT  1.815 0.770 1.870 0.840 ;
        RECT  1.745 0.370 1.815 0.840 ;
        RECT  1.615 0.690 1.640 0.760 ;
        RECT  1.545 0.350 1.615 0.760 ;
        RECT  1.545 0.845 1.615 0.980 ;
        RECT  1.520 0.690 1.545 0.760 ;
        RECT  1.025 0.845 1.545 0.915 ;
        RECT  0.595 0.195 1.470 0.265 ;
        RECT  0.605 0.985 1.450 1.055 ;
        RECT  1.250 0.345 1.320 0.775 ;
        RECT  1.150 0.345 1.250 0.425 ;
        RECT  1.145 0.705 1.250 0.775 ;
        RECT  0.955 0.700 1.025 0.915 ;
        RECT  0.880 0.700 0.955 0.820 ;
        RECT  0.735 0.505 0.805 0.915 ;
        RECT  0.140 0.845 0.735 0.915 ;
        RECT  0.595 0.335 0.665 0.775 ;
        RECT  0.535 0.335 0.595 0.405 ;
        RECT  0.365 0.705 0.595 0.775 ;
        RECT  0.415 0.305 0.535 0.405 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.315 0.525 2.385 0.595 ;
        RECT  1.545 0.525 1.615 0.595 ;
        LAYER M2 ;
        RECT  1.495 0.525 2.435 0.595 ;
    END
END EDFQD2BWP40

MACRO EDFQD4BWP40
    CLASS CORE ;
    FOREIGN EDFQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.195 4.400 0.475 ;
        RECT  4.305 0.710 4.400 1.020 ;
        RECT  4.235 0.355 4.305 0.475 ;
        RECT  4.235 0.710 4.305 0.830 ;
        RECT  4.025 0.355 4.235 0.830 ;
        RECT  4.000 0.355 4.025 0.475 ;
        RECT  4.000 0.710 4.025 0.830 ;
        RECT  3.930 0.195 4.000 0.475 ;
        RECT  3.930 0.710 4.000 1.020 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.700 0.285 0.775 ;
        RECT  0.175 0.470 0.245 0.775 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.525 0.635 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.150 0.625 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 -0.115 4.620 0.115 ;
        RECT  4.490 -0.115 4.570 0.430 ;
        RECT  4.190 -0.115 4.490 0.115 ;
        RECT  4.115 -0.115 4.190 0.270 ;
        RECT  3.805 -0.115 4.115 0.115 ;
        RECT  3.735 -0.115 3.805 0.315 ;
        RECT  3.425 -0.115 3.735 0.115 ;
        RECT  3.355 -0.115 3.425 0.315 ;
        RECT  2.585 -0.115 3.355 0.115 ;
        RECT  2.515 -0.115 2.585 0.260 ;
        RECT  2.010 -0.115 2.515 0.115 ;
        RECT  1.890 -0.115 2.010 0.125 ;
        RECT  1.120 -0.115 1.890 0.115 ;
        RECT  1.000 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.390 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.145 4.620 1.375 ;
        RECT  4.480 0.705 4.570 1.375 ;
        RECT  4.205 1.145 4.480 1.375 ;
        RECT  4.095 0.905 4.205 1.375 ;
        RECT  3.825 1.145 4.095 1.375 ;
        RECT  3.715 0.905 3.825 1.375 ;
        RECT  3.460 1.145 3.715 1.375 ;
        RECT  3.330 1.010 3.460 1.375 ;
        RECT  2.610 1.145 3.330 1.375 ;
        RECT  2.490 1.050 2.610 1.375 ;
        RECT  2.080 1.145 2.490 1.375 ;
        RECT  1.960 1.050 2.080 1.375 ;
        RECT  1.050 1.145 1.960 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.340 1.145 0.930 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.195 4.400 0.475 ;
        RECT  4.305 0.710 4.400 1.020 ;
        RECT  3.930 0.195 3.955 0.475 ;
        RECT  3.930 0.710 3.955 1.020 ;
        RECT  3.825 0.545 3.945 0.615 ;
        RECT  3.755 0.395 3.825 0.810 ;
        RECT  3.615 0.395 3.755 0.465 ;
        RECT  3.615 0.740 3.755 0.810 ;
        RECT  3.465 0.545 3.625 0.615 ;
        RECT  3.545 0.185 3.615 0.465 ;
        RECT  3.545 0.740 3.615 0.965 ;
        RECT  3.325 0.395 3.545 0.465 ;
        RECT  3.395 0.545 3.465 0.920 ;
        RECT  3.015 0.850 3.395 0.920 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.090 0.195 3.165 0.780 ;
        RECT  2.840 0.195 3.090 0.265 ;
        RECT  2.995 0.850 3.015 0.980 ;
        RECT  2.925 0.350 2.995 0.980 ;
        RECT  1.615 0.910 2.925 0.980 ;
        RECT  2.770 0.195 2.840 0.840 ;
        RECT  2.430 0.340 2.770 0.410 ;
        RECT  2.400 0.750 2.770 0.840 ;
        RECT  2.260 0.520 2.690 0.650 ;
        RECT  2.360 0.195 2.430 0.410 ;
        RECT  2.320 0.730 2.400 0.840 ;
        RECT  1.630 0.195 2.360 0.265 ;
        RECT  2.190 0.730 2.235 0.800 ;
        RECT  2.190 0.350 2.210 0.470 ;
        RECT  2.120 0.350 2.190 0.800 ;
        RECT  1.885 0.535 2.120 0.655 ;
        RECT  1.815 0.770 1.870 0.840 ;
        RECT  1.745 0.370 1.815 0.840 ;
        RECT  1.615 0.690 1.640 0.760 ;
        RECT  1.545 0.350 1.615 0.760 ;
        RECT  1.545 0.845 1.615 0.980 ;
        RECT  1.520 0.690 1.545 0.760 ;
        RECT  1.025 0.845 1.545 0.915 ;
        RECT  0.595 0.195 1.470 0.265 ;
        RECT  0.605 0.985 1.450 1.055 ;
        RECT  1.250 0.345 1.320 0.775 ;
        RECT  1.150 0.345 1.250 0.425 ;
        RECT  1.145 0.705 1.250 0.775 ;
        RECT  0.955 0.700 1.025 0.915 ;
        RECT  0.880 0.700 0.955 0.820 ;
        RECT  0.735 0.505 0.805 0.915 ;
        RECT  0.140 0.845 0.735 0.915 ;
        RECT  0.595 0.335 0.665 0.775 ;
        RECT  0.535 0.335 0.595 0.405 ;
        RECT  0.365 0.705 0.595 0.775 ;
        RECT  0.415 0.305 0.535 0.405 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.305 0.525 2.375 0.595 ;
        RECT  1.545 0.525 1.615 0.595 ;
        LAYER M2 ;
        RECT  1.495 0.525 2.425 0.595 ;
    END
END EDFQD4BWP40

MACRO FA1D0BWP40
    CLASS CORE ;
    FOREIGN FA1D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.058000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.185 3.325 1.055 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.066650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.785 ;
        RECT  2.780 0.355 2.835 0.435 ;
        RECT  2.780 0.715 2.835 0.785 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.495 1.505 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.280 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.075 -0.115 3.360 0.115 ;
        RECT  2.965 -0.115 3.075 0.125 ;
        RECT  2.530 -0.115 2.965 0.115 ;
        RECT  2.410 -0.115 2.530 0.125 ;
        RECT  1.550 -0.115 2.410 0.115 ;
        RECT  1.430 -0.115 1.550 0.275 ;
        RECT  0.590 -0.115 1.430 0.115 ;
        RECT  0.470 -0.115 0.590 0.240 ;
        RECT  0.155 -0.115 0.470 0.115 ;
        RECT  0.035 -0.115 0.155 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.095 1.145 3.360 1.375 ;
        RECT  2.975 1.025 3.095 1.375 ;
        RECT  2.510 1.145 2.975 1.375 ;
        RECT  2.390 1.025 2.510 1.375 ;
        RECT  1.550 1.145 2.390 1.375 ;
        RECT  1.430 1.025 1.550 1.375 ;
        RECT  0.590 1.145 1.430 1.375 ;
        RECT  0.470 1.025 0.590 1.375 ;
        RECT  0.155 1.145 0.470 1.375 ;
        RECT  0.035 0.815 0.155 1.375 ;
        RECT  0.000 1.145 0.035 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.085 0.205 3.155 0.955 ;
        RECT  1.990 0.205 3.085 0.275 ;
        RECT  1.990 0.885 3.085 0.955 ;
        RECT  2.665 0.525 2.765 0.635 ;
        RECT  1.240 0.355 2.710 0.425 ;
        RECT  1.885 0.735 2.710 0.805 ;
        RECT  1.675 0.545 2.665 0.615 ;
        RECT  1.815 0.735 1.885 0.940 ;
        RECT  1.240 0.870 1.815 0.940 ;
        RECT  1.605 0.545 1.675 0.790 ;
        RECT  0.925 0.720 1.605 0.790 ;
        RECT  0.740 0.205 1.180 0.275 ;
        RECT  0.260 0.870 1.170 0.940 ;
        RECT  0.925 0.355 0.980 0.425 ;
        RECT  0.855 0.355 0.925 0.790 ;
        RECT  0.670 0.205 0.740 0.390 ;
        RECT  0.260 0.320 0.670 0.390 ;
    END
END FA1D0BWP40

MACRO FA1D1BWP40
    CLASS CORE ;
    FOREIGN FA1D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.113100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.235 0.185 3.325 1.045 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.082500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.785 ;
        RECT  2.780 0.355 2.835 0.435 ;
        RECT  2.780 0.715 2.835 0.785 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.057600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.495 1.505 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.089600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.445 0.495 0.595 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.089600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.255 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.075 -0.115 3.360 0.115 ;
        RECT  2.965 -0.115 3.075 0.125 ;
        RECT  2.530 -0.115 2.965 0.115 ;
        RECT  2.410 -0.115 2.530 0.125 ;
        RECT  1.550 -0.115 2.410 0.115 ;
        RECT  1.430 -0.115 1.550 0.235 ;
        RECT  0.590 -0.115 1.430 0.115 ;
        RECT  0.470 -0.115 0.590 0.255 ;
        RECT  0.155 -0.115 0.470 0.115 ;
        RECT  0.035 -0.115 0.155 0.255 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.095 1.145 3.360 1.375 ;
        RECT  2.975 1.005 3.095 1.375 ;
        RECT  2.510 1.145 2.975 1.375 ;
        RECT  2.390 1.025 2.510 1.375 ;
        RECT  1.550 1.145 2.390 1.375 ;
        RECT  1.430 1.025 1.550 1.375 ;
        RECT  0.590 1.145 1.430 1.375 ;
        RECT  0.470 1.015 0.590 1.375 ;
        RECT  0.130 1.145 0.470 1.375 ;
        RECT  0.060 0.725 0.130 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.085 0.205 3.155 0.935 ;
        RECT  1.990 0.205 3.085 0.275 ;
        RECT  1.990 0.865 3.085 0.935 ;
        RECT  2.665 0.525 2.765 0.635 ;
        RECT  1.240 0.355 2.710 0.425 ;
        RECT  1.885 0.715 2.710 0.785 ;
        RECT  1.675 0.545 2.665 0.615 ;
        RECT  1.815 0.715 1.885 0.935 ;
        RECT  1.240 0.865 1.815 0.935 ;
        RECT  1.605 0.545 1.675 0.785 ;
        RECT  0.925 0.715 1.605 0.785 ;
        RECT  0.740 0.205 1.180 0.275 ;
        RECT  0.265 0.865 1.170 0.935 ;
        RECT  0.925 0.355 0.980 0.425 ;
        RECT  0.855 0.355 0.925 0.785 ;
        RECT  0.670 0.205 0.740 0.405 ;
        RECT  0.260 0.335 0.670 0.405 ;
    END
END FA1D1BWP40

MACRO FA1D2BWP40
    CLASS CORE ;
    FOREIGN FA1D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 0.405 3.465 0.790 ;
        RECT  3.405 0.405 3.410 1.045 ;
        RECT  3.375 0.185 3.405 1.045 ;
        RECT  3.330 0.185 3.375 0.475 ;
        RECT  3.330 0.705 3.375 1.045 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.099000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.355 3.075 0.805 ;
        RECT  2.930 0.355 2.975 0.485 ;
        RECT  2.930 0.705 2.975 0.805 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.057600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.485 0.640 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.089600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.089600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.255 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 -0.115 3.640 0.115 ;
        RECT  3.515 -0.115 3.585 0.340 ;
        RECT  3.205 -0.115 3.515 0.115 ;
        RECT  3.090 -0.115 3.205 0.125 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.125 ;
        RECT  2.490 -0.115 2.690 0.115 ;
        RECT  2.370 -0.115 2.490 0.125 ;
        RECT  1.530 -0.115 2.370 0.115 ;
        RECT  1.410 -0.115 1.530 0.275 ;
        RECT  0.590 -0.115 1.410 0.115 ;
        RECT  0.470 -0.115 0.590 0.255 ;
        RECT  0.155 -0.115 0.470 0.115 ;
        RECT  0.035 -0.115 0.155 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 1.145 3.640 1.375 ;
        RECT  3.515 0.860 3.585 1.375 ;
        RECT  3.230 1.145 3.515 1.375 ;
        RECT  3.110 1.045 3.230 1.375 ;
        RECT  2.855 1.145 3.110 1.375 ;
        RECT  2.730 1.020 2.855 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 1.025 2.470 1.375 ;
        RECT  1.530 1.145 2.350 1.375 ;
        RECT  1.410 1.005 1.530 1.375 ;
        RECT  0.590 1.145 1.410 1.375 ;
        RECT  0.470 1.005 0.590 1.375 ;
        RECT  0.130 1.145 0.470 1.375 ;
        RECT  0.060 0.725 0.130 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.260 0.520 3.270 0.645 ;
        RECT  3.250 0.520 3.260 0.950 ;
        RECT  3.180 0.205 3.250 0.950 ;
        RECT  1.960 0.205 3.180 0.275 ;
        RECT  1.955 0.880 3.180 0.950 ;
        RECT  1.635 0.545 2.835 0.615 ;
        RECT  1.220 0.355 2.670 0.425 ;
        RECT  1.865 0.730 2.670 0.800 ;
        RECT  1.795 0.730 1.865 0.935 ;
        RECT  1.220 0.865 1.795 0.935 ;
        RECT  1.565 0.545 1.635 0.785 ;
        RECT  0.905 0.715 1.565 0.785 ;
        RECT  0.740 0.205 1.160 0.275 ;
        RECT  0.265 0.865 1.150 0.935 ;
        RECT  0.905 0.355 0.960 0.425 ;
        RECT  0.835 0.355 0.905 0.785 ;
        RECT  0.670 0.205 0.740 0.405 ;
        RECT  0.260 0.335 0.670 0.405 ;
    END
END FA1D2BWP40

MACRO FA1D4BWP40
    CLASS CORE ;
    FOREIGN FA1D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.245700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.660 0.185 6.735 0.465 ;
        RECT  6.655 0.730 6.735 1.035 ;
        RECT  6.615 0.355 6.660 0.465 ;
        RECT  6.615 0.730 6.655 0.815 ;
        RECT  6.405 0.355 6.615 0.815 ;
        RECT  6.345 0.355 6.405 0.465 ;
        RECT  6.350 0.730 6.405 0.815 ;
        RECT  6.270 0.730 6.350 1.035 ;
        RECT  6.270 0.185 6.345 0.465 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.198000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.355 5.985 0.445 ;
        RECT  5.915 0.715 5.985 0.805 ;
        RECT  5.705 0.355 5.915 0.805 ;
        RECT  5.470 0.355 5.705 0.485 ;
        RECT  5.470 0.705 5.705 0.805 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.093800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.060 0.485 3.995 0.555 ;
        RECT  2.910 0.355 3.060 0.555 ;
        RECT  2.835 0.355 2.910 0.625 ;
        RECT  1.810 0.540 2.835 0.625 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.151400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.144400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.280 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.945 -0.115 7.000 0.115 ;
        RECT  6.875 -0.115 6.945 0.445 ;
        RECT  6.535 -0.115 6.875 0.115 ;
        RECT  6.465 -0.115 6.535 0.265 ;
        RECT  6.145 -0.115 6.465 0.115 ;
        RECT  6.075 -0.115 6.145 0.460 ;
        RECT  5.755 -0.115 6.075 0.115 ;
        RECT  5.685 -0.115 5.755 0.275 ;
        RECT  5.365 -0.115 5.685 0.115 ;
        RECT  5.280 -0.115 5.365 0.445 ;
        RECT  4.965 -0.115 5.280 0.115 ;
        RECT  4.890 -0.115 4.965 0.265 ;
        RECT  4.580 -0.115 4.890 0.115 ;
        RECT  4.460 -0.115 4.580 0.265 ;
        RECT  4.150 -0.115 4.460 0.115 ;
        RECT  4.030 -0.115 4.150 0.265 ;
        RECT  2.450 -0.115 4.030 0.115 ;
        RECT  2.330 -0.115 2.450 0.300 ;
        RECT  1.510 -0.115 2.330 0.115 ;
        RECT  1.390 -0.115 1.510 0.210 ;
        RECT  0.590 -0.115 1.390 0.115 ;
        RECT  0.470 -0.115 0.590 0.255 ;
        RECT  0.155 -0.115 0.470 0.115 ;
        RECT  0.035 -0.115 0.155 0.275 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.945 1.145 7.000 1.375 ;
        RECT  6.875 0.720 6.945 1.375 ;
        RECT  6.560 1.145 6.875 1.375 ;
        RECT  6.440 0.910 6.560 1.375 ;
        RECT  6.170 1.145 6.440 1.375 ;
        RECT  6.040 1.045 6.170 1.375 ;
        RECT  5.785 1.145 6.040 1.375 ;
        RECT  5.660 1.045 5.785 1.375 ;
        RECT  5.400 1.145 5.660 1.375 ;
        RECT  5.280 1.045 5.400 1.375 ;
        RECT  4.990 1.145 5.280 1.375 ;
        RECT  4.850 1.045 4.990 1.375 ;
        RECT  4.560 1.145 4.850 1.375 ;
        RECT  4.435 1.045 4.560 1.375 ;
        RECT  4.135 1.145 4.435 1.375 ;
        RECT  4.015 1.045 4.135 1.375 ;
        RECT  2.465 1.145 4.015 1.375 ;
        RECT  2.345 1.045 2.465 1.375 ;
        RECT  1.525 1.145 2.345 1.375 ;
        RECT  1.405 1.005 1.525 1.375 ;
        RECT  0.590 1.145 1.405 1.375 ;
        RECT  0.470 1.005 0.590 1.375 ;
        RECT  0.130 1.145 0.470 1.375 ;
        RECT  0.060 0.705 0.130 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.685 0.185 6.735 0.465 ;
        RECT  6.685 0.730 6.735 1.035 ;
        RECT  6.270 0.185 6.335 0.465 ;
        RECT  6.270 0.730 6.335 1.035 ;
        RECT  5.470 0.355 5.635 0.485 ;
        RECT  5.470 0.705 5.635 0.805 ;
        RECT  6.200 0.550 6.310 0.650 ;
        RECT  6.120 0.550 6.200 0.975 ;
        RECT  2.165 0.905 6.120 0.975 ;
        RECT  4.485 0.555 5.625 0.625 ;
        RECT  3.175 0.345 5.190 0.415 ;
        RECT  2.090 0.905 2.165 1.070 ;
        RECT  2.010 0.195 2.130 0.455 ;
        RECT  2.015 0.980 2.090 1.070 ;
        RECT  0.255 0.855 1.965 0.925 ;
        RECT  1.855 0.280 1.935 0.440 ;
        RECT  0.815 0.280 1.855 0.350 ;
        RECT  1.255 0.420 1.745 0.490 ;
        RECT  1.165 0.420 1.255 0.785 ;
        RECT  0.925 0.420 1.165 0.495 ;
        RECT  0.910 0.715 1.165 0.785 ;
        RECT  0.735 0.280 0.815 0.405 ;
        RECT  0.260 0.335 0.735 0.405 ;
        RECT  4.685 0.735 5.190 0.805 ;
        RECT  4.615 0.735 4.685 0.835 ;
        RECT  3.180 0.765 4.615 0.835 ;
        RECT  4.415 0.555 4.485 0.695 ;
        RECT  3.085 0.625 4.415 0.695 ;
        RECT  2.710 0.205 3.555 0.275 ;
        RECT  3.010 0.625 3.085 0.785 ;
        RECT  1.255 0.715 3.010 0.785 ;
        RECT  2.630 0.205 2.710 0.455 ;
        RECT  2.130 0.380 2.630 0.455 ;
    END
END FA1D4BWP40

MACRO FILL16BWP40
    CLASS CORE ;
    FOREIGN FILL16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.240 1.375 ;
        END
    END VDD
END FILL16BWP40

MACRO FILL2BWP40
    CLASS CORE ;
    FOREIGN FILL2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.280 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.280 1.375 ;
        END
    END VDD
END FILL2BWP40

MACRO FILL32BWP40
    CLASS CORE ;
    FOREIGN FILL32BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.480 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 4.480 1.375 ;
        END
    END VDD
END FILL32BWP40

MACRO FILL3BWP40
    CLASS CORE ;
    FOREIGN FILL3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
END FILL3BWP40

MACRO FILL4BWP40
    CLASS CORE ;
    FOREIGN FILL4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.560 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.560 1.375 ;
        END
    END VDD
END FILL4BWP40

MACRO FILL64BWP40
    CLASS CORE ;
    FOREIGN FILL64BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 8.960 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 8.960 1.375 ;
        END
    END VDD
END FILL64BWP40

MACRO FILL8BWP40
    CLASS CORE ;
    FOREIGN FILL8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.120 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 1.120 1.375 ;
        END
    END VDD
END FILL8BWP40

MACRO GAN2D1BWP40
    CLASS CORE ;
    FOREIGN GAN2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.200 1.365 1.060 ;
        RECT  1.170 0.200 1.295 0.280 ;
        RECT  1.190 0.980 1.295 1.060 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.320 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.320 ;
        RECT  0.210 -0.115 0.810 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.890 1.145 0.990 1.375 ;
        RECT  0.810 0.940 0.890 1.375 ;
        RECT  0.610 1.145 0.810 1.375 ;
        RECT  0.490 0.985 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.500 1.225 0.785 ;
        RECT  0.945 0.715 1.155 0.785 ;
        RECT  0.875 0.500 0.945 0.785 ;
        RECT  0.665 0.715 0.875 0.785 ;
        RECT  0.595 0.200 0.665 0.915 ;
        RECT  0.490 0.200 0.595 0.280 ;
        RECT  0.270 0.845 0.595 0.915 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAN2D1BWP40

MACRO GAN2D2BWP40
    CLASS CORE ;
    FOREIGN GAN2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.365 0.920 ;
        RECT  1.100 0.345 1.295 0.415 ;
        RECT  0.980 0.850 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.415 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.210 -0.115 0.790 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.915 1.145 1.190 1.375 ;
        RECT  0.795 0.980 0.915 1.375 ;
        RECT  0.610 1.145 0.795 1.375 ;
        RECT  0.490 0.985 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.520 1.225 0.640 ;
        RECT  0.595 0.200 0.665 0.915 ;
        RECT  0.490 0.200 0.595 0.280 ;
        RECT  0.270 0.845 0.595 0.915 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAN2D2BWP40

MACRO GAOI21D1BWP40
    CLASS CORE ;
    FOREIGN GAOI21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.260250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.190 1.300 0.290 ;
        RECT  1.190 0.190 1.260 0.415 ;
        RECT  0.920 0.345 1.190 0.415 ;
        RECT  0.850 0.205 0.920 0.415 ;
        RECT  0.665 0.205 0.850 0.275 ;
        RECT  0.595 0.205 0.665 0.915 ;
        RECT  0.490 0.205 0.595 0.275 ;
        RECT  0.290 0.845 0.595 0.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 1.250 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.260 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        RECT  0.355 0.495 0.435 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 1.400 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.210 -0.115 0.990 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  0.990 0.850 1.110 1.375 ;
        RECT  0.000 1.145 0.990 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.970 1.310 1.070 ;
        RECT  1.190 0.710 1.260 1.070 ;
        RECT  0.920 0.710 1.190 0.780 ;
        RECT  0.850 0.710 0.920 1.055 ;
        RECT  0.070 0.985 0.850 1.055 ;
        RECT  0.300 0.185 0.400 0.405 ;
    END
END GAOI21D1BWP40

MACRO GAOI21D2BWP40
    CLASS CORE ;
    FOREIGN GAOI21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.398000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.200 2.065 0.915 ;
        RECT  1.890 0.200 1.995 0.280 ;
        RECT  1.505 0.825 1.995 0.915 ;
        RECT  1.505 0.195 1.610 0.290 ;
        RECT  1.435 0.195 1.505 0.915 ;
        RECT  1.285 0.195 1.435 0.270 ;
        RECT  1.190 0.195 1.285 0.415 ;
        RECT  0.885 0.345 1.190 0.415 ;
        RECT  0.815 0.185 0.885 0.415 ;
        RECT  0.665 0.345 0.815 0.415 ;
        RECT  0.595 0.345 0.665 0.915 ;
        RECT  0.385 0.825 0.595 0.915 ;
        RECT  0.290 0.775 0.385 0.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.495 1.250 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.925 0.670 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 2.100 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.610 -0.115 0.990 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 2.100 1.375 ;
        RECT  0.990 0.850 1.110 1.375 ;
        RECT  0.000 1.145 0.990 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.985 2.010 1.055 ;
        RECT  1.700 0.185 1.800 0.415 ;
        RECT  1.190 0.710 1.260 1.055 ;
        RECT  0.920 0.710 1.190 0.780 ;
        RECT  0.850 0.710 0.920 1.055 ;
        RECT  0.070 0.985 0.850 1.055 ;
        RECT  0.300 0.185 0.400 0.405 ;
        LAYER VIA1 ;
        RECT  1.715 0.300 1.785 0.370 ;
        RECT  0.315 0.300 0.385 0.370 ;
        LAYER M2 ;
        RECT  0.265 0.300 1.835 0.370 ;
    END
END GAOI21D2BWP40

MACRO GAOI22D1BWP40
    CLASS CORE ;
    FOREIGN GAOI22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.990 1.365 1.060 ;
        RECT  0.805 0.200 0.910 0.275 ;
        RECT  0.735 0.200 0.805 1.060 ;
        RECT  0.490 0.200 0.735 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.315 0.495 0.595 0.650 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.295 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.445 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.210 -0.115 1.190 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.145 1.400 1.375 ;
        RECT  0.490 0.985 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.845 1.200 0.920 ;
        RECT  1.085 0.185 1.100 0.290 ;
        RECT  1.015 0.185 1.085 0.465 ;
        RECT  1.015 0.755 1.085 0.920 ;
        RECT  1.000 0.185 1.015 0.290 ;
        RECT  0.905 0.845 1.015 0.920 ;
        RECT  0.300 0.185 0.400 0.405 ;
        RECT  0.315 0.745 0.385 1.065 ;
        LAYER VIA1 ;
        RECT  1.015 0.805 1.085 0.875 ;
        RECT  0.315 0.805 0.385 0.875 ;
        LAYER M2 ;
        RECT  0.265 0.805 1.135 0.875 ;
    END
END GAOI22D1BWP40

MACRO GAOI22D2BWP40
    CLASS CORE ;
    FOREIGN GAOI22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.272000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.815 2.625 0.920 ;
        RECT  2.130 0.345 2.135 0.920 ;
        RECT  2.065 0.345 2.130 0.910 ;
        RECT  1.800 0.345 2.065 0.415 ;
        RECT  1.810 0.705 2.065 0.910 ;
        RECT  1.685 0.705 1.810 0.915 ;
        RECT  1.700 0.185 1.800 0.415 ;
        RECT  0.735 0.705 1.685 0.775 ;
        RECT  1.000 0.185 1.100 0.415 ;
        RECT  0.735 0.345 1.000 0.415 ;
        RECT  0.665 0.345 0.735 0.775 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.560 0.650 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.495 1.270 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.495 2.675 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.495 1.955 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.275 ;
        RECT  0.410 -0.115 2.390 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 2.800 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.985 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.555 0.990 2.710 1.060 ;
        RECT  2.600 0.185 2.700 0.425 ;
        RECT  2.310 0.355 2.600 0.425 ;
        RECT  2.240 0.205 2.310 0.425 ;
        RECT  1.890 0.205 2.240 0.275 ;
        RECT  1.500 0.190 1.600 0.410 ;
        RECT  1.475 0.845 1.555 1.060 ;
        RECT  0.280 0.845 1.475 0.915 ;
        RECT  1.200 0.190 1.300 0.410 ;
        RECT  0.560 0.205 0.910 0.275 ;
        RECT  0.490 0.205 0.560 0.425 ;
        RECT  0.200 0.355 0.490 0.425 ;
        RECT  0.100 0.185 0.200 0.425 ;
        LAYER VIA1 ;
        RECT  2.240 0.245 2.310 0.315 ;
        RECT  1.515 0.245 1.585 0.315 ;
        RECT  1.215 0.245 1.285 0.315 ;
        RECT  0.490 0.245 0.560 0.315 ;
        LAYER M2 ;
        RECT  1.465 0.245 2.360 0.315 ;
        RECT  0.440 0.245 1.335 0.315 ;
    END
END GAOI22D2BWP40

MACRO GBUFFD1BWP40
    CLASS CORE ;
    FOREIGN GBUFFD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.200 0.665 1.060 ;
        RECT  0.490 0.200 0.595 0.280 ;
        RECT  0.490 0.980 0.595 1.060 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.265 0.495 0.385 0.640 ;
        RECT  0.175 0.355 0.265 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.400 -0.115 0.700 0.115 ;
        RECT  0.300 -0.115 0.400 0.290 ;
        RECT  0.000 -0.115 0.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.145 0.700 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.455 0.500 0.525 0.780 ;
        RECT  0.105 0.710 0.455 0.780 ;
        RECT  0.105 0.200 0.210 0.280 ;
        RECT  0.105 0.980 0.210 1.060 ;
        RECT  0.035 0.200 0.105 1.060 ;
    END
END GBUFFD1BWP40

MACRO GBUFFD2BWP40
    CLASS CORE ;
    FOREIGN GBUFFD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.360 1.365 0.915 ;
        RECT  1.090 0.360 1.295 0.430 ;
        RECT  0.990 0.845 1.295 0.915 ;
        RECT  1.010 0.185 1.090 0.430 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.525 0.640 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.300 0.290 ;
        RECT  0.900 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.900 0.290 ;
        RECT  0.400 -0.115 0.800 0.115 ;
        RECT  0.300 -0.115 0.400 0.290 ;
        RECT  0.200 -0.115 0.300 0.115 ;
        RECT  0.100 -0.115 0.200 0.290 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.410 1.145 0.790 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.185 1.145 0.290 1.375 ;
        RECT  0.115 0.960 0.185 1.375 ;
        RECT  0.000 1.145 0.115 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.520 1.225 0.640 ;
        RECT  0.595 0.200 0.665 1.060 ;
        RECT  0.490 0.200 0.595 0.280 ;
        RECT  0.490 0.980 0.595 1.060 ;
    END
END GBUFFD2BWP40

MACRO GBUFFD3BWP40
    CLASS CORE ;
    FOREIGN GBUFFD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.276000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.370 1.365 0.920 ;
        RECT  1.085 0.370 1.295 0.440 ;
        RECT  0.665 0.850 1.295 0.920 ;
        RECT  1.015 0.185 1.085 0.440 ;
        RECT  0.610 0.370 1.015 0.440 ;
        RECT  0.565 0.850 0.665 1.060 ;
        RECT  0.540 0.200 0.610 0.440 ;
        RECT  0.490 0.980 0.565 1.060 ;
        RECT  0.490 0.200 0.540 0.280 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.265 0.355 0.385 0.485 ;
        RECT  0.175 0.355 0.265 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.115 1.400 0.115 ;
        RECT  1.200 -0.115 1.300 0.290 ;
        RECT  0.900 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.900 0.290 ;
        RECT  0.410 -0.115 0.800 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.410 1.145 0.790 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.125 0.520 1.225 0.640 ;
        RECT  0.495 0.545 1.125 0.615 ;
        RECT  0.425 0.545 0.495 0.780 ;
        RECT  0.105 0.710 0.425 0.780 ;
        RECT  0.105 0.200 0.210 0.280 ;
        RECT  0.105 0.980 0.210 1.060 ;
        RECT  0.035 0.200 0.105 1.060 ;
    END
END GBUFFD3BWP40

MACRO GBUFFD4BWP40
    CLASS CORE ;
    FOREIGN GBUFFD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.272000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.360 2.065 0.915 ;
        RECT  1.790 0.360 1.995 0.440 ;
        RECT  0.990 0.775 1.995 0.915 ;
        RECT  1.710 0.185 1.790 0.440 ;
        RECT  1.090 0.360 1.710 0.440 ;
        RECT  1.010 0.185 1.090 0.440 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.525 0.640 ;
        RECT  0.150 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.100 0.115 ;
        RECT  1.900 -0.115 2.000 0.290 ;
        RECT  1.600 -0.115 1.900 0.115 ;
        RECT  1.500 -0.115 1.600 0.290 ;
        RECT  1.300 -0.115 1.500 0.115 ;
        RECT  1.200 -0.115 1.300 0.290 ;
        RECT  0.900 -0.115 1.200 0.115 ;
        RECT  0.800 -0.115 0.900 0.290 ;
        RECT  0.610 -0.115 0.800 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.200 -0.115 0.490 0.115 ;
        RECT  0.100 -0.115 0.200 0.290 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.145 2.100 1.375 ;
        RECT  1.890 0.985 2.010 1.375 ;
        RECT  1.610 1.145 1.890 1.375 ;
        RECT  1.490 0.985 1.610 1.375 ;
        RECT  1.310 1.145 1.490 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.520 1.925 0.640 ;
        RECT  0.595 0.355 0.665 0.920 ;
        RECT  0.400 0.355 0.595 0.425 ;
        RECT  0.280 0.850 0.595 0.920 ;
        RECT  0.300 0.190 0.400 0.425 ;
    END
END GBUFFD4BWP40

MACRO GBUFFD8BWP40
    CLASS CORE ;
    FOREIGN GBUFFD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.544000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  2.595 0.305 3.045 0.935 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 1.225 0.640 ;
        RECT  0.160 0.495 0.245 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.100 -0.115 4.200 0.115 ;
        RECT  4.000 -0.115 4.100 0.290 ;
        RECT  3.700 -0.115 4.000 0.115 ;
        RECT  3.600 -0.115 3.700 0.290 ;
        RECT  3.400 -0.115 3.600 0.115 ;
        RECT  3.300 -0.115 3.400 0.290 ;
        RECT  3.000 -0.115 3.300 0.115 ;
        RECT  2.900 -0.115 3.000 0.290 ;
        RECT  2.700 -0.115 2.900 0.115 ;
        RECT  2.600 -0.115 2.700 0.290 ;
        RECT  2.300 -0.115 2.600 0.115 ;
        RECT  2.200 -0.115 2.300 0.290 ;
        RECT  2.000 -0.115 2.200 0.115 ;
        RECT  1.900 -0.115 2.000 0.290 ;
        RECT  1.600 -0.115 1.900 0.115 ;
        RECT  1.500 -0.115 1.600 0.290 ;
        RECT  1.310 -0.115 1.500 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.400 -0.115 0.790 0.115 ;
        RECT  0.300 -0.115 0.400 0.290 ;
        RECT  0.200 -0.115 0.300 0.115 ;
        RECT  0.100 -0.115 0.200 0.290 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.110 1.145 4.200 1.375 ;
        RECT  3.990 0.985 4.110 1.375 ;
        RECT  3.710 1.145 3.990 1.375 ;
        RECT  3.590 0.985 3.710 1.375 ;
        RECT  3.410 1.145 3.590 1.375 ;
        RECT  3.290 0.985 3.410 1.375 ;
        RECT  3.010 1.145 3.290 1.375 ;
        RECT  2.890 0.985 3.010 1.375 ;
        RECT  2.710 1.145 2.890 1.375 ;
        RECT  2.590 0.985 2.710 1.375 ;
        RECT  2.310 1.145 2.590 1.375 ;
        RECT  2.190 0.985 2.310 1.375 ;
        RECT  2.010 1.145 2.190 1.375 ;
        RECT  1.890 0.985 2.010 1.375 ;
        RECT  1.610 1.145 1.890 1.375 ;
        RECT  1.490 0.985 1.610 1.375 ;
        RECT  1.310 1.145 1.490 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.410 1.145 0.790 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.210 1.145 0.290 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.365 0.520 4.165 0.640 ;
        RECT  1.690 0.775 3.975 0.915 ;
        RECT  3.810 0.185 3.890 0.440 ;
        RECT  3.185 0.360 3.810 0.440 ;
        RECT  3.110 0.185 3.185 0.440 ;
        RECT  2.490 0.360 3.110 0.440 ;
        RECT  2.410 0.185 2.490 0.440 ;
        RECT  1.790 0.360 2.410 0.440 ;
        RECT  1.710 0.185 1.790 0.440 ;
        RECT  1.295 0.355 1.365 0.920 ;
        RECT  1.100 0.355 1.295 0.425 ;
        RECT  0.600 0.850 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  0.600 0.355 1.000 0.425 ;
        RECT  0.500 0.190 0.600 0.425 ;
        RECT  0.500 0.850 0.600 1.070 ;
        LAYER VIA1 ;
        RECT  2.880 0.365 2.950 0.435 ;
        RECT  2.880 0.805 2.950 0.875 ;
        RECT  2.650 0.365 2.720 0.435 ;
        RECT  2.650 0.805 2.720 0.875 ;
    END
END GBUFFD8BWP40

MACRO GDCAP10BWP40
    CLASS CORE ;
    FOREIGN GDCAP10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.690 -0.115 7.000 0.115 ;
        RECT  6.610 -0.115 6.690 0.300 ;
        RECT  6.490 -0.115 6.610 0.115 ;
        RECT  6.410 -0.115 6.490 0.300 ;
        RECT  5.990 -0.115 6.410 0.115 ;
        RECT  5.910 -0.115 5.990 0.300 ;
        RECT  5.790 -0.115 5.910 0.115 ;
        RECT  5.710 -0.115 5.790 0.300 ;
        RECT  5.290 -0.115 5.710 0.115 ;
        RECT  5.210 -0.115 5.290 0.300 ;
        RECT  5.090 -0.115 5.210 0.115 ;
        RECT  5.010 -0.115 5.090 0.300 ;
        RECT  4.590 -0.115 5.010 0.115 ;
        RECT  4.510 -0.115 4.590 0.300 ;
        RECT  4.390 -0.115 4.510 0.115 ;
        RECT  4.310 -0.115 4.390 0.300 ;
        RECT  3.890 -0.115 4.310 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.690 -0.115 3.810 0.115 ;
        RECT  3.610 -0.115 3.690 0.300 ;
        RECT  3.190 -0.115 3.610 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.910 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.910 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.900 1.145 7.000 1.375 ;
        RECT  6.810 0.850 6.900 1.375 ;
        RECT  6.590 0.850 6.810 0.920 ;
        RECT  6.190 1.145 6.810 1.375 ;
        RECT  6.110 0.850 6.190 1.375 ;
        RECT  5.890 0.850 6.110 0.920 ;
        RECT  5.490 1.145 6.110 1.375 ;
        RECT  5.410 0.850 5.490 1.375 ;
        RECT  5.190 0.850 5.410 0.920 ;
        RECT  4.790 1.145 5.410 1.375 ;
        RECT  4.710 0.850 4.790 1.375 ;
        RECT  4.490 0.850 4.710 0.920 ;
        RECT  4.090 1.145 4.710 1.375 ;
        RECT  4.010 0.850 4.090 1.375 ;
        RECT  3.790 0.850 4.010 0.920 ;
        RECT  3.390 1.145 4.010 1.375 ;
        RECT  3.310 0.850 3.390 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.690 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.690 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.800 0.190 6.910 0.450 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.555 0.380 6.800 0.450 ;
        RECT  6.500 0.710 6.745 0.780 ;
        RECT  6.470 0.380 6.555 0.640 ;
        RECT  6.390 0.710 6.500 1.070 ;
        RECT  6.210 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.390 0.780 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP10BWP40

MACRO GDCAP12BWP40
    CLASS CORE ;
    FOREIGN GDCAP12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.090 -0.115 8.400 0.115 ;
        RECT  8.010 -0.115 8.090 0.300 ;
        RECT  7.890 -0.115 8.010 0.115 ;
        RECT  7.810 -0.115 7.890 0.300 ;
        RECT  7.390 -0.115 7.810 0.115 ;
        RECT  7.310 -0.115 7.390 0.300 ;
        RECT  7.190 -0.115 7.310 0.115 ;
        RECT  7.100 -0.115 7.190 0.300 ;
        RECT  6.690 -0.115 7.100 0.115 ;
        RECT  6.610 -0.115 6.690 0.300 ;
        RECT  6.490 -0.115 6.610 0.115 ;
        RECT  6.410 -0.115 6.490 0.300 ;
        RECT  5.990 -0.115 6.410 0.115 ;
        RECT  5.910 -0.115 5.990 0.300 ;
        RECT  5.790 -0.115 5.910 0.115 ;
        RECT  5.710 -0.115 5.790 0.300 ;
        RECT  5.290 -0.115 5.710 0.115 ;
        RECT  5.210 -0.115 5.290 0.300 ;
        RECT  5.090 -0.115 5.210 0.115 ;
        RECT  5.010 -0.115 5.090 0.300 ;
        RECT  4.590 -0.115 5.010 0.115 ;
        RECT  4.510 -0.115 4.590 0.300 ;
        RECT  4.390 -0.115 4.510 0.115 ;
        RECT  4.310 -0.115 4.390 0.300 ;
        RECT  3.890 -0.115 4.310 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.690 -0.115 3.810 0.115 ;
        RECT  3.610 -0.115 3.690 0.300 ;
        RECT  3.190 -0.115 3.610 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.910 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.910 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.300 1.145 8.400 1.375 ;
        RECT  8.210 0.850 8.300 1.375 ;
        RECT  7.990 0.850 8.210 0.920 ;
        RECT  7.590 1.145 8.210 1.375 ;
        RECT  7.510 0.850 7.590 1.375 ;
        RECT  7.290 0.850 7.510 0.920 ;
        RECT  6.900 1.145 7.510 1.375 ;
        RECT  6.810 0.850 6.900 1.375 ;
        RECT  6.590 0.850 6.810 0.920 ;
        RECT  6.190 1.145 6.810 1.375 ;
        RECT  6.110 0.850 6.190 1.375 ;
        RECT  5.890 0.850 6.110 0.920 ;
        RECT  5.490 1.145 6.110 1.375 ;
        RECT  5.410 0.850 5.490 1.375 ;
        RECT  5.190 0.850 5.410 0.920 ;
        RECT  4.790 1.145 5.410 1.375 ;
        RECT  4.710 0.850 4.790 1.375 ;
        RECT  4.490 0.850 4.710 0.920 ;
        RECT  4.090 1.145 4.710 1.375 ;
        RECT  4.010 0.850 4.090 1.375 ;
        RECT  3.790 0.850 4.010 0.920 ;
        RECT  3.390 1.145 4.010 1.375 ;
        RECT  3.310 0.850 3.390 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.690 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.690 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.200 0.190 8.310 0.450 ;
        RECT  8.145 0.520 8.230 0.780 ;
        RECT  7.955 0.380 8.200 0.450 ;
        RECT  7.900 0.710 8.145 0.780 ;
        RECT  7.870 0.380 7.955 0.640 ;
        RECT  7.790 0.710 7.900 1.070 ;
        RECT  7.610 0.380 7.870 0.450 ;
        RECT  7.530 0.710 7.790 0.780 ;
        RECT  7.500 0.190 7.610 0.450 ;
        RECT  7.445 0.520 7.530 0.780 ;
        RECT  7.255 0.380 7.500 0.450 ;
        RECT  7.200 0.710 7.445 0.780 ;
        RECT  7.170 0.380 7.255 0.640 ;
        RECT  7.090 0.710 7.200 1.070 ;
        RECT  6.910 0.380 7.170 0.450 ;
        RECT  6.830 0.710 7.090 0.780 ;
        RECT  6.800 0.190 6.910 0.450 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.555 0.380 6.800 0.450 ;
        RECT  6.500 0.710 6.745 0.780 ;
        RECT  6.470 0.380 6.555 0.640 ;
        RECT  6.390 0.710 6.500 1.070 ;
        RECT  6.210 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.390 0.780 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP12BWP40

MACRO GDCAP2BWP40
    CLASS CORE ;
    FOREIGN GDCAP2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.400 1.375 ;
        RECT  1.210 0.850 1.300 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP2BWP40

MACRO GDCAP3BWP40
    CLASS CORE ;
    FOREIGN GDCAP3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 -0.115 2.100 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.145 2.100 1.375 ;
        RECT  1.910 0.850 2.000 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP3BWP40

MACRO GDCAP4BWP40
    CLASS CORE ;
    FOREIGN GDCAP4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.490 -0.115 2.800 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.145 2.800 1.375 ;
        RECT  2.610 0.850 2.700 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP4BWP40

MACRO GDCAP5BWP40
    CLASS CORE ;
    FOREIGN GDCAP5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 -0.115 3.500 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.900 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.900 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.145 3.500 1.375 ;
        RECT  3.310 0.850 3.400 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.700 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.700 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
    END
END GDCAP5BWP40

MACRO GDCAP6BWP40
    CLASS CORE ;
    FOREIGN GDCAP6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.890 -0.115 4.200 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.690 -0.115 3.810 0.115 ;
        RECT  3.610 -0.115 3.690 0.300 ;
        RECT  3.190 -0.115 3.610 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.910 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.910 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.100 1.145 4.200 1.375 ;
        RECT  4.010 0.850 4.100 1.375 ;
        RECT  3.790 0.850 4.010 0.920 ;
        RECT  3.390 1.145 4.010 1.375 ;
        RECT  3.310 0.850 3.390 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.690 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.690 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP6BWP40

MACRO GDCAP8BWP40
    CLASS CORE ;
    FOREIGN GDCAP8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.290 -0.115 5.600 0.115 ;
        RECT  5.210 -0.115 5.290 0.300 ;
        RECT  5.090 -0.115 5.210 0.115 ;
        RECT  5.010 -0.115 5.090 0.300 ;
        RECT  4.590 -0.115 5.010 0.115 ;
        RECT  4.510 -0.115 4.590 0.300 ;
        RECT  4.390 -0.115 4.510 0.115 ;
        RECT  4.310 -0.115 4.390 0.300 ;
        RECT  3.890 -0.115 4.310 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.690 -0.115 3.810 0.115 ;
        RECT  3.610 -0.115 3.690 0.300 ;
        RECT  3.190 -0.115 3.610 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.910 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.910 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.500 1.145 5.600 1.375 ;
        RECT  5.410 0.850 5.500 1.375 ;
        RECT  5.190 0.850 5.410 0.920 ;
        RECT  4.790 1.145 5.410 1.375 ;
        RECT  4.710 0.850 4.790 1.375 ;
        RECT  4.490 0.850 4.710 0.920 ;
        RECT  4.090 1.145 4.710 1.375 ;
        RECT  4.010 0.850 4.090 1.375 ;
        RECT  3.790 0.850 4.010 0.920 ;
        RECT  3.390 1.145 4.010 1.375 ;
        RECT  3.310 0.850 3.390 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.690 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.690 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP8BWP40

MACRO GDCAP9BWP40
    CLASS CORE ;
    FOREIGN GDCAP9BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.990 -0.115 6.300 0.115 ;
        RECT  5.910 -0.115 5.990 0.300 ;
        RECT  5.790 -0.115 5.910 0.115 ;
        RECT  5.700 -0.115 5.790 0.300 ;
        RECT  5.290 -0.115 5.700 0.115 ;
        RECT  5.210 -0.115 5.290 0.300 ;
        RECT  5.090 -0.115 5.210 0.115 ;
        RECT  5.010 -0.115 5.090 0.300 ;
        RECT  4.590 -0.115 5.010 0.115 ;
        RECT  4.510 -0.115 4.590 0.300 ;
        RECT  4.390 -0.115 4.510 0.115 ;
        RECT  4.310 -0.115 4.390 0.300 ;
        RECT  3.890 -0.115 4.310 0.115 ;
        RECT  3.810 -0.115 3.890 0.300 ;
        RECT  3.690 -0.115 3.810 0.115 ;
        RECT  3.610 -0.115 3.690 0.300 ;
        RECT  3.190 -0.115 3.610 0.115 ;
        RECT  3.110 -0.115 3.190 0.300 ;
        RECT  2.990 -0.115 3.110 0.115 ;
        RECT  2.910 -0.115 2.990 0.300 ;
        RECT  2.490 -0.115 2.910 0.115 ;
        RECT  2.410 -0.115 2.490 0.300 ;
        RECT  2.290 -0.115 2.410 0.115 ;
        RECT  2.210 -0.115 2.290 0.300 ;
        RECT  1.790 -0.115 2.210 0.115 ;
        RECT  1.710 -0.115 1.790 0.300 ;
        RECT  1.590 -0.115 1.710 0.115 ;
        RECT  1.510 -0.115 1.590 0.300 ;
        RECT  1.090 -0.115 1.510 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.890 -0.115 1.010 0.115 ;
        RECT  0.810 -0.115 0.890 0.300 ;
        RECT  0.390 -0.115 0.810 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.200 1.145 6.300 1.375 ;
        RECT  6.110 0.850 6.200 1.375 ;
        RECT  5.890 0.850 6.110 0.920 ;
        RECT  5.500 1.145 6.110 1.375 ;
        RECT  5.410 0.850 5.500 1.375 ;
        RECT  5.190 0.850 5.410 0.920 ;
        RECT  4.790 1.145 5.410 1.375 ;
        RECT  4.710 0.850 4.790 1.375 ;
        RECT  4.490 0.850 4.710 0.920 ;
        RECT  4.090 1.145 4.710 1.375 ;
        RECT  4.010 0.850 4.090 1.375 ;
        RECT  3.790 0.850 4.010 0.920 ;
        RECT  3.390 1.145 4.010 1.375 ;
        RECT  3.310 0.850 3.390 1.375 ;
        RECT  3.090 0.850 3.310 0.920 ;
        RECT  2.690 1.145 3.310 1.375 ;
        RECT  2.610 0.850 2.690 1.375 ;
        RECT  2.390 0.850 2.610 0.920 ;
        RECT  1.990 1.145 2.610 1.375 ;
        RECT  1.910 0.850 1.990 1.375 ;
        RECT  1.690 0.850 1.910 0.920 ;
        RECT  1.290 1.145 1.910 1.375 ;
        RECT  1.210 0.850 1.290 1.375 ;
        RECT  0.990 0.850 1.210 0.920 ;
        RECT  0.590 1.145 1.210 1.375 ;
        RECT  0.510 0.850 0.590 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAP9BWP40

MACRO GDCAPBWP40
    CLASS CORE ;
    FOREIGN GDCAPBWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.390 -0.115 0.700 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.190 -0.115 0.310 0.115 ;
        RECT  0.100 -0.115 0.190 0.300 ;
        RECT  0.000 -0.115 0.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.700 1.375 ;
        RECT  0.510 0.850 0.600 1.375 ;
        RECT  0.290 0.850 0.510 0.920 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GDCAPBWP40

MACRO GDFCNQD1BWP40
    CLASS CORE ;
    FOREIGN GDFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.205 5.565 1.055 ;
        RECT  5.390 0.205 5.495 0.275 ;
        RECT  5.390 0.985 5.495 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.960 0.385 1.410 0.455 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.635 0.385 0.765 ;
        RECT  0.175 0.495 0.260 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.400 0.385 4.330 0.455 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.310 -0.115 5.600 0.115 ;
        RECT  5.190 -0.115 5.310 0.275 ;
        RECT  4.385 -0.115 5.190 0.115 ;
        RECT  4.315 -0.115 4.385 0.300 ;
        RECT  2.985 -0.115 4.315 0.115 ;
        RECT  2.915 -0.115 2.985 0.300 ;
        RECT  2.485 -0.115 2.915 0.115 ;
        RECT  2.415 -0.115 2.485 0.300 ;
        RECT  0.885 -0.115 2.415 0.115 ;
        RECT  0.815 -0.115 0.885 0.300 ;
        RECT  0.410 -0.115 0.815 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.305 1.145 5.600 1.375 ;
        RECT  5.215 0.825 5.305 1.375 ;
        RECT  4.810 1.145 5.215 1.375 ;
        RECT  4.690 0.990 4.810 1.375 ;
        RECT  4.410 1.145 4.690 1.375 ;
        RECT  4.290 0.985 4.410 1.375 ;
        RECT  4.085 1.145 4.290 1.375 ;
        RECT  4.015 0.960 4.085 1.375 ;
        RECT  2.480 1.145 4.015 1.375 ;
        RECT  2.410 0.825 2.480 1.375 ;
        RECT  1.810 1.145 2.410 1.375 ;
        RECT  1.690 0.850 1.810 1.375 ;
        RECT  0.410 1.145 1.690 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.520 5.425 0.640 ;
        RECT  4.990 0.900 5.125 1.070 ;
        RECT  4.955 0.200 5.110 0.425 ;
        RECT  4.795 0.205 4.865 0.920 ;
        RECT  4.690 0.205 4.795 0.275 ;
        RECT  4.490 0.850 4.795 0.920 ;
        RECT  4.635 0.505 4.725 0.765 ;
        RECT  4.490 0.185 4.610 0.395 ;
        RECT  4.315 0.545 4.475 0.615 ;
        RECT  4.165 0.385 4.315 0.615 ;
        RECT  3.985 0.200 4.185 0.315 ;
        RECT  3.955 0.475 4.025 0.805 ;
        RECT  3.815 0.185 3.885 0.415 ;
        RECT  3.815 0.820 3.885 1.060 ;
        RECT  3.185 0.345 3.815 0.415 ;
        RECT  3.295 0.985 3.815 1.060 ;
        RECT  3.530 0.520 3.780 0.615 ;
        RECT  3.080 0.205 3.715 0.275 ;
        RECT  3.460 0.520 3.530 0.905 ;
        RECT  3.255 0.520 3.460 0.635 ;
        RECT  3.115 0.345 3.185 0.965 ;
        RECT  2.825 0.520 3.045 0.635 ;
        RECT  2.885 0.875 3.005 1.070 ;
        RECT  2.755 0.520 2.825 0.795 ;
        RECT  2.565 0.185 2.765 0.315 ;
        RECT  2.585 0.880 2.720 1.070 ;
        RECT  2.555 0.385 2.625 0.675 ;
        RECT  2.410 0.385 2.555 0.455 ;
        RECT  2.290 0.540 2.380 0.615 ;
        RECT  2.145 0.205 2.310 0.275 ;
        RECT  2.145 0.985 2.310 1.055 ;
        RECT  2.220 0.540 2.290 0.905 ;
        RECT  2.075 0.205 2.145 1.055 ;
        RECT  1.855 0.520 2.075 0.635 ;
        RECT  1.885 0.185 2.005 0.395 ;
        RECT  1.905 0.705 1.995 1.075 ;
        RECT  1.785 0.705 1.905 0.775 ;
        RECT  1.715 0.185 1.785 0.775 ;
        RECT  1.515 0.510 1.645 0.755 ;
        RECT  1.180 0.985 1.620 1.055 ;
        RECT  1.365 0.200 1.610 0.280 ;
        RECT  1.295 0.200 1.365 0.875 ;
        RECT  1.190 0.200 1.295 0.275 ;
        RECT  1.085 0.805 1.295 0.875 ;
        RECT  1.155 0.355 1.225 0.695 ;
        RECT  0.980 0.185 1.085 0.410 ;
        RECT  1.015 0.805 1.085 0.960 ;
        RECT  0.805 0.495 0.945 0.675 ;
        RECT  0.780 0.805 0.910 1.075 ;
        RECT  0.605 0.205 0.675 1.055 ;
        RECT  0.490 0.205 0.605 0.275 ;
        RECT  0.490 0.985 0.605 1.055 ;
        RECT  0.455 0.345 0.525 0.640 ;
        RECT  0.200 0.345 0.455 0.415 ;
        RECT  0.105 0.985 0.210 1.055 ;
        RECT  0.105 0.190 0.200 0.415 ;
        RECT  0.100 0.190 0.105 1.055 ;
        RECT  0.035 0.345 0.100 1.055 ;
        LAYER VIA1 ;
        RECT  5.020 0.945 5.090 1.015 ;
        RECT  4.980 0.245 5.050 0.315 ;
        RECT  4.655 0.665 4.725 0.735 ;
        RECT  4.210 0.385 4.280 0.455 ;
        RECT  4.045 0.245 4.115 0.315 ;
        RECT  3.955 0.525 4.025 0.595 ;
        RECT  3.460 0.805 3.530 0.875 ;
        RECT  3.115 0.665 3.185 0.735 ;
        RECT  2.915 0.945 2.985 1.015 ;
        RECT  2.755 0.665 2.825 0.735 ;
        RECT  2.625 0.245 2.695 0.315 ;
        RECT  2.610 0.945 2.680 1.015 ;
        RECT  2.450 0.385 2.520 0.455 ;
        RECT  2.220 0.805 2.290 0.875 ;
        RECT  1.915 0.945 1.985 1.015 ;
        RECT  1.910 0.245 1.980 0.315 ;
        RECT  1.550 0.665 1.620 0.735 ;
        RECT  1.200 0.805 1.270 0.875 ;
        RECT  1.155 0.385 1.225 0.455 ;
        RECT  0.865 0.525 0.935 0.595 ;
        RECT  0.820 0.945 0.890 1.015 ;
        RECT  0.605 0.665 0.675 0.735 ;
        RECT  0.455 0.475 0.525 0.545 ;
        LAYER M2 ;
        RECT  2.865 0.945 5.140 1.015 ;
        RECT  3.995 0.245 5.100 0.315 ;
        RECT  3.060 0.665 4.775 0.735 ;
        RECT  0.525 0.525 4.075 0.595 ;
        RECT  1.150 0.805 3.580 0.875 ;
        RECT  0.555 0.665 2.875 0.735 ;
        RECT  1.860 0.245 2.745 0.315 ;
        RECT  0.770 0.945 2.730 1.015 ;
        RECT  0.455 0.425 0.525 0.595 ;
    END
END GDFCNQD1BWP40

MACRO GDFCNQD2BWP40
    CLASS CORE ;
    FOREIGN GDFCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.565 0.205 5.845 0.275 ;
        RECT  5.565 0.930 5.845 1.055 ;
        RECT  5.495 0.205 5.565 1.055 ;
        RECT  5.390 0.205 5.495 0.275 ;
        RECT  5.390 0.930 5.495 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.960 0.385 1.410 0.455 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.635 0.385 0.765 ;
        RECT  0.175 0.495 0.260 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.400 0.385 4.330 0.455 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.185 -0.115 6.300 0.115 ;
        RECT  6.115 -0.115 6.185 0.305 ;
        RECT  5.985 -0.115 6.115 0.115 ;
        RECT  5.915 -0.115 5.985 0.300 ;
        RECT  5.310 -0.115 5.915 0.115 ;
        RECT  5.190 -0.115 5.310 0.275 ;
        RECT  4.385 -0.115 5.190 0.115 ;
        RECT  4.315 -0.115 4.385 0.300 ;
        RECT  2.985 -0.115 4.315 0.115 ;
        RECT  2.915 -0.115 2.985 0.300 ;
        RECT  2.485 -0.115 2.915 0.115 ;
        RECT  2.415 -0.115 2.485 0.300 ;
        RECT  0.885 -0.115 2.415 0.115 ;
        RECT  0.815 -0.115 0.885 0.300 ;
        RECT  0.410 -0.115 0.815 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.185 1.145 6.300 1.375 ;
        RECT  6.115 0.955 6.185 1.375 ;
        RECT  5.985 1.145 6.115 1.375 ;
        RECT  5.915 0.820 5.985 1.375 ;
        RECT  5.305 1.145 5.915 1.375 ;
        RECT  5.215 0.825 5.305 1.375 ;
        RECT  4.810 1.145 5.215 1.375 ;
        RECT  4.690 0.990 4.810 1.375 ;
        RECT  4.410 1.145 4.690 1.375 ;
        RECT  4.290 0.985 4.410 1.375 ;
        RECT  4.085 1.145 4.290 1.375 ;
        RECT  4.015 0.960 4.085 1.375 ;
        RECT  2.480 1.145 4.015 1.375 ;
        RECT  2.410 0.825 2.480 1.375 ;
        RECT  1.810 1.145 2.410 1.375 ;
        RECT  1.690 0.850 1.810 1.375 ;
        RECT  0.410 1.145 1.690 1.375 ;
        RECT  0.290 0.850 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.730 0.520 6.165 0.615 ;
        RECT  4.865 0.520 5.425 0.640 ;
        RECT  4.990 0.900 5.125 1.070 ;
        RECT  4.955 0.200 5.110 0.425 ;
        RECT  4.795 0.205 4.865 0.920 ;
        RECT  4.690 0.205 4.795 0.275 ;
        RECT  4.490 0.850 4.795 0.920 ;
        RECT  4.635 0.505 4.725 0.765 ;
        RECT  4.490 0.185 4.610 0.395 ;
        RECT  4.315 0.545 4.475 0.615 ;
        RECT  4.165 0.385 4.315 0.615 ;
        RECT  3.985 0.200 4.185 0.315 ;
        RECT  3.955 0.475 4.025 0.805 ;
        RECT  3.815 0.185 3.885 0.415 ;
        RECT  3.815 0.820 3.885 1.060 ;
        RECT  3.185 0.345 3.815 0.415 ;
        RECT  3.295 0.985 3.815 1.060 ;
        RECT  3.530 0.520 3.780 0.615 ;
        RECT  3.080 0.205 3.715 0.275 ;
        RECT  3.460 0.520 3.530 0.905 ;
        RECT  3.255 0.520 3.460 0.635 ;
        RECT  3.115 0.345 3.185 0.965 ;
        RECT  2.825 0.520 3.045 0.635 ;
        RECT  2.885 0.875 3.005 1.070 ;
        RECT  2.755 0.520 2.825 0.795 ;
        RECT  2.565 0.185 2.765 0.315 ;
        RECT  2.585 0.880 2.720 1.070 ;
        RECT  2.555 0.385 2.625 0.675 ;
        RECT  2.410 0.385 2.555 0.455 ;
        RECT  2.290 0.540 2.380 0.615 ;
        RECT  2.145 0.205 2.310 0.275 ;
        RECT  2.145 0.985 2.310 1.055 ;
        RECT  2.220 0.540 2.290 0.905 ;
        RECT  2.075 0.205 2.145 1.055 ;
        RECT  1.855 0.520 2.075 0.635 ;
        RECT  1.885 0.185 2.005 0.395 ;
        RECT  1.905 0.705 1.995 1.075 ;
        RECT  1.785 0.705 1.905 0.775 ;
        RECT  1.715 0.185 1.785 0.775 ;
        RECT  1.515 0.510 1.645 0.755 ;
        RECT  1.180 0.985 1.620 1.055 ;
        RECT  1.365 0.200 1.610 0.280 ;
        RECT  1.295 0.200 1.365 0.875 ;
        RECT  1.190 0.200 1.295 0.275 ;
        RECT  1.085 0.805 1.295 0.875 ;
        RECT  1.155 0.355 1.225 0.695 ;
        RECT  0.980 0.185 1.085 0.410 ;
        RECT  1.015 0.805 1.085 0.960 ;
        RECT  0.805 0.495 0.945 0.675 ;
        RECT  0.780 0.805 0.910 1.075 ;
        RECT  0.605 0.205 0.675 1.055 ;
        RECT  0.490 0.205 0.605 0.275 ;
        RECT  0.490 0.985 0.605 1.055 ;
        RECT  0.455 0.345 0.525 0.640 ;
        RECT  0.200 0.345 0.455 0.415 ;
        RECT  0.105 0.985 0.210 1.055 ;
        RECT  0.105 0.190 0.200 0.415 ;
        RECT  0.100 0.190 0.105 1.055 ;
        RECT  0.035 0.345 0.100 1.055 ;
        LAYER VIA1 ;
        RECT  5.875 0.525 5.945 0.595 ;
        RECT  5.195 0.525 5.265 0.595 ;
        RECT  5.020 0.945 5.090 1.015 ;
        RECT  4.980 0.245 5.050 0.315 ;
        RECT  4.655 0.665 4.725 0.735 ;
        RECT  4.210 0.385 4.280 0.455 ;
        RECT  4.045 0.245 4.115 0.315 ;
        RECT  3.955 0.525 4.025 0.595 ;
        RECT  3.460 0.805 3.530 0.875 ;
        RECT  3.115 0.665 3.185 0.735 ;
        RECT  2.915 0.945 2.985 1.015 ;
        RECT  2.755 0.665 2.825 0.735 ;
        RECT  2.625 0.245 2.695 0.315 ;
        RECT  2.610 0.945 2.680 1.015 ;
        RECT  2.450 0.385 2.520 0.455 ;
        RECT  2.220 0.805 2.290 0.875 ;
        RECT  1.915 0.945 1.985 1.015 ;
        RECT  1.910 0.245 1.980 0.315 ;
        RECT  1.550 0.665 1.620 0.735 ;
        RECT  1.200 0.805 1.270 0.875 ;
        RECT  1.155 0.385 1.225 0.455 ;
        RECT  0.865 0.525 0.935 0.595 ;
        RECT  0.820 0.945 0.890 1.015 ;
        RECT  0.605 0.665 0.675 0.735 ;
        RECT  0.455 0.475 0.525 0.545 ;
        LAYER M2 ;
        RECT  5.145 0.525 5.995 0.595 ;
        RECT  2.865 0.945 5.140 1.015 ;
        RECT  3.995 0.245 5.100 0.315 ;
        RECT  3.060 0.665 4.775 0.735 ;
        RECT  0.525 0.525 4.075 0.595 ;
        RECT  1.150 0.805 3.580 0.875 ;
        RECT  0.555 0.665 2.875 0.735 ;
        RECT  1.860 0.245 2.745 0.315 ;
        RECT  0.770 0.945 2.730 1.015 ;
        RECT  0.455 0.425 0.525 0.595 ;
    END
END GDFCNQD2BWP40

MACRO GDFQD1BWP40
    CLASS CORE ;
    FOREIGN GDFQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.205 5.565 1.055 ;
        RECT  5.390 0.205 5.495 0.275 ;
        RECT  5.390 0.985 5.495 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.190 0.665 1.695 0.735 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.355 0.385 0.485 ;
        RECT  0.175 0.355 0.245 0.695 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.310 -0.115 5.600 0.115 ;
        RECT  5.190 -0.115 5.310 0.275 ;
        RECT  4.610 -0.115 5.190 0.115 ;
        RECT  4.490 -0.115 4.610 0.275 ;
        RECT  4.385 -0.115 4.490 0.115 ;
        RECT  4.315 -0.115 4.385 0.300 ;
        RECT  3.385 -0.115 4.315 0.115 ;
        RECT  3.315 -0.115 3.385 0.300 ;
        RECT  3.185 -0.115 3.315 0.115 ;
        RECT  3.115 -0.115 3.185 0.300 ;
        RECT  2.510 -0.115 3.115 0.115 ;
        RECT  2.390 -0.115 2.510 0.275 ;
        RECT  2.010 -0.115 2.390 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  0.410 -0.115 1.890 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.145 5.600 1.375 ;
        RECT  5.190 0.850 5.310 1.375 ;
        RECT  4.610 1.145 5.190 1.375 ;
        RECT  4.490 0.850 4.610 1.375 ;
        RECT  4.385 1.145 4.490 1.375 ;
        RECT  4.315 0.960 4.385 1.375 ;
        RECT  4.110 1.145 4.315 1.375 ;
        RECT  3.990 0.990 4.110 1.375 ;
        RECT  2.510 1.145 3.990 1.375 ;
        RECT  2.390 0.850 2.510 1.375 ;
        RECT  1.085 1.145 2.390 1.375 ;
        RECT  1.015 0.825 1.085 1.375 ;
        RECT  0.910 1.145 1.015 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.385 1.145 0.790 1.375 ;
        RECT  0.315 0.825 0.385 1.375 ;
        RECT  0.000 1.145 0.315 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.355 0.355 5.425 0.655 ;
        RECT  5.110 0.355 5.355 0.425 ;
        RECT  5.075 0.510 5.175 0.770 ;
        RECT  5.005 0.205 5.110 0.425 ;
        RECT  5.005 0.985 5.110 1.055 ;
        RECT  4.990 0.205 5.005 1.055 ;
        RECT  4.935 0.355 4.990 1.055 ;
        RECT  4.725 0.570 4.935 0.640 ;
        RECT  4.795 0.190 4.865 0.485 ;
        RECT  4.690 0.930 4.865 1.055 ;
        RECT  4.700 0.190 4.795 0.290 ;
        RECT  4.375 0.520 4.725 0.640 ;
        RECT  4.095 0.190 4.165 0.485 ;
        RECT  4.025 0.780 4.140 0.875 ;
        RECT  4.000 0.190 4.095 0.290 ;
        RECT  3.955 0.520 4.025 0.875 ;
        RECT  3.885 0.190 3.900 0.290 ;
        RECT  3.815 0.190 3.885 0.455 ;
        RECT  3.815 0.825 3.885 1.065 ;
        RECT  3.800 0.190 3.815 0.290 ;
        RECT  3.185 0.385 3.815 0.455 ;
        RECT  3.290 0.975 3.815 1.065 ;
        RECT  3.665 0.525 3.745 0.635 ;
        RECT  3.480 0.190 3.700 0.315 ;
        RECT  3.335 0.525 3.665 0.595 ;
        RECT  3.255 0.525 3.335 0.635 ;
        RECT  3.115 0.385 3.185 0.945 ;
        RECT  2.975 0.355 3.045 0.680 ;
        RECT  2.905 0.195 3.010 0.275 ;
        RECT  2.895 0.860 3.005 1.070 ;
        RECT  2.835 0.195 2.905 0.395 ;
        RECT  2.695 0.205 2.765 1.055 ;
        RECT  2.590 0.205 2.695 0.275 ;
        RECT  2.590 0.985 2.695 1.055 ;
        RECT  2.535 0.355 2.625 0.640 ;
        RECT  2.260 0.520 2.360 0.765 ;
        RECT  2.180 0.985 2.310 1.055 ;
        RECT  2.180 0.190 2.300 0.350 ;
        RECT  2.110 0.190 2.180 1.055 ;
        RECT  1.890 0.985 2.110 1.055 ;
        RECT  1.925 0.520 1.995 0.905 ;
        RECT  1.855 0.520 1.925 0.640 ;
        RECT  1.505 0.850 1.810 0.920 ;
        RECT  1.695 0.190 1.800 0.400 ;
        RECT  1.645 0.635 1.785 0.765 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.505 0.205 1.610 0.275 ;
        RECT  1.190 0.990 1.610 1.060 ;
        RECT  1.435 0.205 1.505 0.920 ;
        RECT  1.190 0.205 1.435 0.275 ;
        RECT  1.170 0.355 1.260 0.640 ;
        RECT  0.875 0.520 1.170 0.640 ;
        RECT  0.785 0.195 1.105 0.315 ;
        RECT  0.595 0.205 0.665 1.055 ;
        RECT  0.490 0.205 0.595 0.275 ;
        RECT  0.490 0.985 0.595 1.055 ;
        RECT  0.455 0.495 0.525 0.905 ;
        RECT  0.105 0.205 0.210 0.275 ;
        RECT  0.105 0.800 0.200 1.070 ;
        RECT  0.100 0.205 0.105 1.070 ;
        RECT  0.035 0.205 0.100 0.880 ;
        LAYER VIA1 ;
        RECT  5.090 0.665 5.160 0.735 ;
        RECT  4.795 0.385 4.865 0.455 ;
        RECT  4.735 0.945 4.805 1.015 ;
        RECT  4.095 0.385 4.165 0.455 ;
        RECT  4.015 0.805 4.085 0.875 ;
        RECT  3.535 0.245 3.605 0.315 ;
        RECT  3.350 0.525 3.420 0.595 ;
        RECT  3.115 0.665 3.185 0.735 ;
        RECT  2.975 0.385 3.045 0.455 ;
        RECT  2.915 0.945 2.985 1.015 ;
        RECT  2.835 0.245 2.905 0.315 ;
        RECT  2.695 0.665 2.765 0.735 ;
        RECT  2.550 0.525 2.620 0.595 ;
        RECT  2.275 0.665 2.345 0.735 ;
        RECT  2.215 0.245 2.285 0.315 ;
        RECT  1.925 0.805 1.995 0.875 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.435 0.525 1.505 0.595 ;
        RECT  1.180 0.385 1.250 0.455 ;
        RECT  0.910 0.245 0.980 0.315 ;
        RECT  0.595 0.385 0.665 0.455 ;
        RECT  0.455 0.805 0.525 0.875 ;
        RECT  0.100 0.805 0.170 0.875 ;
        LAYER M2 ;
        RECT  3.065 0.665 5.210 0.735 ;
        RECT  4.045 0.385 4.915 0.455 ;
        RECT  2.865 0.945 4.855 1.015 ;
        RECT  0.050 0.805 4.135 0.875 ;
        RECT  2.785 0.245 3.655 0.315 ;
        RECT  1.385 0.525 3.470 0.595 ;
        RECT  0.545 0.385 3.095 0.455 ;
        RECT  2.225 0.665 2.815 0.735 ;
        RECT  0.860 0.245 2.335 0.315 ;
    END
END GDFQD1BWP40

MACRO GDFQD2BWP40
    CLASS CORE ;
    FOREIGN GDFQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Q
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.885 0.205 5.110 0.275 ;
        RECT  4.885 0.985 5.110 1.055 ;
        RECT  4.795 0.205 4.885 1.055 ;
        RECT  4.690 0.205 4.795 0.275 ;
        RECT  4.690 0.985 4.795 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.190 0.665 1.695 0.735 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.355 0.385 0.485 ;
        RECT  0.175 0.355 0.245 0.695 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.310 -0.115 5.600 0.115 ;
        RECT  5.190 -0.115 5.310 0.275 ;
        RECT  4.610 -0.115 5.190 0.115 ;
        RECT  4.490 -0.115 4.610 0.275 ;
        RECT  3.385 -0.115 4.490 0.115 ;
        RECT  3.315 -0.115 3.385 0.300 ;
        RECT  3.185 -0.115 3.315 0.115 ;
        RECT  3.115 -0.115 3.185 0.300 ;
        RECT  2.510 -0.115 3.115 0.115 ;
        RECT  2.390 -0.115 2.510 0.275 ;
        RECT  2.010 -0.115 2.390 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  0.410 -0.115 1.890 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.145 5.600 1.375 ;
        RECT  5.190 0.850 5.310 1.375 ;
        RECT  4.610 1.145 5.190 1.375 ;
        RECT  4.490 0.850 4.610 1.375 ;
        RECT  4.110 1.145 4.490 1.375 ;
        RECT  3.990 0.990 4.110 1.375 ;
        RECT  2.510 1.145 3.990 1.375 ;
        RECT  2.390 0.850 2.510 1.375 ;
        RECT  1.085 1.145 2.390 1.375 ;
        RECT  1.015 0.825 1.085 1.375 ;
        RECT  0.910 1.145 1.015 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.385 1.145 0.790 1.375 ;
        RECT  0.315 0.825 0.385 1.375 ;
        RECT  0.000 1.145 0.315 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.510 0.355 5.565 1.055 ;
        RECT  5.495 0.205 5.510 1.055 ;
        RECT  5.390 0.205 5.495 0.425 ;
        RECT  5.390 0.985 5.495 1.055 ;
        RECT  5.320 0.510 5.425 0.770 ;
        RECT  5.145 0.355 5.390 0.425 ;
        RECT  5.055 0.355 5.145 0.645 ;
        RECT  4.350 0.520 4.725 0.640 ;
        RECT  4.235 0.930 4.410 1.055 ;
        RECT  3.995 0.205 4.405 0.275 ;
        RECT  4.045 0.780 4.140 0.875 ;
        RECT  3.955 0.520 4.045 0.875 ;
        RECT  3.885 0.190 3.900 0.290 ;
        RECT  3.815 0.190 3.885 0.455 ;
        RECT  3.815 0.825 3.885 1.065 ;
        RECT  3.800 0.190 3.815 0.290 ;
        RECT  3.185 0.385 3.815 0.455 ;
        RECT  3.290 0.975 3.815 1.065 ;
        RECT  3.665 0.525 3.745 0.635 ;
        RECT  3.480 0.190 3.700 0.315 ;
        RECT  3.335 0.525 3.665 0.595 ;
        RECT  3.255 0.525 3.335 0.635 ;
        RECT  3.115 0.385 3.185 0.945 ;
        RECT  2.975 0.355 3.045 0.680 ;
        RECT  2.905 0.195 3.010 0.275 ;
        RECT  2.895 0.860 3.005 1.070 ;
        RECT  2.835 0.195 2.905 0.395 ;
        RECT  2.695 0.205 2.765 1.055 ;
        RECT  2.590 0.205 2.695 0.275 ;
        RECT  2.590 0.985 2.695 1.055 ;
        RECT  2.535 0.355 2.625 0.640 ;
        RECT  2.260 0.520 2.360 0.765 ;
        RECT  2.180 0.985 2.310 1.055 ;
        RECT  2.180 0.190 2.300 0.350 ;
        RECT  2.110 0.190 2.180 1.055 ;
        RECT  1.890 0.985 2.110 1.055 ;
        RECT  1.925 0.520 1.995 0.905 ;
        RECT  1.855 0.520 1.925 0.640 ;
        RECT  1.505 0.850 1.810 0.920 ;
        RECT  1.695 0.190 1.800 0.400 ;
        RECT  1.645 0.635 1.785 0.765 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.505 0.205 1.610 0.275 ;
        RECT  1.190 0.990 1.610 1.060 ;
        RECT  1.435 0.205 1.505 0.920 ;
        RECT  1.190 0.205 1.435 0.275 ;
        RECT  1.170 0.355 1.260 0.640 ;
        RECT  0.875 0.520 1.170 0.640 ;
        RECT  0.785 0.195 1.105 0.315 ;
        RECT  0.595 0.205 0.665 1.055 ;
        RECT  0.490 0.205 0.595 0.275 ;
        RECT  0.490 0.985 0.595 1.055 ;
        RECT  0.455 0.495 0.525 0.905 ;
        RECT  0.105 0.205 0.210 0.275 ;
        RECT  0.105 0.800 0.200 1.070 ;
        RECT  0.100 0.205 0.105 1.070 ;
        RECT  0.035 0.205 0.100 0.880 ;
        LAYER VIA1 ;
        RECT  5.330 0.665 5.400 0.735 ;
        RECT  5.075 0.525 5.145 0.595 ;
        RECT  4.525 0.525 4.595 0.595 ;
        RECT  4.280 0.945 4.350 1.015 ;
        RECT  4.015 0.805 4.085 0.875 ;
        RECT  3.535 0.245 3.605 0.315 ;
        RECT  3.350 0.525 3.420 0.595 ;
        RECT  3.115 0.665 3.185 0.735 ;
        RECT  2.975 0.385 3.045 0.455 ;
        RECT  2.915 0.945 2.985 1.015 ;
        RECT  2.835 0.245 2.905 0.315 ;
        RECT  2.695 0.665 2.765 0.735 ;
        RECT  2.550 0.525 2.620 0.595 ;
        RECT  2.275 0.665 2.345 0.735 ;
        RECT  2.215 0.245 2.285 0.315 ;
        RECT  1.925 0.805 1.995 0.875 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.435 0.525 1.505 0.595 ;
        RECT  1.180 0.385 1.250 0.455 ;
        RECT  0.910 0.245 0.980 0.315 ;
        RECT  0.595 0.385 0.665 0.455 ;
        RECT  0.455 0.805 0.525 0.875 ;
        RECT  0.100 0.805 0.170 0.875 ;
        LAYER M2 ;
        RECT  3.065 0.665 5.450 0.735 ;
        RECT  4.475 0.525 5.195 0.595 ;
        RECT  2.865 0.945 4.400 1.015 ;
        RECT  0.050 0.805 4.135 0.875 ;
        RECT  2.785 0.245 3.655 0.315 ;
        RECT  1.385 0.525 3.470 0.595 ;
        RECT  0.545 0.385 3.095 0.455 ;
        RECT  2.225 0.665 2.815 0.735 ;
        RECT  0.860 0.245 2.335 0.315 ;
    END
END GDFQD2BWP40

MACRO GFILL10BWP40
    CLASS CORE ;
    FOREIGN GFILL10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 7.000 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 7.000 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.800 0.190 6.910 0.450 ;
        RECT  6.800 0.850 6.910 1.070 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.555 0.380 6.800 0.450 ;
        RECT  6.590 0.850 6.800 0.920 ;
        RECT  6.500 0.710 6.745 0.780 ;
        RECT  6.370 0.200 6.710 0.280 ;
        RECT  6.470 0.380 6.555 0.640 ;
        RECT  6.390 0.710 6.500 1.070 ;
        RECT  6.210 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.390 0.780 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.100 0.850 6.210 1.070 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.890 0.850 6.100 0.920 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.670 0.200 6.010 0.280 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.400 0.850 5.510 1.070 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.190 0.850 5.400 0.920 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  4.970 0.200 5.310 0.280 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.700 0.850 4.810 1.070 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.490 0.850 4.700 0.920 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.270 0.200 4.610 0.280 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  4.000 0.850 4.110 1.070 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.570 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL10BWP40

MACRO GFILL12BWP40
    CLASS CORE ;
    FOREIGN GFILL12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 8.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 8.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.200 0.190 8.310 0.450 ;
        RECT  8.200 0.850 8.310 1.070 ;
        RECT  8.145 0.520 8.230 0.780 ;
        RECT  7.955 0.380 8.200 0.450 ;
        RECT  7.990 0.850 8.200 0.920 ;
        RECT  7.900 0.710 8.145 0.780 ;
        RECT  7.770 0.200 8.110 0.280 ;
        RECT  7.870 0.380 7.955 0.640 ;
        RECT  7.790 0.710 7.900 1.070 ;
        RECT  7.610 0.380 7.870 0.450 ;
        RECT  7.530 0.710 7.790 0.780 ;
        RECT  7.500 0.190 7.610 0.450 ;
        RECT  7.500 0.850 7.610 1.070 ;
        RECT  7.445 0.520 7.530 0.780 ;
        RECT  7.255 0.380 7.500 0.450 ;
        RECT  7.290 0.850 7.500 0.920 ;
        RECT  7.200 0.710 7.445 0.780 ;
        RECT  7.070 0.200 7.410 0.280 ;
        RECT  7.170 0.380 7.255 0.640 ;
        RECT  7.090 0.710 7.200 1.070 ;
        RECT  6.910 0.380 7.170 0.450 ;
        RECT  6.830 0.710 7.090 0.780 ;
        RECT  6.800 0.190 6.910 0.450 ;
        RECT  6.800 0.850 6.910 1.070 ;
        RECT  6.745 0.520 6.830 0.780 ;
        RECT  6.555 0.380 6.800 0.450 ;
        RECT  6.590 0.850 6.800 0.920 ;
        RECT  6.500 0.710 6.745 0.780 ;
        RECT  6.370 0.200 6.710 0.280 ;
        RECT  6.470 0.380 6.555 0.640 ;
        RECT  6.390 0.710 6.500 1.070 ;
        RECT  6.210 0.380 6.470 0.450 ;
        RECT  6.130 0.710 6.390 0.780 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.100 0.850 6.210 1.070 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.890 0.850 6.100 0.920 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.670 0.200 6.010 0.280 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.400 0.850 5.510 1.070 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.190 0.850 5.400 0.920 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  4.970 0.200 5.310 0.280 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.700 0.850 4.810 1.070 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.490 0.850 4.700 0.920 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.270 0.200 4.610 0.280 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  4.000 0.850 4.110 1.070 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.570 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL12BWP40

MACRO GFILL2BWP40
    CLASS CORE ;
    FOREIGN GFILL2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.400 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 1.400 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL2BWP40

MACRO GFILL3BWP40
    CLASS CORE ;
    FOREIGN GFILL3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.100 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL3BWP40

MACRO GFILL4BWP40
    CLASS CORE ;
    FOREIGN GFILL4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 2.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 2.800 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL4BWP40

MACRO GFILL5BWP40
    CLASS CORE ;
    FOREIGN GFILL5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 3.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 3.500 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL5BWP40

MACRO GFILL6BWP40
    CLASS CORE ;
    FOREIGN GFILL6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 4.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 4.200 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  4.000 0.850 4.110 1.070 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.570 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL6BWP40

MACRO GFILL8BWP40
    CLASS CORE ;
    FOREIGN GFILL8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 5.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 5.600 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.400 0.850 5.510 1.070 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.190 0.850 5.400 0.920 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  4.970 0.200 5.310 0.280 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.700 0.850 4.810 1.070 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.490 0.850 4.700 0.920 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.270 0.200 4.610 0.280 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  4.000 0.850 4.110 1.070 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.570 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL8BWP40

MACRO GFILL9BWP40
    CLASS CORE ;
    FOREIGN GFILL9BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 6.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 6.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.100 0.190 6.210 0.450 ;
        RECT  6.100 0.850 6.210 1.070 ;
        RECT  6.045 0.520 6.130 0.780 ;
        RECT  5.855 0.380 6.100 0.450 ;
        RECT  5.890 0.850 6.100 0.920 ;
        RECT  5.800 0.710 6.045 0.780 ;
        RECT  5.670 0.200 6.010 0.280 ;
        RECT  5.770 0.380 5.855 0.640 ;
        RECT  5.690 0.710 5.800 1.070 ;
        RECT  5.510 0.380 5.770 0.450 ;
        RECT  5.430 0.710 5.690 0.780 ;
        RECT  5.400 0.190 5.510 0.450 ;
        RECT  5.400 0.850 5.510 1.070 ;
        RECT  5.345 0.520 5.430 0.780 ;
        RECT  5.155 0.380 5.400 0.450 ;
        RECT  5.190 0.850 5.400 0.920 ;
        RECT  5.100 0.710 5.345 0.780 ;
        RECT  4.970 0.200 5.310 0.280 ;
        RECT  5.070 0.380 5.155 0.640 ;
        RECT  4.990 0.710 5.100 1.070 ;
        RECT  4.810 0.380 5.070 0.450 ;
        RECT  4.730 0.710 4.990 0.780 ;
        RECT  4.700 0.190 4.810 0.450 ;
        RECT  4.700 0.850 4.810 1.070 ;
        RECT  4.645 0.520 4.730 0.780 ;
        RECT  4.455 0.380 4.700 0.450 ;
        RECT  4.490 0.850 4.700 0.920 ;
        RECT  4.400 0.710 4.645 0.780 ;
        RECT  4.270 0.200 4.610 0.280 ;
        RECT  4.370 0.380 4.455 0.640 ;
        RECT  4.290 0.710 4.400 1.070 ;
        RECT  4.110 0.380 4.370 0.450 ;
        RECT  4.030 0.710 4.290 0.780 ;
        RECT  4.000 0.190 4.110 0.450 ;
        RECT  4.000 0.850 4.110 1.070 ;
        RECT  3.945 0.520 4.030 0.780 ;
        RECT  3.755 0.380 4.000 0.450 ;
        RECT  3.790 0.850 4.000 0.920 ;
        RECT  3.700 0.710 3.945 0.780 ;
        RECT  3.570 0.200 3.910 0.280 ;
        RECT  3.670 0.380 3.755 0.640 ;
        RECT  3.590 0.710 3.700 1.070 ;
        RECT  3.410 0.380 3.670 0.450 ;
        RECT  3.330 0.710 3.590 0.780 ;
        RECT  3.300 0.190 3.410 0.450 ;
        RECT  3.300 0.850 3.410 1.070 ;
        RECT  3.245 0.520 3.330 0.780 ;
        RECT  3.055 0.380 3.300 0.450 ;
        RECT  3.090 0.850 3.300 0.920 ;
        RECT  3.000 0.710 3.245 0.780 ;
        RECT  2.870 0.200 3.210 0.280 ;
        RECT  2.970 0.380 3.055 0.640 ;
        RECT  2.890 0.710 3.000 1.070 ;
        RECT  2.710 0.380 2.970 0.450 ;
        RECT  2.630 0.710 2.890 0.780 ;
        RECT  2.600 0.190 2.710 0.450 ;
        RECT  2.600 0.850 2.710 1.070 ;
        RECT  2.545 0.520 2.630 0.780 ;
        RECT  2.355 0.380 2.600 0.450 ;
        RECT  2.390 0.850 2.600 0.920 ;
        RECT  2.300 0.710 2.545 0.780 ;
        RECT  2.170 0.200 2.510 0.280 ;
        RECT  2.270 0.380 2.355 0.640 ;
        RECT  2.190 0.710 2.300 1.070 ;
        RECT  2.010 0.380 2.270 0.450 ;
        RECT  1.930 0.710 2.190 0.780 ;
        RECT  1.900 0.190 2.010 0.450 ;
        RECT  1.900 0.850 2.010 1.070 ;
        RECT  1.845 0.520 1.930 0.780 ;
        RECT  1.655 0.380 1.900 0.450 ;
        RECT  1.690 0.850 1.900 0.920 ;
        RECT  1.600 0.710 1.845 0.780 ;
        RECT  1.470 0.200 1.810 0.280 ;
        RECT  1.570 0.380 1.655 0.640 ;
        RECT  1.490 0.710 1.600 1.070 ;
        RECT  1.310 0.380 1.570 0.450 ;
        RECT  1.230 0.710 1.490 0.780 ;
        RECT  1.200 0.190 1.310 0.450 ;
        RECT  1.200 0.850 1.310 1.070 ;
        RECT  1.145 0.520 1.230 0.780 ;
        RECT  0.955 0.380 1.200 0.450 ;
        RECT  0.990 0.850 1.200 0.920 ;
        RECT  0.900 0.710 1.145 0.780 ;
        RECT  0.770 0.200 1.110 0.280 ;
        RECT  0.870 0.380 0.955 0.640 ;
        RECT  0.790 0.710 0.900 1.070 ;
        RECT  0.610 0.380 0.870 0.450 ;
        RECT  0.530 0.710 0.790 0.780 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILL9BWP40

MACRO GFILLBWP40
    CLASS CORE ;
    FOREIGN GFILLBWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 0.700 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.145 0.700 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.500 0.190 0.610 0.450 ;
        RECT  0.500 0.850 0.610 1.070 ;
        RECT  0.445 0.520 0.530 0.780 ;
        RECT  0.255 0.380 0.500 0.450 ;
        RECT  0.290 0.850 0.500 0.920 ;
        RECT  0.200 0.710 0.445 0.780 ;
        RECT  0.070 0.200 0.410 0.280 ;
        RECT  0.170 0.380 0.255 0.640 ;
        RECT  0.090 0.710 0.200 1.070 ;
    END
END GFILLBWP40

MACRO GINVD1BWP40
    CLASS CORE ;
    FOREIGN GINVD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.200 0.290 ;
        RECT  0.105 0.970 0.200 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.530 0.765 ;
        RECT  0.175 0.495 0.455 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 -0.115 0.700 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.390 -0.115 0.490 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 0.700 1.375 ;
        RECT  0.500 0.970 0.600 1.375 ;
        RECT  0.410 1.145 0.500 1.375 ;
        RECT  0.290 0.845 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
END GINVD1BWP40

MACRO GINVD2BWP40
    CLASS CORE ;
    FOREIGN GINVD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.845 0.420 0.920 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.275 0.495 0.530 0.645 ;
        RECT  0.175 0.495 0.275 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 -0.115 0.700 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.145 0.700 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
END GINVD2BWP40

MACRO GINVD3BWP40
    CLASS CORE ;
    FOREIGN GINVD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.276000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.190 0.900 0.415 ;
        RECT  0.810 0.775 0.890 1.075 ;
        RECT  0.105 0.775 0.810 0.920 ;
        RECT  0.405 0.345 0.735 0.415 ;
        RECT  0.300 0.190 0.405 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.230 0.765 ;
        RECT  0.175 0.495 1.155 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  1.090 -0.115 1.190 0.115 ;
        RECT  1.010 -0.115 1.090 0.320 ;
        RECT  0.610 -0.115 1.010 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.400 1.375 ;
        RECT  1.200 0.970 1.300 1.375 ;
        RECT  1.110 1.145 1.200 1.375 ;
        RECT  0.990 0.845 1.110 1.375 ;
        RECT  0.610 1.145 0.990 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
END GINVD3BWP40

MACRO GINVD4BWP40
    CLASS CORE ;
    FOREIGN GINVD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.272000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.345 1.365 0.920 ;
        RECT  1.100 0.345 1.295 0.415 ;
        RECT  0.105 0.775 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.300 0.190 0.400 0.415 ;
        RECT  0.105 0.345 0.300 0.415 ;
        RECT  0.035 0.345 0.105 0.920 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.225 0.640 ;
        RECT  0.735 0.355 0.805 0.640 ;
        RECT  0.175 0.495 0.735 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.615 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.615 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
END GINVD4BWP40

MACRO GINVD8BWP40
    CLASS CORE ;
    FOREIGN GINVD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.544000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  1.195 0.285 1.645 0.935 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 2.625 0.640 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 -0.115 2.800 0.115 ;
        RECT  2.590 -0.115 2.710 0.275 ;
        RECT  2.310 -0.115 2.590 0.115 ;
        RECT  2.190 -0.115 2.310 0.275 ;
        RECT  2.010 -0.115 2.190 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  1.610 -0.115 1.890 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  1.310 -0.115 1.490 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.710 1.145 2.800 1.375 ;
        RECT  2.590 0.990 2.710 1.375 ;
        RECT  2.310 1.145 2.590 1.375 ;
        RECT  2.185 0.990 2.310 1.375 ;
        RECT  2.010 1.145 2.185 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.610 1.145 1.890 1.375 ;
        RECT  1.490 0.990 1.610 1.375 ;
        RECT  1.310 1.145 1.490 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.785 0.990 0.910 1.375 ;
        RECT  0.615 1.145 0.785 1.375 ;
        RECT  0.490 0.990 0.615 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.240 0.775 2.555 0.920 ;
        RECT  2.400 0.190 2.500 0.415 ;
        RECT  1.800 0.345 2.400 0.415 ;
        RECT  1.700 0.190 1.800 0.415 ;
        RECT  1.100 0.345 1.700 0.415 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.400 0.345 1.000 0.415 ;
        RECT  0.300 0.190 0.400 0.415 ;
        LAYER VIA1 ;
        RECT  1.480 0.345 1.550 0.415 ;
        RECT  1.480 0.805 1.550 0.875 ;
        RECT  1.250 0.345 1.320 0.415 ;
        RECT  1.250 0.805 1.320 0.875 ;
    END
END GINVD8BWP40

MACRO GMUX2D1BWP40
    CLASS CORE ;
    FOREIGN GMUX2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.205 0.290 ;
        RECT  0.105 0.970 0.200 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.815 0.665 1.975 0.735 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.665 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.670 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.145 2.100 1.375 ;
        RECT  1.740 0.835 1.810 1.375 ;
        RECT  1.700 0.835 1.740 0.935 ;
        RECT  0.410 1.145 1.740 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.005 0.355 2.065 1.070 ;
        RECT  1.995 0.190 2.005 1.070 ;
        RECT  1.900 0.190 1.995 0.425 ;
        RECT  1.890 0.970 1.995 1.070 ;
        RECT  1.835 0.495 1.925 0.765 ;
        RECT  1.225 0.355 1.900 0.425 ;
        RECT  1.190 0.200 1.610 0.275 ;
        RECT  1.500 0.775 1.600 1.075 ;
        RECT  1.200 0.775 1.300 1.075 ;
        RECT  1.155 0.355 1.225 0.660 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.425 ;
        RECT  0.335 0.355 1.000 0.425 ;
        RECT  0.855 0.495 0.945 0.765 ;
        RECT  0.490 0.200 0.910 0.275 ;
        RECT  0.800 0.845 0.900 1.075 ;
        RECT  0.500 0.775 0.600 1.070 ;
        RECT  0.265 0.355 0.335 0.640 ;
        RECT  0.175 0.520 0.265 0.640 ;
        LAYER VIA1 ;
        RECT  1.855 0.665 1.925 0.735 ;
        RECT  1.520 0.945 1.590 1.015 ;
        RECT  1.215 0.805 1.285 0.875 ;
        RECT  0.865 0.665 0.935 0.735 ;
        RECT  0.815 0.945 0.885 1.015 ;
        RECT  0.515 0.805 0.585 0.875 ;
        LAYER M2 ;
        RECT  0.765 0.945 1.640 1.015 ;
        RECT  0.465 0.805 1.335 0.875 ;
    END
END GMUX2D1BWP40

MACRO GMUX2D2BWP40
    CLASS CORE ;
    FOREIGN GMUX2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.195 0.910 0.275 ;
        RECT  0.805 0.970 0.910 1.065 ;
        RECT  0.735 0.195 0.805 1.065 ;
        RECT  0.490 0.195 0.735 0.275 ;
        RECT  0.490 0.970 0.735 1.065 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.515 0.665 2.675 0.735 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.220 0.525 1.965 0.595 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.370 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.390 -0.115 0.990 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.210 -0.115 0.310 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.110 1.145 2.440 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.395 1.145 0.990 1.375 ;
        RECT  0.305 0.810 0.395 1.375 ;
        RECT  0.210 1.145 0.305 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.705 0.355 2.765 1.070 ;
        RECT  2.695 0.190 2.705 1.070 ;
        RECT  2.600 0.190 2.695 0.425 ;
        RECT  2.590 0.970 2.695 1.070 ;
        RECT  2.535 0.495 2.625 0.765 ;
        RECT  1.925 0.355 2.600 0.425 ;
        RECT  1.890 0.200 2.310 0.275 ;
        RECT  2.200 0.775 2.300 1.075 ;
        RECT  1.900 0.775 2.000 1.075 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.425 ;
        RECT  1.035 0.355 1.700 0.425 ;
        RECT  1.555 0.495 1.645 0.765 ;
        RECT  1.190 0.200 1.610 0.275 ;
        RECT  1.500 0.845 1.600 1.075 ;
        RECT  1.135 0.495 1.365 0.625 ;
        RECT  1.200 0.775 1.300 1.070 ;
        RECT  0.965 0.355 1.035 0.640 ;
        RECT  0.875 0.520 0.965 0.640 ;
        RECT  0.115 0.495 0.565 0.625 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.220 0.945 2.290 1.015 ;
        RECT  1.915 0.805 1.985 0.875 ;
        RECT  1.565 0.665 1.635 0.735 ;
        RECT  1.515 0.945 1.585 1.015 ;
        RECT  1.270 0.525 1.340 0.595 ;
        RECT  1.215 0.805 1.285 0.875 ;
        RECT  0.915 0.525 0.985 0.595 ;
        RECT  0.310 0.525 0.380 0.595 ;
        LAYER M2 ;
        RECT  1.465 0.945 2.340 1.015 ;
        RECT  1.165 0.805 2.035 0.875 ;
        RECT  0.260 0.525 1.035 0.595 ;
    END
END GMUX2D2BWP40

MACRO GMUX2ND1BWP40
    CLASS CORE ;
    FOREIGN GMUX2ND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.200 0.290 ;
        RECT  0.105 0.970 0.200 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.525 0.665 2.675 0.735 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.940 0.525 1.390 0.595 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.090 0.525 2.540 0.595 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.390 -0.115 0.990 0.115 ;
        RECT  0.310 -0.115 0.390 0.300 ;
        RECT  0.000 -0.115 0.310 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.290 1.145 2.440 1.375 ;
        RECT  1.210 0.940 1.290 1.375 ;
        RECT  0.890 1.145 1.210 1.375 ;
        RECT  0.810 0.940 0.890 1.375 ;
        RECT  0.410 1.145 0.810 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.705 0.355 2.765 1.070 ;
        RECT  2.695 0.190 2.705 1.070 ;
        RECT  2.600 0.190 2.695 0.425 ;
        RECT  2.600 0.970 2.695 1.070 ;
        RECT  2.535 0.495 2.625 0.765 ;
        RECT  1.925 0.355 2.600 0.425 ;
        RECT  2.135 0.495 2.370 0.625 ;
        RECT  1.890 0.200 2.310 0.275 ;
        RECT  2.200 0.775 2.300 1.075 ;
        RECT  1.900 0.775 2.000 1.075 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.560 0.495 1.645 0.765 ;
        RECT  1.250 0.200 1.610 0.275 ;
        RECT  1.500 0.845 1.600 1.075 ;
        RECT  1.180 0.200 1.250 0.415 ;
        RECT  0.805 0.495 1.250 0.625 ;
        RECT  0.900 0.345 1.180 0.415 ;
        RECT  1.000 0.775 1.100 1.045 ;
        RECT  0.800 0.190 0.900 0.415 ;
        RECT  0.635 0.355 0.705 0.615 ;
        RECT  0.430 0.545 0.635 0.615 ;
        RECT  0.555 0.185 0.605 0.290 ;
        RECT  0.560 0.970 0.605 1.070 ;
        RECT  0.490 0.695 0.560 1.070 ;
        RECT  0.485 0.185 0.555 0.440 ;
        RECT  0.245 0.695 0.490 0.765 ;
        RECT  0.245 0.370 0.485 0.440 ;
        RECT  0.175 0.370 0.245 0.765 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.220 0.945 2.290 1.015 ;
        RECT  2.195 0.525 2.265 0.595 ;
        RECT  1.915 0.805 1.985 0.875 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.575 0.665 1.645 0.735 ;
        RECT  1.515 0.945 1.585 1.015 ;
        RECT  1.020 0.525 1.090 0.595 ;
        RECT  1.015 0.805 1.085 0.875 ;
        RECT  0.635 0.385 0.705 0.455 ;
        LAYER M2 ;
        RECT  1.465 0.945 2.340 1.015 ;
        RECT  0.965 0.805 2.035 0.875 ;
        RECT  0.585 0.385 1.835 0.455 ;
    END
END GMUX2ND1BWP40

MACRO GMUX2ND2BWP40
    CLASS CORE ;
    FOREIGN GMUX2ND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.200 0.910 0.290 ;
        RECT  0.805 0.980 0.910 1.060 ;
        RECT  0.735 0.200 0.805 1.060 ;
        RECT  0.490 0.200 0.735 0.290 ;
        RECT  0.490 0.980 0.735 1.060 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.225 0.665 3.375 0.735 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.495 1.950 0.625 ;
        RECT  1.560 0.495 1.645 0.765 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 3.070 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.210 -0.115 3.500 0.115 ;
        RECT  3.090 -0.115 3.210 0.270 ;
        RECT  1.810 -0.115 3.090 0.115 ;
        RECT  1.690 -0.115 1.810 0.275 ;
        RECT  1.090 -0.115 1.690 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.390 -0.115 1.010 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.210 -0.115 0.310 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.145 3.500 1.375 ;
        RECT  3.140 0.835 3.210 1.375 ;
        RECT  3.100 0.835 3.140 0.935 ;
        RECT  1.990 1.145 3.140 1.375 ;
        RECT  1.910 0.940 1.990 1.375 ;
        RECT  1.590 1.145 1.910 1.375 ;
        RECT  1.510 0.940 1.590 1.375 ;
        RECT  1.110 1.145 1.510 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.200 1.145 0.990 1.375 ;
        RECT  0.200 0.850 0.410 0.920 ;
        RECT  0.100 0.850 0.200 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.405 0.355 3.465 1.070 ;
        RECT  3.395 0.190 3.405 1.070 ;
        RECT  3.300 0.190 3.395 0.425 ;
        RECT  3.300 0.970 3.395 1.070 ;
        RECT  3.235 0.495 3.325 0.765 ;
        RECT  2.625 0.355 3.300 0.425 ;
        RECT  2.590 0.200 3.010 0.275 ;
        RECT  2.900 0.775 3.000 1.075 ;
        RECT  2.600 0.775 2.700 1.075 ;
        RECT  2.555 0.355 2.625 0.660 ;
        RECT  2.485 0.190 2.500 0.290 ;
        RECT  2.415 0.190 2.485 0.965 ;
        RECT  2.400 0.190 2.415 0.290 ;
        RECT  2.260 0.495 2.345 0.765 ;
        RECT  1.950 0.200 2.310 0.275 ;
        RECT  2.200 0.845 2.300 1.075 ;
        RECT  1.880 0.200 1.950 0.415 ;
        RECT  1.600 0.345 1.880 0.415 ;
        RECT  1.715 0.775 1.800 1.045 ;
        RECT  1.500 0.190 1.600 0.415 ;
        RECT  1.335 0.355 1.405 0.615 ;
        RECT  1.130 0.545 1.335 0.615 ;
        RECT  1.255 0.185 1.305 0.290 ;
        RECT  1.260 0.970 1.305 1.070 ;
        RECT  1.190 0.695 1.260 1.070 ;
        RECT  1.185 0.185 1.255 0.440 ;
        RECT  0.945 0.695 1.190 0.765 ;
        RECT  0.945 0.370 1.185 0.440 ;
        RECT  0.875 0.370 0.945 0.765 ;
        RECT  0.135 0.495 0.555 0.655 ;
        LAYER VIA1 ;
        RECT  3.255 0.665 3.325 0.735 ;
        RECT  2.920 0.945 2.990 1.015 ;
        RECT  2.615 0.805 2.685 0.875 ;
        RECT  2.415 0.385 2.485 0.455 ;
        RECT  2.275 0.665 2.345 0.735 ;
        RECT  2.215 0.945 2.285 1.015 ;
        RECT  1.725 0.805 1.795 0.875 ;
        RECT  1.335 0.385 1.405 0.455 ;
        RECT  0.875 0.525 0.945 0.595 ;
        RECT  0.365 0.525 0.435 0.595 ;
        LAYER M2 ;
        RECT  2.165 0.945 3.040 1.015 ;
        RECT  1.675 0.805 2.735 0.875 ;
        RECT  1.285 0.385 2.535 0.455 ;
        RECT  0.285 0.525 0.995 0.595 ;
    END
END GMUX2ND2BWP40

MACRO GND2D1BWP40
    CLASS CORE ;
    FOREIGN GND2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.137750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.190 0.665 0.920 ;
        RECT  0.500 0.190 0.595 0.290 ;
        RECT  0.290 0.845 0.595 0.920 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.145 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.210 -0.115 0.700 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.145 0.700 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.300 0.190 0.400 0.410 ;
    END
END GND2D1BWP40

MACRO GND2D2BWP40
    CLASS CORE ;
    FOREIGN GND2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.212500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.850 1.120 0.920 ;
        RECT  0.595 0.355 0.700 0.920 ;
        RECT  0.400 0.355 0.595 0.425 ;
        RECT  0.280 0.850 0.595 0.920 ;
        RECT  0.300 0.190 0.400 0.425 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        RECT  0.165 0.495 0.435 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  0.840 0.495 1.155 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 1.400 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.000 -0.115 0.990 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.190 1.300 0.425 ;
        RECT  0.910 0.355 1.200 0.425 ;
        RECT  0.840 0.205 0.910 0.425 ;
        RECT  0.490 0.205 0.840 0.275 ;
        RECT  0.100 0.190 0.200 0.415 ;
        LAYER VIA1 ;
        RECT  0.840 0.245 0.910 0.315 ;
        RECT  0.115 0.245 0.185 0.315 ;
        LAYER M2 ;
        RECT  0.065 0.245 0.960 0.315 ;
    END
END GND2D2BWP40

MACRO GND3D1BWP40
    CLASS CORE ;
    FOREIGN GND3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.214250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.850 1.110 0.920 ;
        RECT  0.105 0.190 0.200 0.290 ;
        RECT  0.035 0.190 0.105 0.920 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.495 0.385 0.765 ;
        RECT  0.175 0.495 0.295 0.650 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.570 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.245 0.625 ;
        RECT  0.865 0.495 0.945 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.000 -0.115 0.790 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.600 0.345 1.000 0.415 ;
        RECT  0.500 0.190 0.600 0.415 ;
        RECT  0.300 0.190 0.400 0.410 ;
    END
END GND3D1BWP40

MACRO GND3D2BWP40
    CLASS CORE ;
    FOREIGN GND3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.352000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.850 1.815 0.920 ;
        RECT  0.595 0.190 0.665 0.920 ;
        RECT  0.500 0.190 0.595 0.290 ;
        RECT  0.105 0.850 0.595 0.920 ;
        RECT  0.105 0.190 0.200 0.290 ;
        RECT  0.035 0.190 0.105 0.920 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        RECT  0.265 0.635 0.435 0.765 ;
        RECT  0.175 0.495 0.265 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.245 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.495 1.930 0.765 ;
        RECT  1.575 0.495 1.840 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 -0.115 2.100 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  1.610 -0.115 1.890 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  0.000 -0.115 1.490 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.145 2.100 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.610 1.145 1.890 1.375 ;
        RECT  1.490 0.990 1.610 1.375 ;
        RECT  1.310 1.145 1.490 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.990 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.700 0.190 1.800 0.415 ;
        RECT  1.445 0.345 1.700 0.415 ;
        RECT  1.365 0.345 1.445 0.780 ;
        RECT  1.300 0.345 1.365 0.415 ;
        RECT  0.805 0.710 1.365 0.780 ;
        RECT  1.200 0.190 1.300 0.415 ;
        RECT  1.000 0.190 1.100 0.415 ;
        RECT  0.805 0.190 0.900 0.290 ;
        RECT  0.735 0.190 0.805 0.780 ;
        RECT  0.300 0.190 0.400 0.410 ;
        LAYER VIA1 ;
        RECT  1.015 0.245 1.085 0.315 ;
        RECT  0.315 0.245 0.385 0.315 ;
        LAYER M2 ;
        RECT  0.265 0.245 1.145 0.315 ;
    END
END GND3D2BWP40

MACRO GNR2D1BWP40
    CLASS CORE ;
    FOREIGN GNR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.700 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.138250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.500 0.970 0.595 1.070 ;
        RECT  0.300 0.190 0.400 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.650 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.650 ;
        RECT  0.035 0.355 0.105 0.650 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.610 -0.115 0.700 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.145 0.700 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.850 0.410 1.070 ;
    END
END GNR2D1BWP40

MACRO GNR2D2BWP40
    CLASS CORE ;
    FOREIGN GNR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.195500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.195 1.110 0.280 ;
        RECT  0.990 0.195 1.085 0.415 ;
        RECT  0.665 0.345 0.990 0.415 ;
        RECT  0.595 0.345 0.665 0.915 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.290 0.845 0.595 0.915 ;
        RECT  0.300 0.190 0.400 0.415 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.525 0.765 ;
        RECT  0.135 0.495 0.445 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.250 0.630 ;
        RECT  0.830 0.495 1.155 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  0.990 0.850 1.110 1.375 ;
        RECT  0.000 1.145 0.990 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.710 1.300 1.070 ;
        RECT  0.910 0.710 1.200 0.780 ;
        RECT  0.840 0.710 0.910 1.055 ;
        RECT  0.090 0.985 0.840 1.055 ;
    END
END GNR2D2BWP40

MACRO GNR3D1BWP40
    CLASS CORE ;
    FOREIGN GNR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.197750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  0.400 0.345 1.000 0.425 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.105 0.345 0.300 0.425 ;
        RECT  0.105 0.970 0.245 1.070 ;
        RECT  0.035 0.345 0.105 1.070 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  0.850 0.495 1.155 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.000 1.145 0.790 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.850 1.120 0.920 ;
        RECT  0.640 0.850 0.720 1.055 ;
        RECT  0.490 0.985 0.640 1.055 ;
        RECT  0.315 0.770 0.400 1.055 ;
    END
END GNR3D1BWP40

MACRO GNR3D2BWP40
    CLASS CORE ;
    FOREIGN GNR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.336000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.190 1.800 0.425 ;
        RECT  1.100 0.345 1.700 0.425 ;
        RECT  1.000 0.190 1.100 0.425 ;
        RECT  0.400 0.345 1.000 0.425 ;
        RECT  0.105 0.990 0.610 1.060 ;
        RECT  0.300 0.190 0.400 0.425 ;
        RECT  0.105 0.345 0.300 0.425 ;
        RECT  0.035 0.345 0.105 1.060 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.495 1.930 0.640 ;
        RECT  1.575 0.495 1.645 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.280 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.175 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 -0.115 2.100 0.115 ;
        RECT  1.890 -0.115 2.010 0.275 ;
        RECT  1.610 -0.115 1.890 0.115 ;
        RECT  1.490 -0.115 1.610 0.275 ;
        RECT  1.310 -0.115 1.490 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.145 2.100 1.375 ;
        RECT  1.890 0.990 2.010 1.375 ;
        RECT  1.610 1.145 1.890 1.375 ;
        RECT  1.490 0.990 1.610 1.375 ;
        RECT  0.000 1.145 1.490 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.320 0.850 1.815 0.920 ;
        RECT  1.250 0.850 1.320 1.060 ;
        RECT  0.790 0.990 1.250 1.060 ;
        RECT  0.290 0.850 1.120 0.920 ;
    END
END GNR3D2BWP40

MACRO GOAI21D1BWP40
    CLASS CORE ;
    FOREIGN GOAI21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.277750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M2 ;
        RECT  0.075 0.245 0.715 0.315 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  0.945 0.665 1.155 0.765 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 0.245 0.780 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.445 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.000 -0.115 0.790 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.985 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.210 1.145 0.790 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.685 0.850 1.130 0.920 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.485 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.595 0.190 0.685 1.055 ;
        RECT  0.500 0.190 0.595 0.290 ;
        RECT  0.490 0.985 0.595 1.055 ;
        RECT  0.290 0.850 0.410 1.060 ;
        RECT  0.385 0.190 0.400 0.290 ;
        RECT  0.315 0.190 0.385 0.485 ;
        RECT  0.300 0.190 0.315 0.290 ;
        RECT  0.100 0.190 0.210 0.415 ;
        LAYER VIA1 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.595 0.245 0.665 0.315 ;
        RECT  0.315 0.385 0.385 0.455 ;
        RECT  0.125 0.245 0.195 0.315 ;
        LAYER M2 ;
        RECT  0.265 0.385 1.135 0.455 ;
    END
END GOAI21D1BWP40

MACRO GOAI21D2BWP40
    CLASS CORE ;
    FOREIGN GOAI21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.353000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.990 2.065 1.060 ;
        RECT  1.700 0.190 1.800 0.415 ;
        RECT  1.505 0.345 1.700 0.415 ;
        RECT  1.435 0.345 1.505 1.060 ;
        RECT  1.205 0.775 1.435 0.920 ;
        RECT  0.665 0.845 1.205 0.920 ;
        RECT  0.595 0.355 0.665 0.920 ;
        RECT  0.400 0.355 0.595 0.425 ;
        RECT  0.300 0.190 0.400 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.965 0.495 1.240 0.640 ;
        RECT  0.875 0.495 0.965 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.525 0.640 ;
        RECT  0.035 0.495 0.115 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.495 2.065 0.765 ;
        RECT  1.575 0.495 1.985 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.110 -0.115 2.100 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.000 -0.115 0.990 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 2.100 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.990 0.910 1.375 ;
        RECT  0.610 1.145 0.790 1.375 ;
        RECT  0.490 0.990 0.610 1.375 ;
        RECT  0.210 1.145 0.490 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.190 2.000 0.415 ;
        RECT  1.690 0.735 1.810 0.920 ;
        RECT  1.260 0.205 1.610 0.275 ;
        RECT  1.190 0.205 1.260 0.425 ;
        RECT  0.910 0.355 1.190 0.425 ;
        RECT  0.840 0.205 0.910 0.425 ;
        RECT  0.470 0.205 0.840 0.275 ;
        RECT  0.290 0.735 0.410 0.920 ;
        RECT  0.100 0.190 0.200 0.415 ;
        LAYER VIA1 ;
        RECT  1.915 0.245 1.985 0.315 ;
        RECT  1.715 0.805 1.785 0.875 ;
        RECT  1.190 0.245 1.260 0.315 ;
        RECT  0.315 0.805 0.385 0.875 ;
        RECT  0.115 0.245 0.185 0.315 ;
        LAYER M2 ;
        RECT  0.065 0.245 2.035 0.315 ;
        RECT  0.265 0.805 1.835 0.875 ;
    END
END GOAI21D2BWP40

MACRO GOR2D1BWP40
    CLASS CORE ;
    FOREIGN GOR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.190 1.365 1.070 ;
        RECT  1.200 0.190 1.295 0.290 ;
        RECT  1.200 0.970 1.295 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.315 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.090 0.300 ;
        RECT  0.885 -0.115 1.010 0.115 ;
        RECT  0.815 -0.115 0.885 0.300 ;
        RECT  0.610 -0.115 0.815 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 1.145 1.400 1.375 ;
        RECT  0.885 0.850 1.130 0.920 ;
        RECT  0.815 0.850 0.885 1.375 ;
        RECT  0.210 1.145 0.815 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.500 1.225 0.780 ;
        RECT  0.945 0.710 1.155 0.780 ;
        RECT  0.875 0.500 0.945 0.780 ;
        RECT  0.665 0.710 0.875 0.780 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.500 0.970 0.595 1.070 ;
        RECT  0.290 0.845 0.410 1.055 ;
        RECT  0.300 0.190 0.400 0.415 ;
    END
END GOR2D1BWP40

MACRO GOR2D2BWP40
    CLASS CORE ;
    FOREIGN GOR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.350 1.365 0.920 ;
        RECT  1.100 0.350 1.295 0.420 ;
        RECT  0.980 0.850 1.295 0.920 ;
        RECT  1.000 0.190 1.100 0.420 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.315 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 -0.115 1.400 0.115 ;
        RECT  1.190 -0.115 1.310 0.275 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.275 ;
        RECT  0.610 -0.115 0.790 0.115 ;
        RECT  0.490 -0.115 0.610 0.275 ;
        RECT  0.210 -0.115 0.490 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.145 1.400 1.375 ;
        RECT  1.190 0.990 1.310 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.210 1.145 0.790 1.375 ;
        RECT  0.090 0.985 0.210 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.520 1.225 0.640 ;
        RECT  0.595 0.345 0.665 1.070 ;
        RECT  0.400 0.345 0.595 0.415 ;
        RECT  0.500 0.970 0.595 1.070 ;
        RECT  0.290 0.845 0.410 1.055 ;
        RECT  0.300 0.190 0.400 0.415 ;
    END
END GOR2D2BWP40

MACRO GSDFCNQD1BWP40
    CLASS CORE ;
    FOREIGN GSDFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN SI
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.325 0.525 0.860 0.595 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.065 0.665 0.580 0.735 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.295 0.205 8.365 1.055 ;
        RECT  8.190 0.205 8.295 0.275 ;
        RECT  8.155 0.940 8.295 1.055 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.370 0.525 1.860 0.595 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  4.070 0.245 4.605 0.315 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  3.350 0.385 7.225 0.455 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.110 -0.115 8.400 0.115 ;
        RECT  7.990 -0.115 8.110 0.275 ;
        RECT  7.210 -0.115 7.990 0.115 ;
        RECT  7.090 -0.115 7.210 0.270 ;
        RECT  5.080 -0.115 7.090 0.115 ;
        RECT  4.980 -0.115 5.080 0.300 ;
        RECT  4.610 -0.115 4.980 0.115 ;
        RECT  4.490 -0.115 4.610 0.270 ;
        RECT  3.210 -0.115 4.490 0.115 ;
        RECT  3.090 -0.115 3.210 0.270 ;
        RECT  1.985 -0.115 3.090 0.115 ;
        RECT  1.915 -0.115 1.985 0.300 ;
        RECT  1.810 -0.115 1.915 0.115 ;
        RECT  1.685 -0.115 1.810 0.275 ;
        RECT  0.400 -0.115 1.685 0.115 ;
        RECT  0.300 -0.115 0.400 0.290 ;
        RECT  0.000 -0.115 0.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.085 1.145 8.400 1.375 ;
        RECT  8.015 0.825 8.085 1.375 ;
        RECT  7.610 1.145 8.015 1.375 ;
        RECT  7.490 0.990 7.610 1.375 ;
        RECT  7.210 1.145 7.490 1.375 ;
        RECT  7.090 0.985 7.210 1.375 ;
        RECT  6.910 1.145 7.090 1.375 ;
        RECT  6.790 0.990 6.910 1.375 ;
        RECT  6.685 1.145 6.790 1.375 ;
        RECT  6.615 0.825 6.685 1.375 ;
        RECT  5.500 1.145 6.615 1.375 ;
        RECT  5.400 0.970 5.500 1.375 ;
        RECT  5.300 1.145 5.400 1.375 ;
        RECT  5.200 0.835 5.300 1.375 ;
        RECT  5.100 1.145 5.200 1.375 ;
        RECT  5.000 0.970 5.100 1.375 ;
        RECT  4.610 1.145 5.000 1.375 ;
        RECT  4.490 0.855 4.610 1.375 ;
        RECT  4.080 1.145 4.490 1.375 ;
        RECT  3.995 0.950 4.080 1.375 ;
        RECT  3.890 1.145 3.995 1.375 ;
        RECT  3.815 0.825 3.890 1.375 ;
        RECT  3.210 1.145 3.815 1.375 ;
        RECT  3.090 0.850 3.210 1.375 ;
        RECT  1.985 1.145 3.090 1.375 ;
        RECT  1.915 0.960 1.985 1.375 ;
        RECT  1.810 1.145 1.915 1.375 ;
        RECT  1.690 0.855 1.810 1.375 ;
        RECT  0.415 1.145 1.690 1.375 ;
        RECT  0.290 0.855 0.415 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.945 0.520 8.225 0.640 ;
        RECT  7.875 0.520 7.945 0.820 ;
        RECT  7.790 0.900 7.925 1.070 ;
        RECT  7.805 0.200 7.910 0.280 ;
        RECT  7.665 0.730 7.875 0.820 ;
        RECT  7.735 0.200 7.805 0.640 ;
        RECT  7.595 0.205 7.665 0.920 ;
        RECT  7.490 0.205 7.595 0.275 ;
        RECT  7.290 0.850 7.595 0.920 ;
        RECT  7.435 0.505 7.525 0.765 ;
        RECT  7.290 0.185 7.410 0.395 ;
        RECT  7.170 0.545 7.285 0.615 ;
        RECT  7.100 0.355 7.170 0.615 ;
        RECT  6.765 0.200 6.910 0.280 ;
        RECT  6.765 0.530 6.860 0.625 ;
        RECT  6.695 0.200 6.765 0.625 ;
        RECT  6.585 0.200 6.695 0.280 ;
        RECT  6.455 0.495 6.545 0.905 ;
        RECT  6.380 0.190 6.515 0.290 ;
        RECT  6.080 0.985 6.510 1.055 ;
        RECT  5.985 0.205 6.380 0.290 ;
        RECT  6.145 0.805 6.305 0.875 ;
        RECT  6.055 0.475 6.145 0.875 ;
        RECT  5.915 0.205 5.985 0.965 ;
        RECT  5.505 0.205 5.915 0.290 ;
        RECT  5.645 0.520 5.845 0.635 ;
        RECT  5.685 0.875 5.805 1.070 ;
        RECT  5.575 0.385 5.645 0.635 ;
        RECT  5.180 0.385 5.575 0.455 ;
        RECT  5.500 0.780 5.550 0.900 ;
        RECT  5.400 0.190 5.505 0.290 ;
        RECT  5.430 0.525 5.500 0.900 ;
        RECT  5.330 0.525 5.430 0.640 ;
        RECT  5.150 0.195 5.330 0.315 ;
        RECT  5.100 0.385 5.180 0.635 ;
        RECT  4.885 0.520 5.100 0.635 ;
        RECT  4.815 0.205 4.885 1.055 ;
        RECT  4.680 0.205 4.815 0.275 ;
        RECT  4.680 0.985 4.815 1.055 ;
        RECT  4.650 0.355 4.725 0.770 ;
        RECT  4.400 0.355 4.650 0.425 ;
        RECT  4.410 0.700 4.650 0.770 ;
        RECT  4.230 0.525 4.510 0.620 ;
        RECT  4.300 0.700 4.410 1.070 ;
        RECT  4.300 0.185 4.400 0.425 ;
        RECT  4.160 0.205 4.230 0.620 ;
        RECT  3.990 0.185 4.090 0.295 ;
        RECT  3.960 0.405 4.030 0.640 ;
        RECT  3.895 0.200 3.990 0.295 ;
        RECT  3.705 0.405 3.960 0.475 ;
        RECT  3.775 0.200 3.895 0.335 ;
        RECT  3.725 0.545 3.770 0.695 ;
        RECT  3.650 0.545 3.725 0.780 ;
        RECT  3.290 0.945 3.715 1.065 ;
        RECT  3.635 0.195 3.705 0.475 ;
        RECT  3.185 0.710 3.650 0.780 ;
        RECT  3.290 0.195 3.635 0.300 ;
        RECT  3.430 0.370 3.525 0.465 ;
        RECT  3.330 0.370 3.430 0.640 ;
        RECT  3.260 0.520 3.330 0.640 ;
        RECT  3.110 0.370 3.185 0.780 ;
        RECT  3.010 0.370 3.110 0.440 ;
        RECT  3.020 0.515 3.040 0.640 ;
        RECT  2.950 0.515 3.020 0.905 ;
        RECT  2.890 0.200 3.010 0.440 ;
        RECT  2.880 0.985 3.010 1.055 ;
        RECT  2.880 0.370 2.890 0.440 ;
        RECT  2.810 0.370 2.880 1.055 ;
        RECT  2.570 0.195 2.760 0.315 ;
        RECT  2.555 0.925 2.740 1.070 ;
        RECT  2.555 0.480 2.685 0.695 ;
        RECT  2.485 0.185 2.500 0.285 ;
        RECT  2.415 0.185 2.485 0.960 ;
        RECT  2.400 0.185 2.415 0.285 ;
        RECT  2.225 0.525 2.345 0.785 ;
        RECT  2.175 0.195 2.310 0.455 ;
        RECT  2.135 0.980 2.310 1.060 ;
        RECT  2.065 0.695 2.135 1.060 ;
        RECT  1.735 0.695 2.065 0.765 ;
        RECT  1.550 0.525 1.950 0.625 ;
        RECT  1.460 0.980 1.610 1.050 ;
        RECT  1.460 0.205 1.605 0.275 ;
        RECT  1.390 0.205 1.460 1.050 ;
        RECT  1.180 0.205 1.390 0.275 ;
        RECT  1.200 0.785 1.300 1.070 ;
        RECT  1.180 0.345 1.270 0.615 ;
        RECT  1.130 0.525 1.180 0.615 ;
        RECT  1.000 0.770 1.110 1.075 ;
        RECT  0.975 0.185 1.100 0.385 ;
        RECT  0.880 0.470 0.975 0.700 ;
        RECT  0.485 0.195 0.905 0.290 ;
        RECT  0.810 0.960 0.900 1.070 ;
        RECT  0.670 0.470 0.880 0.540 ;
        RECT  0.740 0.635 0.810 1.070 ;
        RECT  0.595 0.470 0.670 0.785 ;
        RECT  0.500 0.855 0.610 1.070 ;
        RECT  0.265 0.715 0.595 0.785 ;
        RECT  0.455 0.370 0.525 0.635 ;
        RECT  0.390 0.370 0.455 0.440 ;
        RECT  0.175 0.525 0.265 0.785 ;
        RECT  0.105 0.190 0.210 0.455 ;
        RECT  0.105 0.855 0.210 1.070 ;
        RECT  0.100 0.190 0.105 1.070 ;
        RECT  0.035 0.380 0.100 0.930 ;
        LAYER VIA1 ;
        RECT  7.820 0.945 7.890 1.015 ;
        RECT  7.735 0.245 7.805 0.315 ;
        RECT  7.445 0.665 7.515 0.735 ;
        RECT  7.100 0.385 7.170 0.455 ;
        RECT  6.695 0.245 6.765 0.315 ;
        RECT  6.475 0.525 6.545 0.595 ;
        RECT  6.185 0.805 6.255 0.875 ;
        RECT  5.915 0.665 5.985 0.735 ;
        RECT  5.715 0.945 5.785 1.015 ;
        RECT  5.455 0.805 5.525 0.875 ;
        RECT  4.815 0.665 4.885 0.735 ;
        RECT  4.655 0.525 4.725 0.595 ;
        RECT  4.160 0.245 4.230 0.315 ;
        RECT  3.800 0.245 3.870 0.315 ;
        RECT  3.475 0.945 3.545 1.015 ;
        RECT  3.400 0.385 3.470 0.455 ;
        RECT  2.950 0.805 3.020 0.875 ;
        RECT  2.635 0.245 2.705 0.315 ;
        RECT  2.625 0.945 2.695 1.015 ;
        RECT  2.560 0.525 2.630 0.595 ;
        RECT  2.415 0.805 2.485 0.875 ;
        RECT  2.245 0.665 2.315 0.735 ;
        RECT  2.210 0.385 2.280 0.455 ;
        RECT  1.785 0.695 1.855 0.765 ;
        RECT  1.610 0.525 1.680 0.595 ;
        RECT  1.390 0.665 1.460 0.735 ;
        RECT  1.210 0.945 1.280 1.015 ;
        RECT  1.180 0.385 1.250 0.455 ;
        RECT  1.020 0.805 1.090 0.875 ;
        RECT  1.015 0.245 1.085 0.315 ;
        RECT  0.740 0.665 0.810 0.735 ;
        RECT  0.530 0.945 0.600 1.015 ;
        RECT  0.455 0.525 0.525 0.595 ;
        RECT  0.175 0.665 0.245 0.735 ;
        RECT  0.110 0.385 0.180 0.455 ;
        LAYER M2 ;
        RECT  5.665 0.945 7.940 1.015 ;
        RECT  6.645 0.245 7.855 0.315 ;
        RECT  5.860 0.665 7.565 0.735 ;
        RECT  2.510 0.525 6.595 0.595 ;
        RECT  2.365 0.805 6.305 0.875 ;
        RECT  2.195 0.665 4.950 0.735 ;
        RECT  2.950 0.245 3.940 0.315 ;
        RECT  2.095 0.945 3.595 1.015 ;
        RECT  2.880 0.245 2.950 0.455 ;
        RECT  2.095 0.385 2.880 0.455 ;
        RECT  0.965 0.245 2.775 0.315 ;
        RECT  2.025 0.385 2.095 1.015 ;
        RECT  1.690 0.695 1.925 0.765 ;
        RECT  1.620 0.695 1.690 0.875 ;
        RECT  0.970 0.805 1.620 0.875 ;
        RECT  0.690 0.665 1.520 0.735 ;
        RECT  0.480 0.945 1.330 1.015 ;
        RECT  0.060 0.385 1.310 0.455 ;
    END
END GSDFCNQD1BWP40

MACRO GXNR2D1BWP40
    CLASS CORE ;
    FOREIGN GXNR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.190 0.205 0.290 ;
        RECT  0.105 0.970 0.200 1.070 ;
        RECT  0.035 0.190 0.105 1.070 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  0.815 0.665 1.975 0.735 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.275 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.145 2.100 1.375 ;
        RECT  1.740 0.835 1.810 1.375 ;
        RECT  1.700 0.835 1.740 0.935 ;
        RECT  0.410 1.145 1.740 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.005 0.355 2.065 1.070 ;
        RECT  1.995 0.190 2.005 1.070 ;
        RECT  1.900 0.190 1.995 0.425 ;
        RECT  1.900 0.970 1.995 1.070 ;
        RECT  1.835 0.495 1.925 0.765 ;
        RECT  1.225 0.355 1.900 0.425 ;
        RECT  1.365 0.545 1.670 0.615 ;
        RECT  1.190 0.200 1.610 0.275 ;
        RECT  1.500 0.775 1.600 1.075 ;
        RECT  1.295 0.545 1.365 1.055 ;
        RECT  1.190 0.985 1.295 1.055 ;
        RECT  1.155 0.355 1.225 0.660 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.855 0.495 0.945 0.765 ;
        RECT  0.605 0.200 0.675 1.055 ;
        RECT  0.490 0.200 0.605 0.275 ;
        RECT  0.490 0.985 0.605 1.055 ;
        RECT  0.265 0.355 0.335 0.640 ;
        RECT  0.175 0.520 0.265 0.640 ;
        RECT  0.675 0.200 0.910 0.275 ;
        RECT  0.800 0.845 0.900 1.075 ;
        LAYER VIA1 ;
        RECT  1.855 0.665 1.925 0.735 ;
        RECT  1.520 0.945 1.590 1.015 ;
        RECT  1.295 0.805 1.365 0.875 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.865 0.665 0.935 0.735 ;
        RECT  0.815 0.945 0.885 1.015 ;
        RECT  0.605 0.805 0.675 0.875 ;
        RECT  0.265 0.385 0.335 0.455 ;
        LAYER M2 ;
        RECT  0.765 0.945 1.640 1.015 ;
        RECT  0.555 0.805 1.415 0.875 ;
        RECT  0.215 0.385 1.135 0.455 ;
    END
END GXNR2D1BWP40

MACRO GXNR2D2BWP40
    CLASS CORE ;
    FOREIGN GXNR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN ZN
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.200 0.910 0.290 ;
        RECT  0.665 0.970 0.910 1.060 ;
        RECT  0.595 0.200 0.665 1.060 ;
        RECT  0.490 0.200 0.595 0.290 ;
        RECT  0.490 0.970 0.595 1.060 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.225 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  1.515 0.665 2.675 0.735 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.275 ;
        RECT  0.390 -0.115 0.990 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.210 -0.115 0.310 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.145 2.800 1.375 ;
        RECT  2.440 0.835 2.510 1.375 ;
        RECT  2.400 0.835 2.440 0.935 ;
        RECT  1.110 1.145 2.440 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.200 1.145 0.990 1.375 ;
        RECT  0.200 0.850 0.410 0.920 ;
        RECT  0.100 0.850 0.200 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.705 0.355 2.765 1.070 ;
        RECT  2.695 0.190 2.705 1.070 ;
        RECT  2.600 0.190 2.695 0.425 ;
        RECT  2.600 0.970 2.695 1.070 ;
        RECT  2.535 0.495 2.625 0.765 ;
        RECT  1.925 0.355 2.600 0.425 ;
        RECT  2.065 0.545 2.370 0.615 ;
        RECT  1.890 0.200 2.310 0.275 ;
        RECT  2.200 0.775 2.300 1.075 ;
        RECT  1.995 0.545 2.065 1.055 ;
        RECT  1.890 0.985 1.995 1.055 ;
        RECT  1.855 0.355 1.925 0.660 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.555 0.495 1.645 0.765 ;
        RECT  1.375 0.200 1.610 0.275 ;
        RECT  1.500 0.845 1.600 1.075 ;
        RECT  1.305 0.200 1.375 1.055 ;
        RECT  1.190 0.200 1.305 0.275 ;
        RECT  1.190 0.985 1.305 1.055 ;
        RECT  0.965 0.355 1.035 0.640 ;
        RECT  0.755 0.520 0.965 0.640 ;
        RECT  0.190 0.520 0.525 0.640 ;
        RECT  0.120 0.355 0.190 0.640 ;
        LAYER VIA1 ;
        RECT  2.555 0.665 2.625 0.735 ;
        RECT  2.220 0.945 2.290 1.015 ;
        RECT  1.995 0.805 2.065 0.875 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.565 0.665 1.635 0.735 ;
        RECT  1.515 0.945 1.585 1.015 ;
        RECT  1.305 0.805 1.375 0.875 ;
        RECT  0.965 0.385 1.035 0.455 ;
        RECT  0.120 0.385 0.190 0.455 ;
        LAYER M2 ;
        RECT  1.465 0.945 2.340 1.015 ;
        RECT  1.255 0.805 2.115 0.875 ;
        RECT  0.070 0.385 1.835 0.455 ;
    END
END GXNR2D2BWP40

MACRO GXOR2D1BWP40
    CLASS CORE ;
    FOREIGN GXOR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.205 0.210 0.275 ;
        RECT  0.105 0.970 0.200 1.070 ;
        RECT  0.035 0.205 0.105 1.070 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.495 0.550 0.625 ;
        RECT  0.315 0.495 0.390 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.385 1.925 0.640 ;
        RECT  1.225 0.385 1.855 0.455 ;
        RECT  1.155 0.385 1.225 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.810 -0.115 2.100 0.115 ;
        RECT  1.690 -0.115 1.810 0.270 ;
        RECT  0.410 -0.115 1.690 0.115 ;
        RECT  0.290 -0.115 0.410 0.270 ;
        RECT  0.000 -0.115 0.290 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 1.145 2.100 1.375 ;
        RECT  1.715 0.805 1.785 1.375 ;
        RECT  0.410 1.145 1.715 1.375 ;
        RECT  0.290 0.855 0.410 1.375 ;
        RECT  0.000 1.145 0.290 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.205 2.065 0.880 ;
        RECT  1.995 0.205 2.000 1.070 ;
        RECT  1.890 0.205 1.995 0.275 ;
        RECT  1.890 0.800 1.995 1.070 ;
        RECT  1.440 0.545 1.670 0.615 ;
        RECT  1.190 0.200 1.610 0.275 ;
        RECT  1.510 0.855 1.610 1.075 ;
        RECT  1.360 0.545 1.440 1.055 ;
        RECT  1.190 0.985 1.360 1.055 ;
        RECT  1.085 0.190 1.100 0.290 ;
        RECT  1.015 0.190 1.085 0.965 ;
        RECT  1.000 0.190 1.015 0.290 ;
        RECT  0.875 0.495 0.945 0.875 ;
        RECT  0.735 0.200 0.910 0.275 ;
        RECT  0.665 0.945 0.910 1.055 ;
        RECT  0.815 0.805 0.875 0.875 ;
        RECT  0.665 0.200 0.735 0.875 ;
        RECT  0.490 0.200 0.665 0.275 ;
        RECT  0.590 0.805 0.665 0.875 ;
        RECT  0.500 0.805 0.590 1.075 ;
        RECT  0.175 0.355 0.245 0.675 ;
        LAYER VIA1 ;
        RECT  1.925 0.805 1.995 0.875 ;
        RECT  1.525 0.945 1.595 1.015 ;
        RECT  1.365 0.665 1.435 0.735 ;
        RECT  1.015 0.385 1.085 0.455 ;
        RECT  0.845 0.805 0.915 0.875 ;
        RECT  0.695 0.945 0.765 1.015 ;
        RECT  0.665 0.665 0.735 0.735 ;
        RECT  0.175 0.385 0.245 0.455 ;
        LAYER M2 ;
        RECT  0.795 0.805 2.045 0.875 ;
        RECT  0.645 0.945 1.655 1.015 ;
        RECT  0.615 0.665 1.485 0.735 ;
        RECT  0.125 0.385 1.135 0.455 ;
    END
END GXOR2D1BWP40

MACRO GXOR2D2BWP40
    CLASS CORE ;
    FOREIGN GXOR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE gacore ;
    PIN Z
        ANTENNADIFFAREA 0.280000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.205 0.910 0.275 ;
        RECT  0.665 0.970 0.910 1.060 ;
        RECT  0.595 0.205 0.665 1.060 ;
        RECT  0.490 0.205 0.595 0.275 ;
        RECT  0.490 0.970 0.595 1.060 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.495 1.250 0.625 ;
        RECT  1.015 0.495 1.095 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.385 2.625 0.640 ;
        RECT  1.925 0.385 2.555 0.455 ;
        RECT  1.855 0.385 1.925 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.510 -0.115 2.800 0.115 ;
        RECT  2.390 -0.115 2.510 0.270 ;
        RECT  1.110 -0.115 2.390 0.115 ;
        RECT  0.990 -0.115 1.110 0.270 ;
        RECT  0.390 -0.115 0.990 0.115 ;
        RECT  0.310 -0.115 0.390 0.320 ;
        RECT  0.210 -0.115 0.310 0.115 ;
        RECT  0.090 -0.115 0.210 0.275 ;
        RECT  0.000 -0.115 0.090 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.485 1.145 2.800 1.375 ;
        RECT  2.415 0.805 2.485 1.375 ;
        RECT  1.110 1.145 2.415 1.375 ;
        RECT  0.990 0.855 1.110 1.375 ;
        RECT  0.200 1.145 0.990 1.375 ;
        RECT  0.200 0.850 0.410 0.920 ;
        RECT  0.100 0.850 0.200 1.375 ;
        RECT  0.000 1.145 0.100 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.700 0.205 2.765 0.880 ;
        RECT  2.695 0.205 2.700 1.070 ;
        RECT  2.590 0.205 2.695 0.275 ;
        RECT  2.590 0.800 2.695 1.070 ;
        RECT  2.140 0.545 2.370 0.615 ;
        RECT  1.890 0.200 2.310 0.275 ;
        RECT  2.210 0.855 2.310 1.075 ;
        RECT  2.060 0.545 2.140 1.055 ;
        RECT  1.890 0.985 2.060 1.055 ;
        RECT  1.785 0.190 1.800 0.290 ;
        RECT  1.715 0.190 1.785 0.965 ;
        RECT  1.700 0.190 1.715 0.290 ;
        RECT  1.575 0.495 1.645 0.875 ;
        RECT  1.435 0.200 1.610 0.275 ;
        RECT  1.365 0.945 1.610 1.055 ;
        RECT  1.515 0.805 1.575 0.875 ;
        RECT  1.365 0.200 1.435 0.875 ;
        RECT  1.190 0.200 1.365 0.275 ;
        RECT  1.290 0.805 1.365 0.875 ;
        RECT  1.200 0.805 1.290 1.075 ;
        RECT  0.875 0.355 0.945 0.660 ;
        RECT  0.765 0.510 0.875 0.660 ;
        RECT  0.180 0.520 0.525 0.640 ;
        RECT  0.035 0.355 0.180 0.640 ;
        LAYER VIA1 ;
        RECT  2.625 0.805 2.695 0.875 ;
        RECT  2.225 0.945 2.295 1.015 ;
        RECT  2.065 0.665 2.135 0.735 ;
        RECT  1.715 0.385 1.785 0.455 ;
        RECT  1.545 0.805 1.615 0.875 ;
        RECT  1.395 0.945 1.465 1.015 ;
        RECT  1.365 0.665 1.435 0.735 ;
        RECT  0.875 0.385 0.945 0.455 ;
        RECT  0.110 0.385 0.180 0.455 ;
        LAYER M2 ;
        RECT  1.495 0.805 2.745 0.875 ;
        RECT  1.345 0.945 2.355 1.015 ;
        RECT  1.315 0.665 2.185 0.735 ;
        RECT  0.060 0.385 1.835 0.455 ;
    END
END GXOR2D2BWP40

MACRO HA1D0BWP40
    CLASS CORE ;
    FOREIGN HA1D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.054000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.340 2.625 0.905 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.725 0.125 1.065 ;
        RECT  0.035 0.185 0.105 1.065 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.995 2.180 1.075 ;
        RECT  0.945 0.995 2.040 1.065 ;
        RECT  0.850 0.870 0.945 1.065 ;
        RECT  0.665 0.870 0.850 0.940 ;
        RECT  0.595 0.545 0.665 0.940 ;
        RECT  0.350 0.545 0.595 0.615 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.525 0.945 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.390 -0.115 2.660 0.115 ;
        RECT  2.270 -0.115 2.390 0.140 ;
        RECT  1.320 -0.115 2.270 0.115 ;
        RECT  1.240 -0.115 1.320 0.265 ;
        RECT  0.910 -0.115 1.240 0.115 ;
        RECT  0.820 -0.115 0.910 0.270 ;
        RECT  0.345 -0.115 0.820 0.115 ;
        RECT  0.225 -0.115 0.345 0.255 ;
        RECT  0.000 -0.115 0.225 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.145 2.660 1.375 ;
        RECT  2.290 0.735 2.370 1.375 ;
        RECT  1.250 1.145 2.290 1.375 ;
        RECT  1.140 1.135 1.250 1.375 ;
        RECT  0.770 1.145 1.140 1.375 ;
        RECT  0.650 1.010 0.770 1.375 ;
        RECT  0.350 1.145 0.650 1.375 ;
        RECT  0.230 0.940 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.520 2.460 0.640 ;
        RECT  2.320 0.210 2.390 0.640 ;
        RECT  1.695 0.210 2.320 0.280 ;
        RECT  2.075 0.350 2.145 0.860 ;
        RECT  1.930 0.520 2.075 0.600 ;
        RECT  1.860 0.855 1.950 0.925 ;
        RECT  1.860 0.350 1.930 0.420 ;
        RECT  1.780 0.350 1.860 0.925 ;
        RECT  1.260 0.855 1.780 0.925 ;
        RECT  1.620 0.210 1.695 0.785 ;
        RECT  1.460 0.195 1.530 0.785 ;
        RECT  1.435 0.195 1.460 0.315 ;
        RECT  1.370 0.715 1.460 0.785 ;
        RECT  1.260 0.510 1.390 0.630 ;
        RECT  1.190 0.365 1.260 0.925 ;
        RECT  1.095 0.365 1.190 0.455 ;
        RECT  0.935 0.730 1.190 0.800 ;
        RECT  1.005 0.185 1.095 0.455 ;
        RECT  0.560 0.205 0.740 0.275 ;
        RECT  0.490 0.205 0.560 0.415 ;
        RECT  0.455 0.710 0.525 1.060 ;
        RECT  0.275 0.345 0.490 0.415 ;
        RECT  0.275 0.710 0.455 0.780 ;
        RECT  0.195 0.345 0.275 0.780 ;
        RECT  0.180 0.520 0.195 0.640 ;
    END
END HA1D0BWP40

MACRO HA1D1BWP40
    CLASS CORE ;
    FOREIGN HA1D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.106650 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.185 2.625 1.065 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.185 0.125 0.465 ;
        RECT  0.105 0.725 0.125 1.045 ;
        RECT  0.035 0.185 0.105 1.045 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.995 2.180 1.075 ;
        RECT  0.945 0.995 2.040 1.065 ;
        RECT  0.875 0.870 0.945 1.065 ;
        RECT  0.665 0.870 0.875 0.940 ;
        RECT  0.595 0.545 0.665 0.940 ;
        RECT  0.350 0.545 0.595 0.615 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.525 0.945 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.390 -0.115 2.660 0.115 ;
        RECT  2.270 -0.115 2.390 0.140 ;
        RECT  1.320 -0.115 2.270 0.115 ;
        RECT  1.240 -0.115 1.320 0.265 ;
        RECT  0.910 -0.115 1.240 0.115 ;
        RECT  0.820 -0.115 0.910 0.270 ;
        RECT  0.345 -0.115 0.820 0.115 ;
        RECT  0.225 -0.115 0.345 0.275 ;
        RECT  0.000 -0.115 0.225 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 1.145 2.660 1.375 ;
        RECT  2.315 0.710 2.395 1.375 ;
        RECT  1.250 1.145 2.315 1.375 ;
        RECT  1.140 1.135 1.250 1.375 ;
        RECT  0.770 1.145 1.140 1.375 ;
        RECT  0.650 1.010 0.770 1.375 ;
        RECT  0.330 1.145 0.650 1.375 ;
        RECT  0.250 0.845 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.520 2.460 0.640 ;
        RECT  2.320 0.210 2.390 0.640 ;
        RECT  1.695 0.210 2.320 0.280 ;
        RECT  2.075 0.350 2.145 0.860 ;
        RECT  1.930 0.520 2.075 0.600 ;
        RECT  1.860 0.855 1.950 0.925 ;
        RECT  1.860 0.350 1.930 0.420 ;
        RECT  1.780 0.350 1.860 0.925 ;
        RECT  1.260 0.855 1.780 0.925 ;
        RECT  1.620 0.210 1.695 0.785 ;
        RECT  1.460 0.215 1.530 0.785 ;
        RECT  1.435 0.215 1.460 0.335 ;
        RECT  1.370 0.715 1.460 0.785 ;
        RECT  1.260 0.510 1.390 0.630 ;
        RECT  1.190 0.365 1.260 0.925 ;
        RECT  1.095 0.365 1.190 0.455 ;
        RECT  0.935 0.730 1.190 0.800 ;
        RECT  1.005 0.185 1.095 0.455 ;
        RECT  0.560 0.205 0.740 0.275 ;
        RECT  0.490 0.205 0.560 0.415 ;
        RECT  0.455 0.695 0.525 1.060 ;
        RECT  0.275 0.345 0.490 0.415 ;
        RECT  0.275 0.695 0.455 0.765 ;
        RECT  0.195 0.345 0.275 0.765 ;
        RECT  0.180 0.520 0.195 0.640 ;
    END
END HA1D1BWP40

MACRO HA1D2BWP40
    CLASS CORE ;
    FOREIGN HA1D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.118500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.400 0.385 3.465 0.790 ;
        RECT  3.375 0.195 3.400 1.065 ;
        RECT  3.315 0.195 3.375 0.460 ;
        RECT  3.320 0.720 3.375 1.065 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.144000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.210 0.405 0.465 ;
        RECT  0.385 0.725 0.405 1.045 ;
        RECT  0.315 0.210 0.385 1.045 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.995 3.020 1.075 ;
        RECT  1.785 0.995 2.880 1.065 ;
        RECT  1.715 0.870 1.785 1.065 ;
        RECT  1.505 0.870 1.715 0.940 ;
        RECT  1.435 0.545 1.505 0.940 ;
        RECT  0.685 0.545 1.435 0.615 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.525 1.785 0.625 ;
        RECT  1.575 0.355 1.645 0.625 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 -0.115 3.640 0.115 ;
        RECT  3.515 -0.115 3.585 0.280 ;
        RECT  3.230 -0.115 3.515 0.115 ;
        RECT  3.105 -0.115 3.230 0.140 ;
        RECT  2.160 -0.115 3.105 0.115 ;
        RECT  2.080 -0.115 2.160 0.400 ;
        RECT  1.750 -0.115 2.080 0.115 ;
        RECT  1.660 -0.115 1.750 0.270 ;
        RECT  1.055 -0.115 1.660 0.115 ;
        RECT  0.925 -0.115 1.055 0.125 ;
        RECT  0.595 -0.115 0.925 0.115 ;
        RECT  0.520 -0.115 0.595 0.255 ;
        RECT  0.155 -0.115 0.520 0.115 ;
        RECT  0.060 -0.115 0.155 0.420 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 1.145 3.640 1.375 ;
        RECT  3.515 0.865 3.585 1.375 ;
        RECT  3.210 1.145 3.515 1.375 ;
        RECT  3.130 0.710 3.210 1.375 ;
        RECT  2.090 1.145 3.130 1.375 ;
        RECT  1.980 1.135 2.090 1.375 ;
        RECT  1.610 1.145 1.980 1.375 ;
        RECT  1.490 1.010 1.610 1.375 ;
        RECT  1.160 1.145 1.490 1.375 ;
        RECT  1.085 0.975 1.160 1.375 ;
        RECT  0.985 1.145 1.085 1.375 ;
        RECT  0.910 0.975 0.985 1.375 ;
        RECT  0.600 1.145 0.910 1.375 ;
        RECT  0.520 0.865 0.600 1.375 ;
        RECT  0.150 1.145 0.520 1.375 ;
        RECT  0.060 0.720 0.150 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.540 3.300 0.620 ;
        RECT  3.160 0.210 3.230 0.620 ;
        RECT  2.535 0.210 3.160 0.280 ;
        RECT  2.915 0.350 2.985 0.860 ;
        RECT  2.770 0.520 2.915 0.600 ;
        RECT  2.700 0.855 2.790 0.925 ;
        RECT  2.700 0.350 2.770 0.420 ;
        RECT  2.620 0.350 2.700 0.925 ;
        RECT  1.935 0.855 2.620 0.925 ;
        RECT  2.460 0.210 2.535 0.785 ;
        RECT  2.300 0.215 2.370 0.785 ;
        RECT  2.275 0.215 2.300 0.335 ;
        RECT  2.210 0.715 2.300 0.785 ;
        RECT  1.935 0.510 2.230 0.630 ;
        RECT  1.865 0.185 1.935 0.925 ;
        RECT  1.775 0.730 1.865 0.800 ;
        RECT  1.505 0.205 1.580 0.275 ;
        RECT  1.435 0.205 1.505 0.455 ;
        RECT  0.555 0.385 1.435 0.455 ;
        RECT  0.690 0.210 1.365 0.310 ;
        RECT  1.290 0.820 1.360 1.055 ;
        RECT  0.805 0.820 1.290 0.895 ;
        RECT  0.785 0.710 0.805 0.895 ;
        RECT  0.715 0.710 0.785 1.060 ;
        RECT  0.555 0.710 0.715 0.780 ;
        RECT  0.475 0.385 0.555 0.780 ;
        RECT  0.460 0.520 0.475 0.640 ;
    END
END HA1D2BWP40

MACRO HA1D4BWP40
    CLASS CORE ;
    FOREIGN HA1D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN S
        ANTENNADIFFAREA 0.237000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.145 0.765 5.235 1.035 ;
        RECT  5.135 0.195 5.215 0.450 ;
        RECT  5.075 0.765 5.145 0.845 ;
        RECT  5.075 0.355 5.135 0.450 ;
        RECT  4.865 0.355 5.075 0.845 ;
        RECT  4.795 0.355 4.865 0.450 ;
        RECT  4.820 0.755 4.865 0.845 ;
        RECT  4.720 0.755 4.820 1.035 ;
        RECT  4.715 0.195 4.795 0.450 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.215 0.735 0.305 ;
        RECT  0.600 0.725 0.700 1.025 ;
        RECT  0.595 0.215 0.665 0.485 ;
        RECT  0.595 0.725 0.600 0.875 ;
        RECT  0.385 0.325 0.595 0.875 ;
        RECT  0.330 0.325 0.385 0.445 ;
        RECT  0.335 0.720 0.385 0.875 ;
        RECT  0.225 0.720 0.335 1.040 ;
        RECT  0.240 0.195 0.330 0.445 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.280 0.995 4.420 1.075 ;
        RECT  2.920 0.995 4.280 1.065 ;
        RECT  2.835 0.875 2.920 1.065 ;
        RECT  2.640 0.875 2.835 0.945 ;
        RECT  2.570 0.635 2.640 0.945 ;
        RECT  2.485 0.635 2.570 0.765 ;
        RECT  2.415 0.545 2.485 0.765 ;
        RECT  1.025 0.545 2.415 0.615 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 2.905 0.630 ;
        RECT  2.720 0.530 2.835 0.630 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.405 -0.115 5.460 0.115 ;
        RECT  5.330 -0.115 5.405 0.455 ;
        RECT  4.985 -0.115 5.330 0.115 ;
        RECT  4.915 -0.115 4.985 0.280 ;
        RECT  4.630 -0.115 4.915 0.115 ;
        RECT  4.505 -0.115 4.630 0.140 ;
        RECT  3.540 -0.115 4.505 0.115 ;
        RECT  3.415 -0.115 3.540 0.305 ;
        RECT  2.885 -0.115 3.415 0.115 ;
        RECT  2.795 -0.115 2.885 0.270 ;
        RECT  1.670 -0.115 2.795 0.115 ;
        RECT  1.560 -0.115 1.670 0.170 ;
        RECT  1.295 -0.115 1.560 0.115 ;
        RECT  1.175 -0.115 1.295 0.170 ;
        RECT  0.890 -0.115 1.175 0.115 ;
        RECT  0.815 -0.115 0.890 0.260 ;
        RECT  0.515 -0.115 0.815 0.115 ;
        RECT  0.435 -0.115 0.515 0.245 ;
        RECT  0.140 -0.115 0.435 0.115 ;
        RECT  0.045 -0.115 0.140 0.445 ;
        RECT  0.000 -0.115 0.045 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.410 1.145 5.460 1.375 ;
        RECT  5.330 0.720 5.410 1.375 ;
        RECT  5.010 1.145 5.330 1.375 ;
        RECT  4.915 0.940 5.010 1.375 ;
        RECT  4.610 1.145 4.915 1.375 ;
        RECT  4.530 0.710 4.610 1.375 ;
        RECT  3.490 1.145 4.530 1.375 ;
        RECT  3.380 1.135 3.490 1.375 ;
        RECT  2.745 1.145 3.380 1.375 ;
        RECT  2.625 1.015 2.745 1.375 ;
        RECT  2.330 1.145 2.625 1.375 ;
        RECT  2.210 1.045 2.330 1.375 ;
        RECT  1.845 1.145 2.210 1.375 ;
        RECT  1.770 0.975 1.845 1.375 ;
        RECT  1.655 1.145 1.770 1.375 ;
        RECT  1.575 0.975 1.655 1.375 ;
        RECT  1.280 1.145 1.575 1.375 ;
        RECT  1.205 0.975 1.280 1.375 ;
        RECT  0.895 1.145 1.205 1.375 ;
        RECT  0.805 0.860 0.895 1.375 ;
        RECT  0.520 1.145 0.805 1.375 ;
        RECT  0.435 1.000 0.520 1.375 ;
        RECT  0.135 1.145 0.435 1.375 ;
        RECT  0.045 0.720 0.135 1.375 ;
        RECT  0.000 1.145 0.045 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.145 0.765 5.235 1.035 ;
        RECT  5.145 0.195 5.215 0.450 ;
        RECT  4.715 0.195 4.795 0.450 ;
        RECT  4.720 0.755 4.795 1.035 ;
        RECT  0.665 0.215 0.735 0.305 ;
        RECT  0.665 0.725 0.700 1.025 ;
        RECT  0.240 0.195 0.315 0.445 ;
        RECT  0.225 0.720 0.315 1.040 ;
        RECT  4.630 0.535 4.700 0.630 ;
        RECT  4.560 0.210 4.630 0.630 ;
        RECT  3.935 0.210 4.560 0.280 ;
        RECT  4.315 0.350 4.385 0.860 ;
        RECT  4.170 0.520 4.315 0.600 ;
        RECT  4.100 0.855 4.190 0.925 ;
        RECT  4.100 0.350 4.170 0.420 ;
        RECT  4.020 0.350 4.100 0.925 ;
        RECT  3.075 0.855 4.020 0.925 ;
        RECT  3.860 0.210 3.935 0.785 ;
        RECT  3.700 0.215 3.770 0.785 ;
        RECT  3.675 0.215 3.700 0.460 ;
        RECT  3.155 0.715 3.700 0.785 ;
        RECT  3.295 0.385 3.675 0.460 ;
        RECT  3.075 0.540 3.595 0.615 ;
        RECT  3.215 0.210 3.295 0.460 ;
        RECT  3.005 0.185 3.075 0.925 ;
        RECT  2.890 0.710 3.005 0.800 ;
        RECT  2.610 0.245 2.705 0.455 ;
        RECT  0.850 0.385 2.610 0.455 ;
        RECT  0.985 0.240 2.520 0.310 ;
        RECT  2.425 0.895 2.495 1.025 ;
        RECT  2.110 0.895 2.425 0.965 ;
        RECT  2.025 0.820 2.110 1.045 ;
        RECT  1.460 0.820 2.025 0.895 ;
        RECT  1.390 0.820 1.460 1.070 ;
        RECT  1.100 0.820 1.390 0.895 ;
        RECT  1.080 0.710 1.100 0.895 ;
        RECT  1.010 0.710 1.080 1.065 ;
        RECT  0.850 0.710 1.010 0.780 ;
        RECT  0.770 0.385 0.850 0.780 ;
        RECT  0.735 0.530 0.770 0.640 ;
    END
END HA1D4BWP40

MACRO IAO21D0BWP40
    CLASS CORE ;
    FOREIGN IAO21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.054375 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 1.075 ;
        RECT  0.725 0.355 0.875 0.425 ;
        RECT  0.830 0.975 0.875 1.075 ;
        RECT  0.655 0.185 0.725 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.635 0.805 0.905 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.420 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.545 0.225 0.625 ;
        RECT  0.035 0.355 0.115 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.920 0.280 ;
        RECT  0.550 -0.115 0.840 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.060 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.980 1.375 ;
        RECT  0.430 1.000 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.515 0.345 0.585 0.915 ;
        RECT  0.330 0.345 0.515 0.415 ;
        RECT  0.140 0.845 0.515 0.915 ;
        RECT  0.250 0.185 0.330 0.415 ;
        RECT  0.060 0.845 0.140 1.055 ;
    END
END IAO21D0BWP40

MACRO IAO21D1BWP40
    CLASS CORE ;
    FOREIGN IAO21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.108750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 1.075 ;
        RECT  0.725 0.355 0.875 0.425 ;
        RECT  0.830 0.835 0.875 1.075 ;
        RECT  0.655 0.245 0.725 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.420 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.545 0.225 0.625 ;
        RECT  0.035 0.355 0.115 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.920 0.280 ;
        RECT  0.550 -0.115 0.840 0.115 ;
        RECT  0.430 -0.115 0.550 0.255 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.060 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.980 1.375 ;
        RECT  0.430 1.000 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.515 0.345 0.585 0.915 ;
        RECT  0.330 0.345 0.515 0.415 ;
        RECT  0.140 0.845 0.515 0.915 ;
        RECT  0.250 0.185 0.330 0.415 ;
        RECT  0.060 0.845 0.140 1.055 ;
    END
END IAO21D1BWP40

MACRO IAO21D2BWP40
    CLASS CORE ;
    FOREIGN IAO21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.200500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.185 1.150 0.425 ;
        RECT  0.805 0.355 1.050 0.425 ;
        RECT  0.805 0.705 0.945 0.805 ;
        RECT  0.735 0.355 0.805 0.805 ;
        RECT  0.635 0.185 0.735 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.875 0.495 1.015 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.495 0.390 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.215 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.425 ;
        RECT  0.955 -0.115 1.270 0.115 ;
        RECT  0.835 -0.115 0.955 0.215 ;
        RECT  0.530 -0.115 0.835 0.115 ;
        RECT  0.410 -0.115 0.530 0.215 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.365 1.145 1.400 1.375 ;
        RECT  1.255 1.025 1.365 1.375 ;
        RECT  0.525 1.145 1.255 1.375 ;
        RECT  0.410 1.030 0.525 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.195 0.520 1.265 0.950 ;
        RECT  0.545 0.880 1.195 0.950 ;
        RECT  0.545 0.545 0.635 0.615 ;
        RECT  0.475 0.355 0.545 0.950 ;
        RECT  0.330 0.355 0.475 0.425 ;
        RECT  0.130 0.880 0.475 0.950 ;
        RECT  0.230 0.185 0.330 0.425 ;
        RECT  0.050 0.790 0.130 1.040 ;
    END
END IAO21D2BWP40

MACRO IAO21D4BWP40
    CLASS CORE ;
    FOREIGN IAO21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.345000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.455 0.425 ;
        RECT  2.415 0.775 2.455 0.905 ;
        RECT  2.340 0.185 2.415 0.905 ;
        RECT  2.205 0.355 2.340 0.905 ;
        RECT  2.040 0.355 2.205 0.425 ;
        RECT  1.965 0.775 2.205 0.905 ;
        RECT  1.960 0.195 2.040 0.425 ;
        RECT  1.660 0.355 1.960 0.425 ;
        RECT  1.580 0.195 1.660 0.425 ;
        RECT  1.280 0.355 1.580 0.425 ;
        RECT  1.200 0.265 1.280 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.495 2.105 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.255 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.545 0.650 0.615 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.605 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.605 0.465 ;
        RECT  2.230 -0.115 2.530 0.115 ;
        RECT  2.150 -0.115 2.230 0.285 ;
        RECT  1.850 -0.115 2.150 0.115 ;
        RECT  1.770 -0.115 1.850 0.285 ;
        RECT  1.470 -0.115 1.770 0.115 ;
        RECT  1.390 -0.115 1.470 0.285 ;
        RECT  1.090 -0.115 1.390 0.115 ;
        RECT  1.015 -0.115 1.090 0.465 ;
        RECT  0.710 -0.115 1.015 0.115 ;
        RECT  0.610 -0.115 0.710 0.255 ;
        RECT  0.330 -0.115 0.610 0.115 ;
        RECT  0.230 -0.115 0.330 0.255 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.655 1.145 2.660 1.375 ;
        RECT  1.585 0.835 1.655 1.375 ;
        RECT  1.275 1.145 1.585 1.375 ;
        RECT  1.205 0.835 1.275 1.375 ;
        RECT  0.345 1.145 1.205 1.375 ;
        RECT  0.215 1.040 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.040 0.355 2.135 0.425 ;
        RECT  1.965 0.775 2.135 0.905 ;
        RECT  1.960 0.195 2.040 0.425 ;
        RECT  1.660 0.355 1.960 0.425 ;
        RECT  1.580 0.195 1.660 0.425 ;
        RECT  1.280 0.355 1.580 0.425 ;
        RECT  1.200 0.265 1.280 0.425 ;
        RECT  2.535 0.740 2.605 1.055 ;
        RECT  1.845 0.985 2.535 1.055 ;
        RECT  1.775 0.695 1.845 1.055 ;
        RECT  1.465 0.695 1.775 0.765 ;
        RECT  0.885 0.545 1.680 0.615 ;
        RECT  1.395 0.695 1.465 1.030 ;
        RECT  1.085 0.695 1.395 0.765 ;
        RECT  1.015 0.695 1.085 1.030 ;
        RECT  0.035 0.890 0.910 0.970 ;
        RECT  0.815 0.185 0.885 0.805 ;
        RECT  0.505 0.335 0.815 0.415 ;
        RECT  0.605 0.735 0.815 0.805 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.125 0.335 0.435 0.415 ;
        RECT  0.035 0.185 0.125 0.415 ;
    END
END IAO21D4BWP40

MACRO IAO22D0BWP40
    CLASS CORE ;
    FOREIGN IAO22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.064375 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.210 0.945 0.415 ;
        RECT  0.805 0.345 0.830 0.415 ;
        RECT  0.715 0.345 0.805 0.800 ;
        RECT  0.685 0.725 0.715 0.800 ;
        RECT  0.615 0.725 0.685 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.525 1.270 0.635 ;
        RECT  1.155 0.355 1.225 0.635 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.495 1.085 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.215 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.635 0.390 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.350 0.275 ;
        RECT  0.690 -0.115 1.270 0.115 ;
        RECT  0.610 -0.115 0.690 0.275 ;
        RECT  0.510 -0.115 0.610 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.145 1.400 1.375 ;
        RECT  1.040 1.045 1.160 1.375 ;
        RECT  0.130 1.145 1.040 1.375 ;
        RECT  0.050 0.995 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.905 1.345 1.025 ;
        RECT  0.800 0.905 1.275 0.975 ;
        RECT  0.545 0.525 0.590 0.635 ;
        RECT  0.475 0.345 0.545 1.050 ;
        RECT  0.320 0.345 0.475 0.415 ;
        RECT  0.410 0.980 0.475 1.050 ;
        RECT  0.240 0.185 0.320 0.415 ;
    END
END IAO22D0BWP40

MACRO IAO22D1BWP40
    CLASS CORE ;
    FOREIGN IAO22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.128750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.185 0.945 0.435 ;
        RECT  0.805 0.355 0.865 0.435 ;
        RECT  0.735 0.355 0.805 0.775 ;
        RECT  0.685 0.700 0.735 0.775 ;
        RECT  0.615 0.700 0.685 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.270 0.635 ;
        RECT  1.155 0.495 1.225 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.635 ;
        RECT  0.985 0.525 1.015 0.635 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.215 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.635 0.390 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.400 ;
        RECT  0.690 -0.115 1.260 0.115 ;
        RECT  0.610 -0.115 0.690 0.275 ;
        RECT  0.510 -0.115 0.610 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.275 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.145 1.400 1.375 ;
        RECT  1.040 0.985 1.160 1.375 ;
        RECT  0.130 1.145 1.040 1.375 ;
        RECT  0.050 0.995 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.845 1.345 0.965 ;
        RECT  0.895 0.845 1.275 0.915 ;
        RECT  0.805 0.845 0.895 1.075 ;
        RECT  0.545 0.540 0.615 0.620 ;
        RECT  0.475 0.345 0.545 1.050 ;
        RECT  0.320 0.345 0.475 0.415 ;
        RECT  0.410 0.980 0.475 1.050 ;
        RECT  0.240 0.185 0.320 0.415 ;
    END
END IAO22D1BWP40

MACRO IAO22D2BWP40
    CLASS CORE ;
    FOREIGN IAO22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.204450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.195 1.925 0.425 ;
        RECT  1.065 0.355 1.805 0.425 ;
        RECT  0.995 0.195 1.065 0.425 ;
        RECT  0.945 0.355 0.995 0.425 ;
        RECT  0.875 0.355 0.945 0.795 ;
        RECT  0.695 0.355 0.875 0.425 ;
        RECT  0.785 0.725 0.875 0.795 ;
        RECT  0.615 0.285 0.695 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.300 0.495 1.645 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.495 1.810 0.840 ;
        RECT  1.225 0.770 1.730 0.840 ;
        RECT  1.115 0.495 1.225 0.840 ;
        RECT  1.015 0.495 1.115 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.405 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 -0.115 1.960 0.115 ;
        RECT  1.350 -0.115 1.480 0.145 ;
        RECT  0.900 -0.115 1.350 0.115 ;
        RECT  0.780 -0.115 0.900 0.235 ;
        RECT  0.530 -0.115 0.780 0.115 ;
        RECT  0.410 -0.115 0.530 0.270 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.145 1.960 1.375 ;
        RECT  1.540 1.050 1.670 1.375 ;
        RECT  1.285 1.145 1.540 1.375 ;
        RECT  1.165 1.050 1.285 1.375 ;
        RECT  0.130 1.145 1.165 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.685 0.910 1.900 0.980 ;
        RECT  1.155 0.215 1.675 0.285 ;
        RECT  0.545 0.540 0.795 0.620 ;
        RECT  0.615 0.725 0.685 0.980 ;
        RECT  0.475 0.345 0.545 1.055 ;
        RECT  0.320 0.345 0.475 0.415 ;
        RECT  0.410 0.985 0.475 1.055 ;
        RECT  0.240 0.255 0.320 0.415 ;
    END
END IAO22D2BWP40

MACRO IAO22D4BWP40
    CLASS CORE ;
    FOREIGN IAO22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.374750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.355 2.650 0.425 ;
        RECT  1.795 0.195 1.865 0.425 ;
        RECT  1.575 0.355 1.795 0.425 ;
        RECT  1.575 0.715 1.705 0.800 ;
        RECT  1.485 0.355 1.575 0.800 ;
        RECT  1.415 0.195 1.485 0.800 ;
        RECT  1.365 0.355 1.415 0.800 ;
        RECT  1.105 0.355 1.365 0.425 ;
        RECT  1.195 0.715 1.365 0.800 ;
        RECT  1.015 0.195 1.105 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.045 0.495 3.325 0.625 ;
        RECT  2.975 0.495 3.045 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.485 0.765 ;
        RECT  2.065 0.545 2.415 0.615 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.675 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 -0.115 3.640 0.115 ;
        RECT  3.290 -0.115 3.415 0.215 ;
        RECT  3.035 -0.115 3.290 0.115 ;
        RECT  2.905 -0.115 3.035 0.215 ;
        RECT  1.705 -0.115 2.905 0.115 ;
        RECT  1.575 -0.115 1.705 0.235 ;
        RECT  1.320 -0.115 1.575 0.115 ;
        RECT  1.200 -0.115 1.320 0.235 ;
        RECT  0.735 -0.115 1.200 0.115 ;
        RECT  0.665 -0.115 0.735 0.275 ;
        RECT  0.360 -0.115 0.665 0.115 ;
        RECT  0.280 -0.115 0.360 0.275 ;
        RECT  0.000 -0.115 0.280 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.145 3.640 1.375 ;
        RECT  3.285 1.050 3.415 1.375 ;
        RECT  3.035 1.145 3.285 1.375 ;
        RECT  2.905 1.050 3.035 1.375 ;
        RECT  2.465 1.145 2.905 1.375 ;
        RECT  2.345 1.050 2.465 1.375 ;
        RECT  2.090 1.145 2.345 1.375 ;
        RECT  1.960 1.050 2.090 1.375 ;
        RECT  0.360 1.145 1.960 1.375 ;
        RECT  0.280 1.015 0.360 1.375 ;
        RECT  0.000 1.145 0.280 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.865 0.355 2.650 0.425 ;
        RECT  1.795 0.195 1.865 0.425 ;
        RECT  1.645 0.355 1.795 0.425 ;
        RECT  1.645 0.715 1.705 0.800 ;
        RECT  1.105 0.355 1.295 0.425 ;
        RECT  1.195 0.715 1.295 0.800 ;
        RECT  1.015 0.195 1.105 0.425 ;
        RECT  3.505 0.185 3.595 0.415 ;
        RECT  3.505 0.705 3.575 0.980 ;
        RECT  3.195 0.345 3.505 0.415 ;
        RECT  3.195 0.910 3.505 0.980 ;
        RECT  3.125 0.185 3.195 0.415 ;
        RECT  3.125 0.705 3.195 0.980 ;
        RECT  2.815 0.345 3.125 0.415 ;
        RECT  2.810 0.910 3.125 0.980 ;
        RECT  2.745 0.205 2.815 0.415 ;
        RECT  2.740 0.705 2.810 0.980 ;
        RECT  1.960 0.205 2.745 0.275 ;
        RECT  2.630 0.910 2.740 0.980 ;
        RECT  2.560 0.705 2.630 0.980 ;
        RECT  2.250 0.910 2.560 0.980 ;
        RECT  2.180 0.705 2.250 0.980 ;
        RECT  1.870 0.910 2.180 0.980 ;
        RECT  1.800 0.705 1.870 0.980 ;
        RECT  1.105 0.910 1.800 0.980 ;
        RECT  0.925 0.540 1.255 0.620 ;
        RECT  1.035 0.705 1.105 0.980 ;
        RECT  0.545 0.995 0.955 1.065 ;
        RECT  0.855 0.185 0.925 0.915 ;
        RECT  0.850 0.345 0.855 0.915 ;
        RECT  0.545 0.345 0.850 0.415 ;
        RECT  0.635 0.845 0.850 0.915 ;
        RECT  0.475 0.185 0.545 0.415 ;
        RECT  0.475 0.845 0.545 1.065 ;
        RECT  0.160 0.345 0.475 0.415 ;
        RECT  0.165 0.845 0.475 0.915 ;
        RECT  0.075 0.845 0.165 1.075 ;
        RECT  0.070 0.185 0.160 0.415 ;
    END
END IAO22D4BWP40

MACRO IIND4D0BWP40
    CLASS CORE ;
    FOREIGN IIND4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.092125 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.100 0.445 ;
        RECT  0.945 0.355 1.015 0.445 ;
        RECT  0.875 0.355 0.945 1.045 ;
        RECT  0.845 0.745 0.875 1.045 ;
        RECT  0.525 0.745 0.845 0.815 ;
        RECT  0.450 0.745 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.355 0.805 0.665 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.495 1.435 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.390 -0.115 1.490 0.275 ;
        RECT  0.340 -0.115 1.390 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.145 1.540 1.375 ;
        RECT  1.400 0.930 1.480 1.375 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  1.030 0.980 1.110 1.375 ;
        RECT  0.740 1.145 1.030 1.375 ;
        RECT  0.620 0.995 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.055 ;
        RECT  1.025 0.540 1.210 0.620 ;
        RECT  0.300 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.190 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END IIND4D0BWP40

MACRO IIND4D1BWP40
    CLASS CORE ;
    FOREIGN IIND4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.184250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.185 1.100 0.445 ;
        RECT  0.945 0.355 1.015 0.445 ;
        RECT  0.875 0.355 0.945 1.045 ;
        RECT  0.845 0.745 0.875 1.045 ;
        RECT  0.525 0.745 0.845 0.815 ;
        RECT  0.450 0.745 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.355 0.525 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.355 0.805 0.665 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.505 0.640 ;
        RECT  1.350 0.495 1.435 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.390 -0.115 1.490 0.275 ;
        RECT  0.340 -0.115 1.390 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.145 1.540 1.375 ;
        RECT  1.400 0.930 1.480 1.375 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  1.030 0.705 1.110 1.375 ;
        RECT  0.720 1.145 1.030 1.375 ;
        RECT  0.640 0.885 0.720 1.375 ;
        RECT  0.340 1.145 0.640 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.055 ;
        RECT  1.025 0.540 1.210 0.620 ;
        RECT  0.300 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.190 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END IIND4D1BWP40

MACRO IIND4D2BWP40
    CLASS CORE ;
    FOREIGN IIND4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.341750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.745 2.065 1.045 ;
        RECT  1.990 0.355 2.060 1.045 ;
        RECT  1.950 0.355 1.990 0.460 ;
        RECT  1.975 0.745 1.990 1.045 ;
        RECT  1.505 0.745 1.975 0.815 ;
        RECT  1.405 0.745 1.505 1.045 ;
        RECT  1.095 0.745 1.405 0.815 ;
        RECT  1.000 0.745 1.095 1.045 ;
        RECT  0.525 0.745 1.000 0.815 ;
        RECT  0.450 0.745 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.520 1.225 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 0.520 1.715 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.230 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.355 2.625 0.640 ;
        RECT  2.400 0.550 2.555 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.275 ;
        RECT  0.715 -0.115 2.520 0.115 ;
        RECT  0.605 -0.115 0.715 0.275 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.625 1.145 2.660 1.375 ;
        RECT  2.515 0.745 2.625 1.375 ;
        RECT  2.255 1.145 2.515 1.375 ;
        RECT  2.145 0.885 2.255 1.375 ;
        RECT  1.865 1.145 2.145 1.375 ;
        RECT  1.755 0.885 1.865 1.375 ;
        RECT  1.685 1.145 1.755 1.375 ;
        RECT  1.575 0.885 1.685 1.375 ;
        RECT  1.305 1.145 1.575 1.375 ;
        RECT  1.195 0.885 1.305 1.375 ;
        RECT  0.910 1.145 1.195 1.375 ;
        RECT  0.800 0.885 0.910 1.375 ;
        RECT  0.725 1.145 0.800 1.375 ;
        RECT  0.615 0.885 0.725 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.185 2.420 0.475 ;
        RECT  2.340 0.730 2.410 1.055 ;
        RECT  2.275 0.405 2.350 0.475 ;
        RECT  2.275 0.730 2.340 0.800 ;
        RECT  2.200 0.405 2.275 0.800 ;
        RECT  1.850 0.195 2.260 0.275 ;
        RECT  2.130 0.520 2.200 0.640 ;
        RECT  1.780 0.195 1.850 0.435 ;
        RECT  1.365 0.355 1.780 0.435 ;
        RECT  0.795 0.195 1.695 0.275 ;
        RECT  0.525 0.355 1.115 0.435 ;
        RECT  0.450 0.195 0.525 0.435 ;
        RECT  0.380 0.530 0.495 0.630 ;
        RECT  0.300 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.190 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
    END
END IIND4D2BWP40

MACRO IIND4D4BWP40
    CLASS CORE ;
    FOREIGN IIND4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.675000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.370 3.810 0.440 ;
        RECT  3.680 0.745 3.790 1.045 ;
        RECT  3.535 0.745 3.680 0.815 ;
        RECT  3.390 0.370 3.535 0.815 ;
        RECT  3.325 0.370 3.390 1.045 ;
        RECT  3.285 0.370 3.325 0.495 ;
        RECT  3.320 0.745 3.325 1.045 ;
        RECT  2.840 0.745 3.320 0.815 ;
        RECT  2.735 0.745 2.840 1.035 ;
        RECT  2.455 0.745 2.735 0.815 ;
        RECT  2.360 0.745 2.455 1.045 ;
        RECT  2.065 0.745 2.360 0.815 ;
        RECT  1.985 0.745 2.065 1.045 ;
        RECT  1.675 0.745 1.985 0.815 ;
        RECT  1.575 0.745 1.675 1.045 ;
        RECT  1.105 0.745 1.575 0.815 ;
        RECT  1.015 0.745 1.105 1.045 ;
        RECT  0.715 0.745 1.015 0.815 ;
        RECT  0.640 0.745 0.715 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.520 2.065 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.520 2.905 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.385 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.585 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.545 -0.115 4.620 0.115 ;
        RECT  4.445 -0.115 4.545 0.400 ;
        RECT  4.160 -0.115 4.445 0.115 ;
        RECT  4.075 -0.115 4.160 0.265 ;
        RECT  1.295 -0.115 4.075 0.115 ;
        RECT  1.185 -0.115 1.295 0.275 ;
        RECT  0.905 -0.115 1.185 0.115 ;
        RECT  0.795 -0.115 0.905 0.275 ;
        RECT  0.530 -0.115 0.795 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.140 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.145 4.620 1.375 ;
        RECT  4.455 0.720 4.535 1.375 ;
        RECT  4.160 1.145 4.455 1.375 ;
        RECT  4.075 0.925 4.160 1.375 ;
        RECT  3.970 1.145 4.075 1.375 ;
        RECT  3.900 0.855 3.970 1.375 ;
        RECT  3.610 1.145 3.900 1.375 ;
        RECT  3.490 0.905 3.610 1.375 ;
        RECT  3.195 1.145 3.490 1.375 ;
        RECT  3.115 0.915 3.195 1.375 ;
        RECT  3.015 1.145 3.115 1.375 ;
        RECT  2.920 0.915 3.015 1.375 ;
        RECT  2.655 1.145 2.920 1.375 ;
        RECT  2.535 0.905 2.655 1.375 ;
        RECT  2.270 1.145 2.535 1.375 ;
        RECT  2.150 0.905 2.270 1.375 ;
        RECT  1.890 1.145 2.150 1.375 ;
        RECT  1.770 0.905 1.890 1.375 ;
        RECT  1.475 1.145 1.770 1.375 ;
        RECT  1.395 0.945 1.475 1.375 ;
        RECT  1.295 1.145 1.395 1.375 ;
        RECT  1.205 0.945 1.295 1.375 ;
        RECT  0.920 1.145 1.205 1.375 ;
        RECT  0.800 0.905 0.920 1.375 ;
        RECT  0.530 1.145 0.800 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.050 0.720 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.370 3.810 0.440 ;
        RECT  3.680 0.745 3.790 1.045 ;
        RECT  3.605 0.745 3.680 0.815 ;
        RECT  2.840 0.745 3.255 0.815 ;
        RECT  2.735 0.745 2.840 1.035 ;
        RECT  2.455 0.745 2.735 0.815 ;
        RECT  2.360 0.745 2.455 1.045 ;
        RECT  2.065 0.745 2.360 0.815 ;
        RECT  1.985 0.745 2.065 1.045 ;
        RECT  1.675 0.745 1.985 0.815 ;
        RECT  1.575 0.745 1.675 1.045 ;
        RECT  1.105 0.745 1.575 0.815 ;
        RECT  1.015 0.745 1.105 1.045 ;
        RECT  0.715 0.745 1.015 0.815 ;
        RECT  0.640 0.745 0.715 1.045 ;
        RECT  4.265 0.230 4.335 0.425 ;
        RECT  4.265 0.735 4.335 1.055 ;
        RECT  4.100 0.355 4.265 0.425 ;
        RECT  4.100 0.735 4.265 0.805 ;
        RECT  4.030 0.355 4.100 0.805 ;
        RECT  3.665 0.540 4.030 0.620 ;
        RECT  3.195 0.195 3.995 0.275 ;
        RECT  3.125 0.195 3.195 0.425 ;
        RECT  2.335 0.345 3.125 0.425 ;
        RECT  1.375 0.195 3.040 0.275 ;
        RECT  0.715 0.345 2.080 0.425 ;
        RECT  0.640 0.195 0.715 0.425 ;
        RECT  0.570 0.530 0.685 0.630 ;
        RECT  0.490 0.345 0.570 0.915 ;
        RECT  0.320 0.345 0.490 0.415 ;
        RECT  0.320 0.845 0.490 0.915 ;
        RECT  0.240 0.190 0.320 0.415 ;
        RECT  0.240 0.845 0.320 1.045 ;
    END
END IIND4D4BWP40

MACRO IINR4D0BWP40
    CLASS CORE ;
    FOREIGN IINR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.081875 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.775 1.100 1.075 ;
        RECT  0.945 0.775 1.015 0.905 ;
        RECT  0.875 0.215 0.945 0.905 ;
        RECT  0.845 0.215 0.875 0.415 ;
        RECT  0.525 0.345 0.845 0.415 ;
        RECT  0.450 0.215 0.525 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.645 0.230 0.765 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.620 1.505 0.905 ;
        RECT  1.350 0.620 1.435 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.390 -0.115 1.490 0.305 ;
        RECT  1.125 -0.115 1.390 0.115 ;
        RECT  1.035 -0.115 1.125 0.300 ;
        RECT  0.730 -0.115 1.035 0.115 ;
        RECT  0.625 -0.115 0.730 0.230 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.145 1.540 1.375 ;
        RECT  1.400 0.990 1.480 1.375 ;
        RECT  0.340 1.145 1.400 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.075 ;
        RECT  1.025 0.540 1.210 0.620 ;
        RECT  0.300 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.070 ;
    END
END IINR4D0BWP40

MACRO IINR4D1BWP40
    CLASS CORE ;
    FOREIGN IINR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.163750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.775 1.100 1.075 ;
        RECT  0.945 0.775 1.015 0.905 ;
        RECT  0.875 0.185 0.945 0.905 ;
        RECT  0.845 0.185 0.875 0.415 ;
        RECT  0.525 0.345 0.845 0.415 ;
        RECT  0.450 0.215 0.525 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.570 0.640 ;
        RECT  0.455 0.495 0.525 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.645 0.230 0.765 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.620 1.505 0.905 ;
        RECT  1.350 0.620 1.435 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 -0.115 1.540 0.115 ;
        RECT  1.390 -0.115 1.490 0.305 ;
        RECT  1.125 -0.115 1.390 0.115 ;
        RECT  1.035 -0.115 1.125 0.460 ;
        RECT  0.730 -0.115 1.035 0.115 ;
        RECT  0.625 -0.115 0.730 0.230 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.145 1.540 1.375 ;
        RECT  1.400 0.990 1.480 1.375 ;
        RECT  0.340 1.145 1.400 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.185 1.280 1.075 ;
        RECT  1.025 0.540 1.210 0.620 ;
        RECT  0.300 0.345 0.380 0.915 ;
        RECT  0.130 0.345 0.300 0.415 ;
        RECT  0.130 0.845 0.300 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.070 ;
    END
END IINR4D1BWP40

MACRO IINR4D2BWP40
    CLASS CORE ;
    FOREIGN IINR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.294250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.185 2.065 0.905 ;
        RECT  1.975 0.185 1.990 0.415 ;
        RECT  1.950 0.800 1.990 0.905 ;
        RECT  1.505 0.345 1.975 0.415 ;
        RECT  1.405 0.185 1.505 0.415 ;
        RECT  1.085 0.345 1.405 0.415 ;
        RECT  1.015 0.185 1.085 0.415 ;
        RECT  0.525 0.345 1.015 0.415 ;
        RECT  0.450 0.205 0.525 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.090 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.510 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.230 0.665 ;
        RECT  0.035 0.435 0.105 0.790 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.520 2.625 0.905 ;
        RECT  2.440 0.520 2.555 0.610 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.400 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.160 -0.115 2.260 0.285 ;
        RECT  1.850 -0.115 2.160 0.115 ;
        RECT  1.770 -0.115 1.850 0.270 ;
        RECT  1.670 -0.115 1.770 0.115 ;
        RECT  1.590 -0.115 1.670 0.270 ;
        RECT  1.295 -0.115 1.590 0.115 ;
        RECT  1.205 -0.115 1.295 0.270 ;
        RECT  0.895 -0.115 1.205 0.115 ;
        RECT  0.815 -0.115 0.895 0.270 ;
        RECT  0.715 -0.115 0.815 0.115 ;
        RECT  0.605 -0.115 0.715 0.275 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.215 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.995 2.610 1.375 ;
        RECT  0.720 1.145 2.530 1.375 ;
        RECT  0.620 1.000 0.720 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 1.040 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.785 2.420 1.075 ;
        RECT  2.340 0.250 2.410 0.435 ;
        RECT  2.275 0.785 2.350 0.855 ;
        RECT  2.275 0.365 2.340 0.435 ;
        RECT  2.200 0.365 2.275 0.855 ;
        RECT  1.850 0.985 2.260 1.065 ;
        RECT  2.135 0.520 2.200 0.640 ;
        RECT  1.780 0.845 1.850 1.065 ;
        RECT  1.380 0.845 1.780 0.915 ;
        RECT  0.800 0.995 1.695 1.065 ;
        RECT  0.525 0.845 1.115 0.915 ;
        RECT  0.380 0.545 0.565 0.615 ;
        RECT  0.450 0.750 0.525 1.010 ;
        RECT  0.300 0.285 0.380 0.970 ;
        RECT  0.130 0.285 0.300 0.355 ;
        RECT  0.130 0.900 0.300 0.970 ;
        RECT  0.050 0.215 0.130 0.355 ;
        RECT  0.050 0.900 0.130 1.070 ;
    END
END IINR4D2BWP40

MACRO IINR4D4BWP40
    CLASS CORE ;
    FOREIGN IINR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.581000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.820 3.810 0.890 ;
        RECT  3.705 0.185 3.795 0.415 ;
        RECT  3.535 0.345 3.705 0.415 ;
        RECT  3.390 0.345 3.535 0.890 ;
        RECT  3.325 0.185 3.390 0.890 ;
        RECT  3.320 0.185 3.325 0.415 ;
        RECT  3.285 0.765 3.325 0.890 ;
        RECT  2.820 0.345 3.320 0.415 ;
        RECT  2.750 0.185 2.820 0.415 ;
        RECT  2.440 0.345 2.750 0.415 ;
        RECT  2.370 0.185 2.440 0.415 ;
        RECT  2.055 0.345 2.370 0.415 ;
        RECT  1.985 0.185 2.055 0.415 ;
        RECT  1.665 0.345 1.985 0.415 ;
        RECT  1.595 0.185 1.665 0.415 ;
        RECT  1.095 0.345 1.595 0.415 ;
        RECT  1.025 0.185 1.095 0.415 ;
        RECT  0.715 0.345 1.025 0.415 ;
        RECT  0.640 0.215 0.715 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 0.495 1.975 0.615 ;
        RECT  1.710 0.495 1.790 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.690 0.495 2.770 0.765 ;
        RECT  2.445 0.495 2.690 0.615 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.385 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.495 4.585 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.545 -0.115 4.620 0.115 ;
        RECT  4.445 -0.115 4.545 0.410 ;
        RECT  4.160 -0.115 4.445 0.115 ;
        RECT  4.075 -0.115 4.160 0.260 ;
        RECT  3.975 -0.115 4.075 0.115 ;
        RECT  3.895 -0.115 3.975 0.260 ;
        RECT  3.595 -0.115 3.895 0.115 ;
        RECT  3.495 -0.115 3.595 0.275 ;
        RECT  3.205 -0.115 3.495 0.115 ;
        RECT  3.115 -0.115 3.205 0.275 ;
        RECT  3.015 -0.115 3.115 0.115 ;
        RECT  2.935 -0.115 3.015 0.275 ;
        RECT  2.640 -0.115 2.935 0.115 ;
        RECT  2.550 -0.115 2.640 0.275 ;
        RECT  2.255 -0.115 2.550 0.115 ;
        RECT  2.175 -0.115 2.255 0.275 ;
        RECT  1.880 -0.115 2.175 0.115 ;
        RECT  1.785 -0.115 1.880 0.275 ;
        RECT  1.485 -0.115 1.785 0.115 ;
        RECT  1.395 -0.115 1.485 0.275 ;
        RECT  1.295 -0.115 1.395 0.115 ;
        RECT  1.185 -0.115 1.295 0.275 ;
        RECT  0.905 -0.115 1.185 0.115 ;
        RECT  0.795 -0.115 0.905 0.275 ;
        RECT  0.530 -0.115 0.795 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.145 4.620 1.375 ;
        RECT  4.455 0.720 4.535 1.375 ;
        RECT  4.160 1.145 4.455 1.375 ;
        RECT  4.075 0.970 4.160 1.375 ;
        RECT  1.295 1.145 4.075 1.375 ;
        RECT  1.205 0.995 1.295 1.375 ;
        RECT  0.905 1.145 1.205 1.375 ;
        RECT  0.815 1.005 0.905 1.375 ;
        RECT  0.530 1.145 0.815 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.050 0.720 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.820 3.810 0.890 ;
        RECT  3.705 0.185 3.795 0.415 ;
        RECT  3.605 0.345 3.705 0.415 ;
        RECT  2.820 0.345 3.255 0.415 ;
        RECT  2.750 0.185 2.820 0.415 ;
        RECT  2.440 0.345 2.750 0.415 ;
        RECT  2.370 0.185 2.440 0.415 ;
        RECT  2.055 0.345 2.370 0.415 ;
        RECT  1.985 0.185 2.055 0.415 ;
        RECT  1.665 0.345 1.985 0.415 ;
        RECT  1.595 0.185 1.665 0.415 ;
        RECT  1.095 0.345 1.595 0.415 ;
        RECT  1.025 0.185 1.095 0.415 ;
        RECT  0.715 0.345 1.025 0.415 ;
        RECT  0.640 0.215 0.715 0.415 ;
        RECT  4.265 0.205 4.335 0.410 ;
        RECT  4.265 0.795 4.335 1.075 ;
        RECT  4.085 0.340 4.265 0.410 ;
        RECT  4.085 0.795 4.265 0.880 ;
        RECT  4.015 0.340 4.085 0.880 ;
        RECT  3.665 0.540 4.015 0.620 ;
        RECT  3.195 0.985 3.995 1.065 ;
        RECT  3.125 0.845 3.195 1.065 ;
        RECT  2.335 0.845 3.125 0.915 ;
        RECT  1.375 0.985 3.040 1.065 ;
        RECT  1.095 0.845 2.080 0.915 ;
        RECT  0.570 0.530 1.120 0.630 ;
        RECT  1.025 0.750 1.095 1.010 ;
        RECT  0.715 0.845 1.025 0.915 ;
        RECT  0.640 0.750 0.715 1.010 ;
        RECT  0.490 0.345 0.570 0.915 ;
        RECT  0.320 0.345 0.490 0.415 ;
        RECT  0.320 0.845 0.490 0.915 ;
        RECT  0.240 0.215 0.320 0.415 ;
        RECT  0.240 0.845 0.320 1.070 ;
    END
END IINR4D4BWP40

MACRO IND2D0BWP40
    CLASS CORE ;
    FOREIGN IND2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.061750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 0.780 ;
        RECT  0.635 0.215 0.735 0.285 ;
        RECT  0.555 0.710 0.735 0.780 ;
        RECT  0.455 0.710 0.555 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.665 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.385 -0.115 0.840 0.115 ;
        RECT  0.265 -0.115 0.385 0.275 ;
        RECT  0.000 -0.115 0.265 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.145 0.840 1.375 ;
        RECT  0.655 0.985 0.755 1.375 ;
        RECT  0.375 1.145 0.655 1.375 ;
        RECT  0.275 0.985 0.375 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.385 0.545 0.465 0.615 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.175 0.345 0.315 0.415 ;
        RECT  0.175 0.845 0.315 0.915 ;
        RECT  0.100 0.185 0.175 0.415 ;
        RECT  0.100 0.845 0.175 1.070 ;
    END
END IND2D0BWP40

MACRO IND2D1BWP40
    CLASS CORE ;
    FOREIGN IND2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.123500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.215 0.805 0.780 ;
        RECT  0.635 0.215 0.735 0.285 ;
        RECT  0.555 0.710 0.735 0.780 ;
        RECT  0.455 0.710 0.555 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.355 0.665 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.385 -0.115 0.840 0.115 ;
        RECT  0.265 -0.115 0.385 0.275 ;
        RECT  0.000 -0.115 0.265 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.145 0.840 1.375 ;
        RECT  0.655 0.860 0.755 1.375 ;
        RECT  0.375 1.145 0.655 1.375 ;
        RECT  0.275 0.985 0.375 1.375 ;
        RECT  0.000 1.145 0.275 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.385 0.545 0.465 0.615 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.175 0.345 0.315 0.415 ;
        RECT  0.175 0.845 0.315 0.915 ;
        RECT  0.100 0.185 0.175 0.415 ;
        RECT  0.100 0.845 0.175 1.070 ;
    END
END IND2D1BWP40

MACRO IND2D2BWP40
    CLASS CORE ;
    FOREIGN IND2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.187500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.355 1.130 0.435 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.960 0.355 1.030 0.530 ;
        RECT  0.685 0.710 1.010 0.800 ;
        RECT  0.685 0.440 0.960 0.530 ;
        RECT  0.595 0.440 0.685 0.800 ;
        RECT  0.535 0.710 0.595 0.800 ;
        RECT  0.435 0.710 0.535 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.350 1.365 0.640 ;
        RECT  1.100 0.520 1.275 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.225 0.625 ;
        RECT  0.035 0.495 0.130 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 1.400 0.115 ;
        RECT  0.600 -0.115 0.730 0.230 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.400 1.375 ;
        RECT  1.220 0.720 1.320 1.375 ;
        RECT  0.890 1.145 1.220 1.375 ;
        RECT  0.810 0.935 0.890 1.375 ;
        RECT  0.720 1.145 0.810 1.375 ;
        RECT  0.625 0.925 0.720 1.375 ;
        RECT  0.330 1.145 0.625 1.375 ;
        RECT  0.230 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.890 0.195 1.315 0.270 ;
        RECT  0.820 0.195 0.890 0.370 ;
        RECT  0.520 0.300 0.820 0.370 ;
        RECT  0.440 0.300 0.520 0.440 ;
        RECT  0.365 0.545 0.490 0.615 ;
        RECT  0.295 0.345 0.365 0.915 ;
        RECT  0.130 0.345 0.295 0.415 ;
        RECT  0.130 0.845 0.295 0.915 ;
        RECT  0.055 0.185 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.070 ;
    END
END IND2D2BWP40

MACRO IND2D3BWP40
    CLASS CORE ;
    FOREIGN IND2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.303250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.195 1.505 0.445 ;
        RECT  1.105 0.355 1.405 0.445 ;
        RECT  1.200 0.710 1.300 1.045 ;
        RECT  1.105 0.710 1.200 0.800 ;
        RECT  1.015 0.355 1.105 0.800 ;
        RECT  0.920 0.710 1.015 0.800 ;
        RECT  0.820 0.710 0.920 1.045 ;
        RECT  0.535 0.710 0.820 0.800 ;
        RECT  0.435 0.710 0.535 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.520 1.505 0.905 ;
        RECT  1.195 0.520 1.410 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.495 0.225 0.625 ;
        RECT  0.035 0.495 0.130 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.115 1.540 0.115 ;
        RECT  0.590 -0.115 0.720 0.230 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 1.010 1.500 1.375 ;
        RECT  1.110 1.145 1.400 1.375 ;
        RECT  1.010 0.900 1.110 1.375 ;
        RECT  0.710 1.145 1.010 1.375 ;
        RECT  0.615 0.900 0.710 1.375 ;
        RECT  0.330 1.145 0.615 1.375 ;
        RECT  0.230 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.890 0.195 1.315 0.270 ;
        RECT  0.820 0.195 0.890 0.370 ;
        RECT  0.520 0.300 0.820 0.370 ;
        RECT  0.440 0.300 0.520 0.440 ;
        RECT  0.365 0.545 0.490 0.615 ;
        RECT  0.295 0.345 0.365 0.915 ;
        RECT  0.130 0.345 0.295 0.415 ;
        RECT  0.130 0.845 0.295 0.915 ;
        RECT  0.055 0.185 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.070 ;
    END
END IND2D3BWP40

MACRO IND2D4BWP40
    CLASS CORE ;
    FOREIGN IND2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.399500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.355 2.090 0.445 ;
        RECT  1.980 0.710 2.080 1.045 ;
        RECT  1.855 0.710 1.980 0.800 ;
        RECT  1.700 0.355 1.855 0.800 ;
        RECT  1.645 0.355 1.700 1.045 ;
        RECT  1.595 0.355 1.645 0.485 ;
        RECT  1.600 0.710 1.645 1.045 ;
        RECT  1.110 0.710 1.600 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
        RECT  0.625 0.710 0.725 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.520 2.345 0.905 ;
        RECT  1.980 0.520 2.250 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.415 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 2.380 0.115 ;
        RECT  1.200 -0.115 1.320 0.230 ;
        RECT  0.910 -0.115 1.200 0.115 ;
        RECT  0.780 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.780 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.135 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.135 0.410 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.145 2.380 1.375 ;
        RECT  2.240 1.010 2.340 1.375 ;
        RECT  1.890 1.145 2.240 1.375 ;
        RECT  1.790 0.985 1.890 1.375 ;
        RECT  1.510 1.145 1.790 1.375 ;
        RECT  1.410 0.985 1.510 1.375 ;
        RECT  1.300 1.145 1.410 1.375 ;
        RECT  1.205 0.965 1.300 1.375 ;
        RECT  0.900 1.145 1.205 1.375 ;
        RECT  0.805 0.925 0.900 1.375 ;
        RECT  0.520 1.145 0.805 1.375 ;
        RECT  0.420 0.985 0.520 1.375 ;
        RECT  0.135 1.145 0.420 1.375 ;
        RECT  0.050 0.860 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.625 0.710 0.725 1.045 ;
        RECT  2.240 0.195 2.315 0.450 ;
        RECT  1.480 0.195 2.240 0.270 ;
        RECT  1.410 0.195 1.480 0.370 ;
        RECT  0.710 0.300 1.410 0.370 ;
        RECT  0.555 0.545 1.115 0.615 ;
        RECT  0.630 0.300 0.710 0.440 ;
        RECT  0.485 0.345 0.555 0.915 ;
        RECT  0.320 0.345 0.485 0.415 ;
        RECT  0.320 0.845 0.485 0.915 ;
        RECT  0.245 0.185 0.320 0.415 ;
        RECT  0.245 0.845 0.320 1.070 ;
        RECT  1.925 0.355 2.090 0.445 ;
        RECT  1.980 0.710 2.080 1.045 ;
        RECT  1.925 0.710 1.980 0.800 ;
        RECT  1.110 0.710 1.575 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
    END
END IND2D4BWP40

MACRO IND2D6BWP40
    CLASS CORE ;
    FOREIGN IND2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.576000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.860 0.445 ;
        RECT  2.750 0.710 2.850 1.045 ;
        RECT  2.470 0.710 2.750 0.800 ;
        RECT  2.370 0.710 2.470 1.045 ;
        RECT  2.275 0.710 2.370 0.800 ;
        RECT  2.090 0.355 2.275 0.800 ;
        RECT  2.065 0.355 2.090 1.045 ;
        RECT  1.985 0.355 2.065 0.485 ;
        RECT  1.990 0.710 2.065 1.045 ;
        RECT  1.510 0.710 1.990 0.800 ;
        RECT  1.410 0.710 1.510 1.045 ;
        RECT  1.110 0.710 1.410 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
        RECT  0.625 0.710 0.725 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 0.520 3.045 0.905 ;
        RECT  2.370 0.520 2.950 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.415 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.115 3.080 0.115 ;
        RECT  1.600 -0.115 1.720 0.230 ;
        RECT  1.325 -0.115 1.600 0.115 ;
        RECT  1.195 -0.115 1.325 0.230 ;
        RECT  0.910 -0.115 1.195 0.115 ;
        RECT  0.780 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.780 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.135 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.135 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 1.145 3.080 1.375 ;
        RECT  2.940 1.010 3.040 1.375 ;
        RECT  2.660 1.145 2.940 1.375 ;
        RECT  2.560 0.870 2.660 1.375 ;
        RECT  2.280 1.145 2.560 1.375 ;
        RECT  2.180 0.870 2.280 1.375 ;
        RECT  1.900 1.145 2.180 1.375 ;
        RECT  1.800 0.870 1.900 1.375 ;
        RECT  1.700 1.145 1.800 1.375 ;
        RECT  1.600 0.870 1.700 1.375 ;
        RECT  1.310 1.145 1.600 1.375 ;
        RECT  1.215 0.870 1.310 1.375 ;
        RECT  0.900 1.145 1.215 1.375 ;
        RECT  0.805 0.870 0.900 1.375 ;
        RECT  0.520 1.145 0.805 1.375 ;
        RECT  0.420 0.985 0.520 1.375 ;
        RECT  0.135 1.145 0.420 1.375 ;
        RECT  0.050 0.860 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.355 2.860 0.445 ;
        RECT  2.750 0.710 2.850 1.045 ;
        RECT  2.470 0.710 2.750 0.800 ;
        RECT  2.370 0.710 2.470 1.045 ;
        RECT  2.345 0.710 2.370 0.800 ;
        RECT  1.985 0.355 1.995 0.485 ;
        RECT  1.990 0.710 1.995 1.045 ;
        RECT  1.510 0.710 1.990 0.800 ;
        RECT  1.410 0.710 1.510 1.045 ;
        RECT  1.110 0.710 1.410 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
        RECT  0.625 0.710 0.725 1.045 ;
        RECT  2.950 0.195 3.030 0.370 ;
        RECT  1.880 0.195 2.950 0.270 ;
        RECT  1.810 0.195 1.880 0.440 ;
        RECT  1.485 0.370 1.810 0.440 ;
        RECT  1.415 0.210 1.485 0.440 ;
        RECT  1.085 0.370 1.415 0.440 ;
        RECT  0.320 0.845 0.485 0.915 ;
        RECT  0.245 0.185 0.320 0.415 ;
        RECT  0.245 0.845 0.320 1.070 ;
        RECT  0.555 0.545 1.350 0.615 ;
        RECT  1.015 0.210 1.085 0.440 ;
        RECT  0.700 0.370 1.015 0.440 ;
        RECT  0.630 0.255 0.700 0.440 ;
        RECT  0.485 0.345 0.555 0.915 ;
        RECT  0.320 0.345 0.485 0.415 ;
    END
END IND2D6BWP40

MACRO IND2D8BWP40
    CLASS CORE ;
    FOREIGN IND2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.763500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.355 3.820 0.445 ;
        RECT  3.710 0.710 3.810 1.045 ;
        RECT  3.430 0.710 3.710 0.800 ;
        RECT  3.330 0.710 3.430 1.045 ;
        RECT  3.050 0.710 3.330 0.800 ;
        RECT  2.950 0.710 3.050 1.045 ;
        RECT  2.835 0.710 2.950 0.800 ;
        RECT  2.670 0.355 2.835 0.800 ;
        RECT  2.625 0.355 2.670 1.045 ;
        RECT  2.565 0.355 2.625 0.485 ;
        RECT  2.570 0.710 2.625 1.045 ;
        RECT  2.090 0.710 2.570 0.800 ;
        RECT  1.990 0.710 2.090 1.045 ;
        RECT  1.700 0.710 1.990 0.800 ;
        RECT  1.600 0.710 1.700 1.045 ;
        RECT  1.300 0.710 1.600 0.800 ;
        RECT  1.200 0.710 1.300 1.045 ;
        RECT  0.915 0.710 1.200 0.800 ;
        RECT  0.815 0.710 0.915 1.045 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 0.520 4.025 0.905 ;
        RECT  2.950 0.520 3.930 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.555 0.765 ;
        RECT  0.300 0.495 0.455 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.115 4.060 0.115 ;
        RECT  2.180 -0.115 2.300 0.230 ;
        RECT  1.905 -0.115 2.180 0.115 ;
        RECT  1.775 -0.115 1.905 0.230 ;
        RECT  1.515 -0.115 1.775 0.115 ;
        RECT  1.385 -0.115 1.515 0.230 ;
        RECT  1.100 -0.115 1.385 0.115 ;
        RECT  0.970 -0.115 1.100 0.230 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.275 ;
        RECT  0.325 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.325 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.020 1.145 4.060 1.375 ;
        RECT  3.920 1.010 4.020 1.375 ;
        RECT  3.620 1.145 3.920 1.375 ;
        RECT  3.520 0.900 3.620 1.375 ;
        RECT  3.240 1.145 3.520 1.375 ;
        RECT  3.140 0.900 3.240 1.375 ;
        RECT  2.860 1.145 3.140 1.375 ;
        RECT  2.760 0.900 2.860 1.375 ;
        RECT  2.480 1.145 2.760 1.375 ;
        RECT  2.390 0.900 2.480 1.375 ;
        RECT  2.280 1.145 2.390 1.375 ;
        RECT  2.185 0.900 2.280 1.375 ;
        RECT  1.890 1.145 2.185 1.375 ;
        RECT  1.795 0.900 1.890 1.375 ;
        RECT  1.500 1.145 1.795 1.375 ;
        RECT  1.405 0.900 1.500 1.375 ;
        RECT  1.090 1.145 1.405 1.375 ;
        RECT  0.995 0.900 1.090 1.375 ;
        RECT  0.710 1.145 0.995 1.375 ;
        RECT  0.610 0.985 0.710 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.225 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.355 3.820 0.445 ;
        RECT  3.710 0.710 3.810 1.045 ;
        RECT  3.430 0.710 3.710 0.800 ;
        RECT  3.330 0.710 3.430 1.045 ;
        RECT  3.050 0.710 3.330 0.800 ;
        RECT  2.950 0.710 3.050 1.045 ;
        RECT  2.905 0.710 2.950 0.800 ;
        RECT  2.090 0.710 2.555 0.800 ;
        RECT  1.990 0.710 2.090 1.045 ;
        RECT  1.700 0.710 1.990 0.800 ;
        RECT  1.600 0.710 1.700 1.045 ;
        RECT  1.300 0.710 1.600 0.800 ;
        RECT  1.200 0.710 1.300 1.045 ;
        RECT  0.915 0.710 1.200 0.800 ;
        RECT  0.815 0.710 0.915 1.045 ;
        RECT  3.930 0.195 4.010 0.370 ;
        RECT  2.460 0.195 3.930 0.270 ;
        RECT  2.390 0.195 2.460 0.415 ;
        RECT  2.075 0.345 2.390 0.415 ;
        RECT  0.745 0.525 2.080 0.615 ;
        RECT  2.005 0.185 2.075 0.415 ;
        RECT  1.680 0.345 2.005 0.415 ;
        RECT  1.610 0.185 1.680 0.415 ;
        RECT  1.285 0.345 1.610 0.415 ;
        RECT  1.215 0.185 1.285 0.415 ;
        RECT  0.885 0.345 1.215 0.415 ;
        RECT  0.815 0.250 0.885 0.415 ;
        RECT  0.675 0.345 0.745 0.915 ;
        RECT  0.505 0.345 0.675 0.415 ;
        RECT  0.505 0.845 0.675 0.915 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.435 0.845 0.505 1.075 ;
        RECT  0.125 0.345 0.435 0.415 ;
        RECT  0.125 0.845 0.435 0.915 ;
        RECT  0.055 0.250 0.125 0.415 ;
        RECT  0.055 0.755 0.125 1.010 ;
    END
END IND2D8BWP40

MACRO IND3D0BWP40
    CLASS CORE ;
    FOREIGN IND3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.082000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.195 0.945 0.265 ;
        RECT  0.855 0.845 0.925 1.045 ;
        RECT  0.545 0.845 0.855 0.915 ;
        RECT  0.525 0.740 0.545 1.045 ;
        RECT  0.455 0.195 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.345 0.685 0.660 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 -0.115 0.980 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 1.020 0.760 1.375 ;
        RECT  0.340 1.145 0.640 1.375 ;
        RECT  0.260 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.345 0.385 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END IND3D0BWP40

MACRO IND3D1BWP40
    CLASS CORE ;
    FOREIGN IND3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.164000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.195 0.945 0.405 ;
        RECT  0.855 0.845 0.925 1.045 ;
        RECT  0.545 0.845 0.855 0.915 ;
        RECT  0.525 0.195 0.835 0.265 ;
        RECT  0.525 0.740 0.545 1.045 ;
        RECT  0.455 0.195 0.525 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.345 0.685 0.660 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 -0.115 0.980 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.980 1.375 ;
        RECT  0.640 1.020 0.760 1.375 ;
        RECT  0.340 1.145 0.640 1.375 ;
        RECT  0.260 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.345 0.385 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END IND3D1BWP40

MACRO IND3D2BWP40
    CLASS CORE ;
    FOREIGN IND3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.287000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.845 1.505 1.075 ;
        RECT  1.365 0.345 1.500 0.415 ;
        RECT  1.365 0.845 1.405 0.925 ;
        RECT  1.295 0.345 1.365 0.925 ;
        RECT  1.105 0.845 1.295 0.925 ;
        RECT  1.015 0.845 1.105 1.075 ;
        RECT  0.535 0.845 1.015 0.925 ;
        RECT  0.445 0.760 0.535 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.645 0.630 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.090 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.115 1.820 0.115 ;
        RECT  0.620 -0.115 0.715 0.270 ;
        RECT  0.355 -0.115 0.620 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.145 1.820 1.375 ;
        RECT  1.635 0.720 1.725 1.375 ;
        RECT  1.290 1.145 1.635 1.375 ;
        RECT  1.205 0.995 1.290 1.375 ;
        RECT  0.900 1.145 1.205 1.375 ;
        RECT  0.820 0.995 0.900 1.375 ;
        RECT  0.720 1.145 0.820 1.375 ;
        RECT  0.640 0.995 0.720 1.375 ;
        RECT  0.340 1.145 0.640 1.375 ;
        RECT  0.260 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.615 0.195 1.725 0.405 ;
        RECT  0.800 0.195 1.615 0.265 ;
        RECT  0.535 0.345 1.145 0.415 ;
        RECT  0.450 0.250 0.535 0.415 ;
        RECT  0.375 0.530 0.500 0.640 ;
        RECT  0.290 0.345 0.375 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.250 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.040 ;
    END
END IND3D2BWP40

MACRO IND3D3BWP40
    CLASS CORE ;
    FOREIGN IND3D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.414500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.185 2.065 0.415 ;
        RECT  1.975 0.845 2.065 1.075 ;
        RECT  1.505 0.345 1.975 0.415 ;
        RECT  1.665 0.845 1.975 0.915 ;
        RECT  1.575 0.845 1.665 1.075 ;
        RECT  1.505 0.845 1.575 0.915 ;
        RECT  1.435 0.345 1.505 0.915 ;
        RECT  1.285 0.845 1.435 0.915 ;
        RECT  1.215 0.845 1.285 1.075 ;
        RECT  0.945 0.845 1.215 0.915 ;
        RECT  0.835 0.760 0.945 1.045 ;
        RECT  0.525 0.845 0.835 0.915 ;
        RECT  0.455 0.760 0.525 1.010 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.495 1.790 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.495 1.230 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.115 2.100 0.115 ;
        RECT  0.645 -0.115 0.715 0.270 ;
        RECT  0.355 -0.115 0.645 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.855 1.145 2.100 1.375 ;
        RECT  1.785 0.995 1.855 1.375 ;
        RECT  1.475 1.145 1.785 1.375 ;
        RECT  1.405 0.995 1.475 1.375 ;
        RECT  1.095 1.145 1.405 1.375 ;
        RECT  1.025 0.995 1.095 1.375 ;
        RECT  0.715 1.145 1.025 1.375 ;
        RECT  0.645 0.995 0.715 1.375 ;
        RECT  0.335 1.145 0.645 1.375 ;
        RECT  0.265 0.985 0.335 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.195 1.890 0.265 ;
        RECT  0.905 0.345 1.320 0.415 ;
        RECT  0.835 0.185 0.905 0.415 ;
        RECT  0.525 0.345 0.835 0.415 ;
        RECT  0.375 0.545 0.640 0.615 ;
        RECT  0.455 0.260 0.525 0.415 ;
        RECT  0.290 0.345 0.375 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END IND3D3BWP40

MACRO IND3D4BWP40
    CLASS CORE ;
    FOREIGN IND3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.564000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.845 3.045 1.075 ;
        RECT  2.605 0.845 2.955 0.915 ;
        RECT  2.415 0.355 2.815 0.425 ;
        RECT  2.535 0.845 2.605 1.075 ;
        RECT  2.415 0.845 2.535 0.915 ;
        RECT  2.225 0.355 2.415 0.915 ;
        RECT  2.205 0.355 2.225 1.075 ;
        RECT  2.135 0.845 2.205 1.075 ;
        RECT  1.845 0.845 2.135 0.915 ;
        RECT  1.775 0.845 1.845 1.075 ;
        RECT  1.465 0.845 1.775 0.915 ;
        RECT  1.395 0.760 1.465 1.010 ;
        RECT  1.095 0.845 1.395 0.915 ;
        RECT  1.025 0.760 1.095 1.010 ;
        RECT  0.715 0.845 1.025 0.915 ;
        RECT  0.645 0.760 0.715 1.010 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.830 0.495 2.910 0.765 ;
        RECT  2.555 0.495 2.830 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.495 1.960 0.625 ;
        RECT  1.570 0.495 1.650 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.390 0.645 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.115 3.080 0.115 ;
        RECT  1.215 -0.115 1.285 0.275 ;
        RECT  0.905 -0.115 1.215 0.115 ;
        RECT  0.835 -0.115 0.905 0.275 ;
        RECT  0.545 -0.115 0.835 0.115 ;
        RECT  0.425 -0.115 0.545 0.270 ;
        RECT  0.145 -0.115 0.425 0.115 ;
        RECT  0.050 -0.115 0.145 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.795 1.145 3.080 1.375 ;
        RECT  2.725 0.995 2.795 1.375 ;
        RECT  2.415 1.145 2.725 1.375 ;
        RECT  2.345 0.995 2.415 1.375 ;
        RECT  2.035 1.145 2.345 1.375 ;
        RECT  1.965 0.995 2.035 1.375 ;
        RECT  1.655 1.145 1.965 1.375 ;
        RECT  1.585 0.995 1.655 1.375 ;
        RECT  1.285 1.145 1.585 1.375 ;
        RECT  1.215 0.995 1.285 1.375 ;
        RECT  0.905 1.145 1.215 1.375 ;
        RECT  0.835 0.995 0.905 1.375 ;
        RECT  0.530 1.145 0.835 1.375 ;
        RECT  0.450 0.985 0.530 1.375 ;
        RECT  0.140 1.145 0.450 1.375 ;
        RECT  0.050 0.860 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.955 0.845 3.045 1.075 ;
        RECT  2.605 0.845 2.955 0.915 ;
        RECT  2.485 0.355 2.815 0.425 ;
        RECT  2.535 0.845 2.605 1.075 ;
        RECT  2.485 0.845 2.535 0.915 ;
        RECT  1.845 0.845 2.135 0.915 ;
        RECT  1.775 0.845 1.845 1.075 ;
        RECT  1.465 0.845 1.775 0.915 ;
        RECT  1.395 0.760 1.465 1.010 ;
        RECT  1.095 0.845 1.395 0.915 ;
        RECT  1.025 0.760 1.095 1.010 ;
        RECT  0.715 0.845 1.025 0.915 ;
        RECT  0.645 0.760 0.715 1.010 ;
        RECT  2.915 0.195 3.005 0.425 ;
        RECT  1.370 0.195 2.915 0.265 ;
        RECT  1.095 0.345 2.070 0.415 ;
        RECT  1.025 0.185 1.095 0.415 ;
        RECT  0.715 0.345 1.025 0.415 ;
        RECT  0.565 0.545 1.025 0.615 ;
        RECT  0.645 0.255 0.715 0.415 ;
        RECT  0.480 0.345 0.565 0.915 ;
        RECT  0.310 0.345 0.480 0.415 ;
        RECT  0.310 0.845 0.480 0.915 ;
        RECT  0.240 0.195 0.310 0.415 ;
        RECT  0.240 0.845 0.310 1.065 ;
    END
END IND3D4BWP40

MACRO IND3D6BWP40
    CLASS CORE ;
    FOREIGN IND3D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.778500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.355 3.980 0.445 ;
        RECT  3.870 0.710 3.970 1.045 ;
        RECT  3.590 0.710 3.870 0.800 ;
        RECT  3.490 0.710 3.590 1.045 ;
        RECT  3.395 0.710 3.490 0.800 ;
        RECT  3.210 0.355 3.395 0.800 ;
        RECT  3.185 0.355 3.210 1.045 ;
        RECT  3.105 0.355 3.185 0.485 ;
        RECT  3.110 0.710 3.185 1.045 ;
        RECT  2.830 0.710 3.110 0.800 ;
        RECT  2.730 0.710 2.830 1.045 ;
        RECT  2.450 0.710 2.730 0.800 ;
        RECT  2.350 0.710 2.450 1.045 ;
        RECT  2.070 0.710 2.350 0.800 ;
        RECT  1.970 0.710 2.070 1.045 ;
        RECT  1.510 0.710 1.970 0.800 ;
        RECT  1.410 0.710 1.510 1.045 ;
        RECT  1.110 0.710 1.410 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
        RECT  0.625 0.710 0.725 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.070 0.520 4.165 0.905 ;
        RECT  3.490 0.520 4.070 0.620 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.495 2.745 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.400 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.685 -0.115 4.200 0.115 ;
        RECT  1.590 -0.115 1.685 0.260 ;
        RECT  1.325 -0.115 1.590 0.115 ;
        RECT  1.195 -0.115 1.325 0.230 ;
        RECT  0.910 -0.115 1.195 0.115 ;
        RECT  0.780 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.780 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.135 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.135 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.145 4.200 1.375 ;
        RECT  4.060 1.010 4.160 1.375 ;
        RECT  3.780 1.145 4.060 1.375 ;
        RECT  3.680 0.905 3.780 1.375 ;
        RECT  3.400 1.145 3.680 1.375 ;
        RECT  3.300 0.905 3.400 1.375 ;
        RECT  3.020 1.145 3.300 1.375 ;
        RECT  2.930 0.905 3.020 1.375 ;
        RECT  2.640 1.145 2.930 1.375 ;
        RECT  2.540 0.905 2.640 1.375 ;
        RECT  2.260 1.145 2.540 1.375 ;
        RECT  2.160 0.905 2.260 1.375 ;
        RECT  1.880 1.145 2.160 1.375 ;
        RECT  1.790 0.905 1.880 1.375 ;
        RECT  1.690 1.145 1.790 1.375 ;
        RECT  1.595 0.905 1.690 1.375 ;
        RECT  1.310 1.145 1.595 1.375 ;
        RECT  1.215 0.905 1.310 1.375 ;
        RECT  0.900 1.145 1.215 1.375 ;
        RECT  0.805 0.905 0.900 1.375 ;
        RECT  0.520 1.145 0.805 1.375 ;
        RECT  0.420 0.985 0.520 1.375 ;
        RECT  0.135 1.145 0.420 1.375 ;
        RECT  0.050 0.860 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.355 3.980 0.445 ;
        RECT  3.870 0.710 3.970 1.045 ;
        RECT  3.590 0.710 3.870 0.800 ;
        RECT  3.490 0.710 3.590 1.045 ;
        RECT  3.465 0.710 3.490 0.800 ;
        RECT  3.105 0.355 3.115 0.485 ;
        RECT  3.110 0.710 3.115 1.045 ;
        RECT  2.830 0.710 3.110 0.800 ;
        RECT  2.730 0.710 2.830 1.045 ;
        RECT  2.450 0.710 2.730 0.800 ;
        RECT  2.350 0.710 2.450 1.045 ;
        RECT  2.070 0.710 2.350 0.800 ;
        RECT  1.970 0.710 2.070 1.045 ;
        RECT  1.510 0.710 1.970 0.800 ;
        RECT  1.410 0.710 1.510 1.045 ;
        RECT  1.110 0.710 1.410 0.800 ;
        RECT  1.010 0.710 1.110 1.045 ;
        RECT  0.725 0.710 1.010 0.800 ;
        RECT  0.625 0.710 0.725 1.045 ;
        RECT  4.070 0.195 4.150 0.370 ;
        RECT  1.770 0.195 4.070 0.270 ;
        RECT  1.485 0.345 2.870 0.415 ;
        RECT  1.415 0.185 1.485 0.415 ;
        RECT  1.085 0.345 1.415 0.415 ;
        RECT  0.540 0.545 1.350 0.615 ;
        RECT  1.015 0.185 1.085 0.415 ;
        RECT  0.700 0.345 1.015 0.415 ;
        RECT  0.620 0.260 0.700 0.415 ;
        RECT  0.470 0.345 0.540 0.915 ;
        RECT  0.320 0.345 0.470 0.415 ;
        RECT  0.320 0.845 0.470 0.915 ;
        RECT  0.245 0.185 0.320 0.415 ;
        RECT  0.245 0.845 0.320 1.070 ;
    END
END IND3D6BWP40

MACRO IND3D8BWP40
    CLASS CORE ;
    FOREIGN IND3D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.033500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.355 5.360 0.445 ;
        RECT  5.250 0.710 5.350 1.045 ;
        RECT  4.970 0.710 5.250 0.800 ;
        RECT  4.870 0.710 4.970 1.045 ;
        RECT  4.590 0.710 4.870 0.800 ;
        RECT  4.490 0.710 4.590 1.045 ;
        RECT  4.375 0.710 4.490 0.800 ;
        RECT  4.210 0.355 4.375 0.800 ;
        RECT  4.165 0.355 4.210 1.045 ;
        RECT  4.105 0.355 4.165 0.485 ;
        RECT  4.110 0.710 4.165 1.045 ;
        RECT  3.810 0.710 4.110 0.800 ;
        RECT  3.710 0.710 3.810 1.045 ;
        RECT  3.430 0.710 3.710 0.800 ;
        RECT  3.330 0.710 3.430 1.045 ;
        RECT  3.050 0.710 3.330 0.800 ;
        RECT  2.950 0.710 3.050 1.045 ;
        RECT  2.670 0.710 2.950 0.800 ;
        RECT  2.570 0.710 2.670 1.045 ;
        RECT  2.090 0.710 2.570 0.800 ;
        RECT  1.990 0.710 2.090 1.045 ;
        RECT  1.700 0.710 1.990 0.800 ;
        RECT  1.600 0.710 1.700 1.045 ;
        RECT  1.300 0.710 1.600 0.800 ;
        RECT  1.200 0.710 1.300 1.045 ;
        RECT  0.915 0.710 1.200 0.800 ;
        RECT  0.815 0.710 0.915 1.045 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.470 0.520 5.565 0.905 ;
        RECT  4.490 0.520 5.470 0.620 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.670 0.520 3.745 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.555 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 -0.115 5.600 0.115 ;
        RECT  2.180 -0.115 2.280 0.275 ;
        RECT  1.905 -0.115 2.180 0.115 ;
        RECT  1.775 -0.115 1.905 0.230 ;
        RECT  1.515 -0.115 1.775 0.115 ;
        RECT  1.385 -0.115 1.515 0.230 ;
        RECT  1.100 -0.115 1.385 0.115 ;
        RECT  0.970 -0.115 1.100 0.230 ;
        RECT  0.720 -0.115 0.970 0.115 ;
        RECT  0.600 -0.115 0.720 0.275 ;
        RECT  0.325 -0.115 0.600 0.115 ;
        RECT  0.240 -0.115 0.325 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.560 1.145 5.600 1.375 ;
        RECT  5.460 1.010 5.560 1.375 ;
        RECT  5.160 1.145 5.460 1.375 ;
        RECT  5.060 0.895 5.160 1.375 ;
        RECT  4.780 1.145 5.060 1.375 ;
        RECT  4.680 0.895 4.780 1.375 ;
        RECT  4.400 1.145 4.680 1.375 ;
        RECT  4.300 0.895 4.400 1.375 ;
        RECT  4.020 1.145 4.300 1.375 ;
        RECT  3.920 0.895 4.020 1.375 ;
        RECT  3.620 1.145 3.920 1.375 ;
        RECT  3.520 0.895 3.620 1.375 ;
        RECT  3.240 1.145 3.520 1.375 ;
        RECT  3.140 0.895 3.240 1.375 ;
        RECT  2.860 1.145 3.140 1.375 ;
        RECT  2.760 0.895 2.860 1.375 ;
        RECT  2.485 1.145 2.760 1.375 ;
        RECT  2.390 0.895 2.485 1.375 ;
        RECT  2.280 1.145 2.390 1.375 ;
        RECT  2.185 0.895 2.280 1.375 ;
        RECT  1.890 1.145 2.185 1.375 ;
        RECT  1.795 0.895 1.890 1.375 ;
        RECT  1.500 1.145 1.795 1.375 ;
        RECT  1.405 0.895 1.500 1.375 ;
        RECT  1.090 1.145 1.405 1.375 ;
        RECT  0.995 0.895 1.090 1.375 ;
        RECT  0.710 1.145 0.995 1.375 ;
        RECT  0.610 0.985 0.710 1.375 ;
        RECT  0.340 1.145 0.610 1.375 ;
        RECT  0.225 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.355 5.360 0.445 ;
        RECT  5.250 0.710 5.350 1.045 ;
        RECT  4.970 0.710 5.250 0.800 ;
        RECT  4.870 0.710 4.970 1.045 ;
        RECT  4.590 0.710 4.870 0.800 ;
        RECT  4.490 0.710 4.590 1.045 ;
        RECT  4.445 0.710 4.490 0.800 ;
        RECT  3.810 0.710 4.095 0.800 ;
        RECT  3.710 0.710 3.810 1.045 ;
        RECT  3.430 0.710 3.710 0.800 ;
        RECT  3.330 0.710 3.430 1.045 ;
        RECT  3.050 0.710 3.330 0.800 ;
        RECT  2.950 0.710 3.050 1.045 ;
        RECT  2.670 0.710 2.950 0.800 ;
        RECT  2.570 0.710 2.670 1.045 ;
        RECT  2.090 0.710 2.570 0.800 ;
        RECT  1.990 0.710 2.090 1.045 ;
        RECT  1.700 0.710 1.990 0.800 ;
        RECT  1.600 0.710 1.700 1.045 ;
        RECT  1.300 0.710 1.600 0.800 ;
        RECT  1.200 0.710 1.300 1.045 ;
        RECT  0.915 0.710 1.200 0.800 ;
        RECT  0.815 0.710 0.915 1.045 ;
        RECT  5.470 0.195 5.550 0.370 ;
        RECT  2.370 0.195 5.470 0.270 ;
        RECT  2.075 0.375 3.820 0.445 ;
        RECT  0.745 0.525 2.080 0.615 ;
        RECT  2.005 0.185 2.075 0.445 ;
        RECT  1.675 0.375 2.005 0.445 ;
        RECT  1.605 0.185 1.675 0.445 ;
        RECT  1.275 0.375 1.605 0.445 ;
        RECT  1.205 0.185 1.275 0.445 ;
        RECT  0.890 0.375 1.205 0.445 ;
        RECT  0.820 0.185 0.890 0.445 ;
        RECT  0.675 0.345 0.745 0.915 ;
        RECT  0.510 0.345 0.675 0.415 ;
        RECT  0.510 0.845 0.675 0.915 ;
        RECT  0.435 0.185 0.510 0.415 ;
        RECT  0.435 0.845 0.510 1.070 ;
        RECT  0.130 0.345 0.435 0.415 ;
        RECT  0.130 0.845 0.435 0.915 ;
        RECT  0.055 0.185 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.070 ;
    END
END IND3D8BWP40

MACRO IND4D0BWP40
    CLASS CORE ;
    FOREIGN IND4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.105375 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.195 1.225 0.855 ;
        RECT  1.015 0.195 1.155 0.275 ;
        RECT  0.950 0.775 1.155 0.855 ;
        RECT  0.870 0.775 0.950 1.055 ;
        RECT  0.565 0.775 0.870 0.855 ;
        RECT  0.455 0.775 0.565 1.055 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.355 0.945 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.340 0.805 0.690 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 -0.115 1.260 0.115 ;
        RECT  0.250 -0.115 0.330 0.265 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.145 1.260 1.375 ;
        RECT  1.080 0.935 1.160 1.375 ;
        RECT  0.760 1.145 1.080 1.375 ;
        RECT  0.680 0.935 0.760 1.375 ;
        RECT  0.330 1.145 0.680 1.375 ;
        RECT  0.250 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.075 ;
    END
END IND4D0BWP40

MACRO IND4D1BWP40
    CLASS CORE ;
    FOREIGN IND4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.210750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.205 1.225 0.855 ;
        RECT  1.115 0.205 1.155 0.415 ;
        RECT  0.950 0.775 1.155 0.855 ;
        RECT  0.870 0.775 0.950 1.055 ;
        RECT  0.565 0.775 0.870 0.855 ;
        RECT  0.455 0.775 0.565 1.055 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.355 0.945 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.340 0.805 0.690 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.355 0.525 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.330 -0.115 1.260 0.115 ;
        RECT  0.250 -0.115 0.330 0.265 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.145 1.260 1.375 ;
        RECT  1.080 0.935 1.160 1.375 ;
        RECT  0.760 1.145 1.080 1.375 ;
        RECT  0.680 0.935 0.760 1.375 ;
        RECT  0.330 1.145 0.680 1.375 ;
        RECT  0.250 0.985 0.330 1.375 ;
        RECT  0.000 1.145 0.250 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.075 ;
    END
END IND4D1BWP40

MACRO IND4D2BWP40
    CLASS CORE ;
    FOREIGN IND4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.358500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.345 2.205 0.915 ;
        RECT  1.975 0.345 2.135 0.415 ;
        RECT  2.065 0.845 2.135 0.915 ;
        RECT  1.995 0.845 2.065 1.075 ;
        RECT  1.505 0.845 1.995 0.915 ;
        RECT  1.405 0.845 1.505 1.075 ;
        RECT  1.095 0.845 1.405 0.915 ;
        RECT  1.015 0.845 1.095 1.075 ;
        RECT  0.525 0.845 1.015 0.915 ;
        RECT  0.455 0.750 0.525 1.010 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.495 2.000 0.625 ;
        RECT  1.850 0.495 1.930 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.495 1.510 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.090 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.115 2.380 0.115 ;
        RECT  0.620 -0.115 0.715 0.270 ;
        RECT  0.355 -0.115 0.620 0.115 ;
        RECT  0.235 -0.115 0.355 0.270 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 1.145 2.380 1.375 ;
        RECT  2.225 0.995 2.295 1.375 ;
        RECT  1.845 1.145 2.225 1.375 ;
        RECT  1.775 0.995 1.845 1.375 ;
        RECT  1.665 1.145 1.775 1.375 ;
        RECT  1.595 0.995 1.665 1.375 ;
        RECT  1.285 1.145 1.595 1.375 ;
        RECT  1.215 0.995 1.285 1.375 ;
        RECT  0.895 1.145 1.215 1.375 ;
        RECT  0.825 0.995 0.895 1.375 ;
        RECT  0.715 1.145 0.825 1.375 ;
        RECT  0.645 0.995 0.715 1.375 ;
        RECT  0.340 1.145 0.645 1.375 ;
        RECT  0.260 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.845 0.195 2.320 0.265 ;
        RECT  1.775 0.195 1.845 0.415 ;
        RECT  1.380 0.345 1.775 0.415 ;
        RECT  0.800 0.195 1.690 0.265 ;
        RECT  0.525 0.345 1.145 0.415 ;
        RECT  0.375 0.545 0.550 0.615 ;
        RECT  0.455 0.255 0.525 0.415 ;
        RECT  0.290 0.345 0.375 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END IND4D2BWP40

MACRO IND4D4BWP40
    CLASS CORE ;
    FOREIGN IND4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.709000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.770 0.445 ;
        RECT  3.665 0.775 3.745 1.045 ;
        RECT  3.535 0.775 3.665 0.905 ;
        RECT  3.355 0.355 3.535 0.905 ;
        RECT  3.325 0.355 3.355 1.045 ;
        RECT  3.260 0.355 3.325 0.495 ;
        RECT  3.285 0.775 3.325 1.045 ;
        RECT  2.995 0.775 3.285 0.905 ;
        RECT  2.915 0.775 2.995 1.045 ;
        RECT  2.605 0.775 2.915 0.905 ;
        RECT  2.535 0.775 2.605 1.045 ;
        RECT  2.225 0.775 2.535 0.905 ;
        RECT  2.155 0.775 2.225 1.045 ;
        RECT  1.845 0.775 2.155 0.905 ;
        RECT  1.775 0.775 1.845 1.045 ;
        RECT  1.465 0.775 1.775 0.905 ;
        RECT  1.395 0.775 1.465 1.045 ;
        RECT  1.105 0.775 1.395 0.905 ;
        RECT  1.015 0.775 1.105 1.045 ;
        RECT  0.725 0.775 1.015 0.865 ;
        RECT  0.635 0.775 0.725 1.045 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.525 3.885 0.920 ;
        RECT  3.630 0.525 3.815 0.640 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.515 0.525 2.940 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.325 0.515 1.945 0.620 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.390 0.645 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 -0.115 4.060 0.115 ;
        RECT  1.190 -0.115 1.285 0.285 ;
        RECT  0.905 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.905 0.285 ;
        RECT  0.545 -0.115 0.810 0.115 ;
        RECT  0.425 -0.115 0.545 0.270 ;
        RECT  0.145 -0.115 0.425 0.115 ;
        RECT  0.050 -0.115 0.145 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.990 1.145 4.060 1.375 ;
        RECT  3.865 1.020 3.990 1.375 ;
        RECT  3.575 1.145 3.865 1.375 ;
        RECT  3.450 1.020 3.575 1.375 ;
        RECT  3.195 1.145 3.450 1.375 ;
        RECT  3.070 1.020 3.195 1.375 ;
        RECT  2.825 1.145 3.070 1.375 ;
        RECT  2.700 1.020 2.825 1.375 ;
        RECT  2.445 1.145 2.700 1.375 ;
        RECT  2.320 1.020 2.445 1.375 ;
        RECT  2.060 1.145 2.320 1.375 ;
        RECT  1.940 0.990 2.060 1.375 ;
        RECT  1.680 1.145 1.940 1.375 ;
        RECT  1.560 0.990 1.680 1.375 ;
        RECT  1.290 1.145 1.560 1.375 ;
        RECT  1.190 0.980 1.290 1.375 ;
        RECT  0.910 1.145 1.190 1.375 ;
        RECT  0.810 0.980 0.910 1.375 ;
        RECT  0.530 1.145 0.810 1.375 ;
        RECT  0.450 0.985 0.530 1.375 ;
        RECT  0.140 1.145 0.450 1.375 ;
        RECT  0.050 0.810 0.140 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.355 3.770 0.445 ;
        RECT  3.665 0.775 3.745 1.045 ;
        RECT  3.605 0.775 3.665 0.905 ;
        RECT  2.995 0.775 3.255 0.905 ;
        RECT  2.915 0.775 2.995 1.045 ;
        RECT  2.605 0.775 2.915 0.905 ;
        RECT  2.535 0.775 2.605 1.045 ;
        RECT  2.225 0.775 2.535 0.905 ;
        RECT  2.155 0.775 2.225 1.045 ;
        RECT  1.845 0.775 2.155 0.905 ;
        RECT  1.775 0.775 1.845 1.045 ;
        RECT  1.465 0.775 1.775 0.905 ;
        RECT  1.395 0.775 1.465 1.045 ;
        RECT  1.105 0.775 1.395 0.905 ;
        RECT  1.015 0.775 1.105 1.045 ;
        RECT  0.725 0.775 1.015 0.865 ;
        RECT  0.635 0.775 0.725 1.045 ;
        RECT  3.895 0.195 3.965 0.455 ;
        RECT  3.190 0.195 3.895 0.265 ;
        RECT  3.100 0.195 3.190 0.435 ;
        RECT  2.315 0.365 3.100 0.435 ;
        RECT  1.370 0.195 3.010 0.265 ;
        RECT  1.095 0.365 2.070 0.435 ;
        RECT  1.025 0.210 1.095 0.435 ;
        RECT  0.725 0.365 1.025 0.435 ;
        RECT  0.565 0.530 0.995 0.640 ;
        RECT  0.640 0.250 0.725 0.435 ;
        RECT  0.480 0.345 0.565 0.915 ;
        RECT  0.310 0.345 0.480 0.415 ;
        RECT  0.310 0.845 0.480 0.915 ;
        RECT  0.240 0.195 0.310 0.415 ;
        RECT  0.240 0.845 0.310 1.065 ;
    END
END IND4D4BWP40

MACRO INR2D0BWP40
    CLASS CORE ;
    FOREIGN INR2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.064375 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.845 0.805 1.065 ;
        RECT  0.525 0.845 0.700 0.925 ;
        RECT  0.525 0.185 0.580 0.285 ;
        RECT  0.455 0.185 0.525 0.925 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 -0.115 0.840 0.115 ;
        RECT  0.700 -0.115 0.800 0.275 ;
        RECT  0.340 -0.115 0.700 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.345 1.145 0.840 1.375 ;
        RECT  0.225 0.985 0.345 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.055 ;
    END
END INR2D0BWP40

MACRO INR2D1BWP40
    CLASS CORE ;
    FOREIGN INR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.128750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.775 0.805 1.045 ;
        RECT  0.525 0.775 0.700 0.855 ;
        RECT  0.525 0.185 0.580 0.425 ;
        RECT  0.455 0.185 0.525 0.855 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.625 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 -0.115 0.840 0.115 ;
        RECT  0.700 -0.115 0.800 0.275 ;
        RECT  0.340 -0.115 0.700 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.345 1.145 0.840 1.375 ;
        RECT  0.225 0.985 0.345 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.915 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.845 0.315 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.055 ;
    END
END INR2D1BWP40

MACRO INR2D2BWP40
    CLASS CORE ;
    FOREIGN INR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.172500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.730 1.130 0.905 ;
        RECT  1.010 0.215 1.110 0.475 ;
        RECT  0.685 0.385 1.010 0.475 ;
        RECT  0.685 0.730 0.960 0.820 ;
        RECT  0.595 0.385 0.685 0.820 ;
        RECT  0.535 0.385 0.595 0.475 ;
        RECT  0.435 0.215 0.535 0.475 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.545 1.365 0.910 ;
        RECT  1.040 0.545 1.275 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 0.520 0.225 0.650 ;
        RECT  0.035 0.495 0.130 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.400 0.115 ;
        RECT  1.220 -0.115 1.320 0.415 ;
        RECT  0.890 -0.115 1.220 0.115 ;
        RECT  0.810 -0.115 0.890 0.270 ;
        RECT  0.720 -0.115 0.810 0.115 ;
        RECT  0.625 -0.115 0.720 0.280 ;
        RECT  0.330 -0.115 0.625 0.115 ;
        RECT  0.230 -0.115 0.330 0.275 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.145 1.400 1.375 ;
        RECT  0.600 1.030 0.730 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.890 0.990 1.315 1.065 ;
        RECT  0.820 0.890 0.890 1.065 ;
        RECT  0.520 0.890 0.820 0.960 ;
        RECT  0.440 0.820 0.520 0.960 ;
        RECT  0.365 0.545 0.490 0.615 ;
        RECT  0.295 0.345 0.365 0.915 ;
        RECT  0.130 0.345 0.295 0.415 ;
        RECT  0.130 0.845 0.295 0.915 ;
        RECT  0.055 0.190 0.130 0.415 ;
        RECT  0.055 0.845 0.130 1.075 ;
    END
END INR2D2BWP40

MACRO INR2D4BWP40
    CLASS CORE ;
    FOREIGN INR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.368500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.815 2.090 0.905 ;
        RECT  1.980 0.215 2.080 0.465 ;
        RECT  1.855 0.375 1.980 0.465 ;
        RECT  1.700 0.375 1.855 0.905 ;
        RECT  1.645 0.215 1.700 0.905 ;
        RECT  1.600 0.215 1.645 0.465 ;
        RECT  1.595 0.775 1.645 0.905 ;
        RECT  1.110 0.375 1.600 0.465 ;
        RECT  1.010 0.215 1.110 0.465 ;
        RECT  0.725 0.375 1.010 0.465 ;
        RECT  0.625 0.215 0.725 0.465 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.355 2.345 0.640 ;
        RECT  1.980 0.540 2.250 0.640 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.415 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 -0.115 2.380 0.115 ;
        RECT  2.240 -0.115 2.340 0.250 ;
        RECT  1.890 -0.115 2.240 0.115 ;
        RECT  1.790 -0.115 1.890 0.275 ;
        RECT  1.510 -0.115 1.790 0.115 ;
        RECT  1.410 -0.115 1.510 0.275 ;
        RECT  1.300 -0.115 1.410 0.115 ;
        RECT  1.205 -0.115 1.300 0.295 ;
        RECT  0.905 -0.115 1.205 0.115 ;
        RECT  0.800 -0.115 0.905 0.275 ;
        RECT  0.520 -0.115 0.800 0.115 ;
        RECT  0.420 -0.115 0.520 0.275 ;
        RECT  0.135 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.135 0.490 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 2.380 1.375 ;
        RECT  1.200 1.030 1.320 1.375 ;
        RECT  0.910 1.145 1.200 1.375 ;
        RECT  0.780 1.030 0.910 1.375 ;
        RECT  0.530 1.145 0.780 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.135 1.145 0.410 1.375 ;
        RECT  0.050 0.800 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.815 2.090 0.905 ;
        RECT  1.980 0.215 2.080 0.465 ;
        RECT  1.925 0.375 1.980 0.465 ;
        RECT  1.110 0.375 1.575 0.465 ;
        RECT  1.010 0.215 1.110 0.465 ;
        RECT  0.725 0.375 1.010 0.465 ;
        RECT  0.625 0.215 0.725 0.465 ;
        RECT  2.245 0.805 2.315 1.065 ;
        RECT  1.480 0.990 2.245 1.065 ;
        RECT  1.410 0.700 1.480 1.065 ;
        RECT  1.085 0.890 1.410 0.960 ;
        RECT  1.015 0.700 1.085 0.960 ;
        RECT  0.555 0.545 1.065 0.615 ;
        RECT  0.710 0.890 1.015 0.960 ;
        RECT  0.630 0.700 0.710 0.960 ;
        RECT  0.485 0.345 0.555 0.915 ;
        RECT  0.320 0.345 0.485 0.415 ;
        RECT  0.320 0.845 0.485 0.915 ;
        RECT  0.245 0.190 0.320 0.415 ;
        RECT  0.245 0.845 0.320 1.075 ;
    END
END INR2D4BWP40

MACRO INR3D0BWP40
    CLASS CORE ;
    FOREIGN INR3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.074000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.205 0.945 0.415 ;
        RECT  0.840 0.875 0.945 1.065 ;
        RECT  0.545 0.345 0.840 0.415 ;
        RECT  0.525 0.995 0.840 1.065 ;
        RECT  0.525 0.215 0.545 0.415 ;
        RECT  0.455 0.215 0.525 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.915 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.250 ;
        RECT  0.355 -0.115 0.640 0.115 ;
        RECT  0.235 -0.115 0.355 0.220 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.980 1.375 ;
        RECT  0.260 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.345 0.385 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.190 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END INR3D0BWP40

MACRO INR3D1BWP40
    CLASS CORE ;
    FOREIGN INR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.148000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.875 0.945 1.065 ;
        RECT  0.855 0.215 0.925 0.415 ;
        RECT  0.545 0.345 0.855 0.415 ;
        RECT  0.525 0.995 0.840 1.065 ;
        RECT  0.525 0.215 0.545 0.415 ;
        RECT  0.455 0.215 0.525 1.065 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.685 0.915 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.250 ;
        RECT  0.355 -0.115 0.640 0.115 ;
        RECT  0.235 -0.115 0.355 0.220 ;
        RECT  0.000 -0.115 0.235 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.980 1.375 ;
        RECT  0.260 0.995 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.345 0.385 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.190 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END INR3D1BWP40

MACRO INR3D2BWP40
    CLASS CORE ;
    FOREIGN INR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.257000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.825 1.505 0.915 ;
        RECT  1.405 0.245 1.475 0.415 ;
        RECT  1.365 0.340 1.405 0.415 ;
        RECT  1.295 0.340 1.365 0.915 ;
        RECT  1.105 0.340 1.295 0.415 ;
        RECT  1.015 0.185 1.105 0.415 ;
        RECT  0.535 0.340 1.015 0.415 ;
        RECT  0.445 0.215 0.535 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.335 1.645 0.635 ;
        RECT  1.440 0.530 1.565 0.635 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.090 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.740 -0.115 1.820 0.115 ;
        RECT  1.610 -0.115 1.740 0.240 ;
        RECT  1.310 -0.115 1.610 0.115 ;
        RECT  1.190 -0.115 1.310 0.270 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.830 -0.115 0.930 0.270 ;
        RECT  0.720 -0.115 0.830 0.115 ;
        RECT  0.620 -0.115 0.720 0.270 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.260 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.145 1.820 1.375 ;
        RECT  0.620 0.985 0.715 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.235 0.990 0.355 1.375 ;
        RECT  0.000 1.145 0.235 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.635 0.805 1.705 1.065 ;
        RECT  0.800 0.995 1.635 1.065 ;
        RECT  0.535 0.845 1.145 0.915 ;
        RECT  0.450 0.845 0.535 1.010 ;
        RECT  0.375 0.520 0.500 0.630 ;
        RECT  0.290 0.345 0.375 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END INR3D2BWP40

MACRO INR3D4BWP40
    CLASS CORE ;
    FOREIGN INR3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.492000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.215 3.045 0.425 ;
        RECT  2.605 0.335 2.955 0.425 ;
        RECT  2.415 0.815 2.810 0.925 ;
        RECT  2.535 0.215 2.605 0.425 ;
        RECT  2.415 0.335 2.535 0.425 ;
        RECT  2.225 0.335 2.415 0.925 ;
        RECT  2.205 0.215 2.225 0.925 ;
        RECT  2.155 0.215 2.205 0.425 ;
        RECT  1.845 0.335 2.155 0.425 ;
        RECT  1.775 0.195 1.845 0.425 ;
        RECT  1.465 0.335 1.775 0.425 ;
        RECT  1.395 0.195 1.465 0.425 ;
        RECT  1.105 0.335 1.395 0.425 ;
        RECT  1.015 0.195 1.105 0.425 ;
        RECT  0.725 0.335 1.015 0.425 ;
        RECT  0.635 0.215 0.725 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.525 2.905 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.520 1.925 0.625 ;
        RECT  1.435 0.520 1.505 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.385 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.825 -0.115 3.080 0.115 ;
        RECT  2.700 -0.115 2.825 0.240 ;
        RECT  2.445 -0.115 2.700 0.115 ;
        RECT  2.320 -0.115 2.445 0.240 ;
        RECT  2.060 -0.115 2.320 0.115 ;
        RECT  1.940 -0.115 2.060 0.250 ;
        RECT  1.680 -0.115 1.940 0.115 ;
        RECT  1.560 -0.115 1.680 0.250 ;
        RECT  1.310 -0.115 1.560 0.115 ;
        RECT  1.190 -0.115 1.310 0.250 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.260 ;
        RECT  0.530 -0.115 0.810 0.115 ;
        RECT  0.450 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.450 0.115 ;
        RECT  0.050 -0.115 0.140 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 1.145 3.080 1.375 ;
        RECT  1.190 0.985 1.285 1.375 ;
        RECT  0.905 1.145 1.190 1.375 ;
        RECT  0.810 0.985 0.905 1.375 ;
        RECT  0.545 1.145 0.810 1.375 ;
        RECT  0.425 0.990 0.545 1.375 ;
        RECT  0.145 1.145 0.425 1.375 ;
        RECT  0.050 0.860 0.145 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.955 0.215 3.045 0.425 ;
        RECT  2.605 0.335 2.955 0.425 ;
        RECT  2.485 0.815 2.810 0.925 ;
        RECT  2.535 0.215 2.605 0.425 ;
        RECT  2.485 0.335 2.535 0.425 ;
        RECT  1.845 0.335 2.135 0.425 ;
        RECT  1.775 0.195 1.845 0.425 ;
        RECT  1.465 0.335 1.775 0.425 ;
        RECT  1.395 0.195 1.465 0.425 ;
        RECT  1.105 0.335 1.395 0.425 ;
        RECT  1.015 0.195 1.105 0.425 ;
        RECT  0.725 0.335 1.015 0.425 ;
        RECT  0.635 0.215 0.725 0.425 ;
        RECT  2.935 0.760 3.030 1.065 ;
        RECT  1.370 0.995 2.935 1.065 ;
        RECT  0.725 0.845 2.070 0.915 ;
        RECT  0.565 0.520 0.995 0.630 ;
        RECT  0.640 0.845 0.725 1.010 ;
        RECT  0.485 0.345 0.565 0.915 ;
        RECT  0.310 0.345 0.485 0.415 ;
        RECT  0.310 0.845 0.485 0.915 ;
        RECT  0.240 0.195 0.310 0.415 ;
        RECT  0.240 0.845 0.310 1.065 ;
    END
END INR3D4BWP40

MACRO INR4D0BWP40
    CLASS CORE ;
    FOREIGN INR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.096625 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.305 1.225 1.050 ;
        RECT  0.950 0.305 1.155 0.385 ;
        RECT  1.015 0.980 1.155 1.050 ;
        RECT  0.870 0.205 0.950 0.385 ;
        RECT  0.565 0.305 0.870 0.385 ;
        RECT  0.455 0.205 0.565 0.385 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.470 0.805 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.655 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 -0.115 1.260 0.115 ;
        RECT  1.060 -0.115 1.180 0.220 ;
        RECT  0.780 -0.115 1.060 0.115 ;
        RECT  0.655 -0.115 0.780 0.215 ;
        RECT  0.330 -0.115 0.655 0.115 ;
        RECT  0.250 -0.115 0.330 0.270 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.145 1.260 1.375 ;
        RECT  0.230 1.020 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.950 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.880 0.315 0.950 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.880 0.130 1.075 ;
    END
END INR4D0BWP40

MACRO INR4D1BWP40
    CLASS CORE ;
    FOREIGN INR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.193250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.305 1.225 0.905 ;
        RECT  1.155 0.305 1.170 1.065 ;
        RECT  0.565 0.305 1.155 0.385 ;
        RECT  1.090 0.800 1.155 1.065 ;
        RECT  0.455 0.205 0.565 0.385 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.470 0.805 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 -0.115 1.260 0.115 ;
        RECT  1.060 -0.115 1.180 0.220 ;
        RECT  0.780 -0.115 1.060 0.115 ;
        RECT  0.655 -0.115 0.780 0.215 ;
        RECT  0.330 -0.115 0.655 0.115 ;
        RECT  0.250 -0.115 0.330 0.270 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.145 1.260 1.375 ;
        RECT  0.230 1.020 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.950 ;
        RECT  0.130 0.345 0.315 0.415 ;
        RECT  0.130 0.880 0.315 0.950 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.880 0.130 1.075 ;
    END
END INR4D1BWP40

MACRO INR4D2BWP40
    CLASS CORE ;
    FOREIGN INR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.313500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.360 2.205 0.900 ;
        RECT  2.065 0.360 2.135 0.450 ;
        RECT  1.995 0.810 2.135 0.900 ;
        RECT  1.975 0.215 2.065 0.450 ;
        RECT  1.505 0.360 1.975 0.450 ;
        RECT  1.405 0.215 1.505 0.450 ;
        RECT  1.105 0.360 1.405 0.450 ;
        RECT  1.015 0.215 1.105 0.450 ;
        RECT  0.535 0.360 1.015 0.450 ;
        RECT  0.445 0.215 0.535 0.450 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.520 2.040 0.625 ;
        RECT  1.685 0.520 1.785 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.520 1.570 0.625 ;
        RECT  1.265 0.520 1.365 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.520 1.155 0.625 ;
        RECT  0.840 0.520 0.950 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 -0.115 2.380 0.115 ;
        RECT  2.230 -0.115 2.315 0.275 ;
        RECT  1.865 -0.115 2.230 0.115 ;
        RECT  1.780 -0.115 1.865 0.275 ;
        RECT  1.680 -0.115 1.780 0.115 ;
        RECT  1.575 -0.115 1.680 0.275 ;
        RECT  1.310 -0.115 1.575 0.115 ;
        RECT  1.190 -0.115 1.310 0.270 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.830 -0.115 0.930 0.280 ;
        RECT  0.720 -0.115 0.830 0.115 ;
        RECT  0.620 -0.115 0.720 0.280 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.260 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.145 2.380 1.375 ;
        RECT  0.620 0.985 0.715 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.235 0.990 0.355 1.375 ;
        RECT  0.000 1.145 0.235 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.870 0.995 2.320 1.065 ;
        RECT  1.780 0.845 1.870 1.065 ;
        RECT  1.380 0.845 1.780 0.915 ;
        RECT  0.800 0.995 1.690 1.065 ;
        RECT  0.535 0.845 1.145 0.915 ;
        RECT  0.450 0.845 0.535 1.010 ;
        RECT  0.375 0.520 0.500 0.630 ;
        RECT  0.290 0.345 0.375 0.915 ;
        RECT  0.120 0.345 0.290 0.415 ;
        RECT  0.120 0.845 0.290 0.915 ;
        RECT  0.050 0.195 0.120 0.415 ;
        RECT  0.050 0.845 0.120 1.065 ;
    END
END INR4D2BWP40

MACRO INR4D4BWP40
    CLASS CORE ;
    FOREIGN INR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.611000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.835 3.770 0.905 ;
        RECT  3.665 0.215 3.745 0.445 ;
        RECT  3.535 0.355 3.665 0.445 ;
        RECT  3.355 0.355 3.535 0.905 ;
        RECT  3.325 0.215 3.355 0.905 ;
        RECT  3.285 0.215 3.325 0.445 ;
        RECT  3.260 0.765 3.325 0.905 ;
        RECT  2.995 0.355 3.285 0.445 ;
        RECT  2.915 0.215 2.995 0.445 ;
        RECT  2.605 0.355 2.915 0.445 ;
        RECT  2.535 0.215 2.605 0.445 ;
        RECT  2.225 0.355 2.535 0.445 ;
        RECT  2.155 0.215 2.225 0.445 ;
        RECT  1.845 0.355 2.155 0.445 ;
        RECT  1.775 0.215 1.845 0.445 ;
        RECT  1.465 0.355 1.775 0.445 ;
        RECT  1.395 0.215 1.465 0.445 ;
        RECT  1.105 0.355 1.395 0.445 ;
        RECT  1.015 0.215 1.105 0.445 ;
        RECT  0.725 0.355 1.015 0.445 ;
        RECT  0.635 0.215 0.725 0.445 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.805 0.520 3.915 0.765 ;
        RECT  3.630 0.520 3.805 0.635 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.515 2.935 0.765 ;
        RECT  2.515 0.515 2.835 0.620 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.515 1.945 0.620 ;
        RECT  1.405 0.515 1.505 0.765 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.390 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.970 -0.115 4.060 0.115 ;
        RECT  3.890 -0.115 3.970 0.435 ;
        RECT  3.575 -0.115 3.890 0.115 ;
        RECT  3.450 -0.115 3.575 0.240 ;
        RECT  3.195 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.195 0.240 ;
        RECT  2.825 -0.115 3.070 0.115 ;
        RECT  2.700 -0.115 2.825 0.240 ;
        RECT  2.445 -0.115 2.700 0.115 ;
        RECT  2.320 -0.115 2.445 0.240 ;
        RECT  2.060 -0.115 2.320 0.115 ;
        RECT  1.940 -0.115 2.060 0.270 ;
        RECT  1.680 -0.115 1.940 0.115 ;
        RECT  1.560 -0.115 1.680 0.270 ;
        RECT  1.290 -0.115 1.560 0.115 ;
        RECT  1.190 -0.115 1.290 0.280 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.910 0.280 ;
        RECT  0.530 -0.115 0.810 0.115 ;
        RECT  0.450 -0.115 0.530 0.275 ;
        RECT  0.140 -0.115 0.450 0.115 ;
        RECT  0.050 -0.115 0.140 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.285 1.145 4.060 1.375 ;
        RECT  1.190 0.985 1.285 1.375 ;
        RECT  0.905 1.145 1.190 1.375 ;
        RECT  0.810 0.985 0.905 1.375 ;
        RECT  0.545 1.145 0.810 1.375 ;
        RECT  0.425 0.990 0.545 1.375 ;
        RECT  0.145 1.145 0.425 1.375 ;
        RECT  0.050 0.860 0.145 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.835 3.770 0.905 ;
        RECT  3.665 0.215 3.745 0.445 ;
        RECT  3.605 0.355 3.665 0.445 ;
        RECT  2.995 0.355 3.255 0.445 ;
        RECT  2.915 0.215 2.995 0.445 ;
        RECT  2.605 0.355 2.915 0.445 ;
        RECT  2.535 0.215 2.605 0.445 ;
        RECT  2.225 0.355 2.535 0.445 ;
        RECT  2.155 0.215 2.225 0.445 ;
        RECT  1.845 0.355 2.155 0.445 ;
        RECT  1.775 0.215 1.845 0.445 ;
        RECT  1.465 0.355 1.775 0.445 ;
        RECT  1.395 0.215 1.465 0.445 ;
        RECT  1.105 0.355 1.395 0.445 ;
        RECT  1.015 0.215 1.105 0.445 ;
        RECT  0.725 0.355 1.015 0.445 ;
        RECT  0.635 0.215 0.725 0.445 ;
        RECT  3.870 0.860 3.985 1.065 ;
        RECT  3.190 0.995 3.870 1.065 ;
        RECT  3.100 0.845 3.190 1.065 ;
        RECT  2.315 0.845 3.100 0.915 ;
        RECT  1.370 0.995 3.010 1.065 ;
        RECT  1.095 0.845 2.070 0.915 ;
        RECT  1.025 0.845 1.095 1.070 ;
        RECT  0.725 0.845 1.025 0.915 ;
        RECT  0.565 0.520 0.995 0.630 ;
        RECT  0.640 0.845 0.725 1.010 ;
        RECT  0.480 0.345 0.565 0.915 ;
        RECT  0.310 0.345 0.480 0.415 ;
        RECT  0.310 0.845 0.480 0.915 ;
        RECT  0.240 0.195 0.310 0.415 ;
        RECT  0.240 0.845 0.310 1.065 ;
    END
END INR4D4BWP40

MACRO INVD0BWP40
    CLASS CORE ;
    FOREIGN INVD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.056000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.185 0.385 1.075 ;
        RECT  0.280 0.185 0.315 0.300 ;
        RECT  0.290 0.965 0.315 1.075 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.080 -0.115 0.150 0.300 ;
        RECT  0.000 -0.115 0.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.145 0.420 1.375 ;
        RECT  0.080 0.965 0.150 1.375 ;
        RECT  0.000 1.145 0.080 1.375 ;
        END
    END VDD
END INVD0BWP40

MACRO INVD10BWP40
    CLASS CORE ;
    FOREIGN INVD10BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.600000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.475 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.435 0.695 1.505 1.045 ;
        RECT  1.435 0.185 1.475 0.465 ;
        RECT  1.405 0.185 1.435 1.045 ;
        RECT  1.225 0.300 1.405 0.885 ;
        RECT  1.095 0.300 1.225 0.465 ;
        RECT  1.095 0.695 1.225 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.320000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.045 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 -0.115 2.100 0.115 ;
        RECT  1.975 -0.115 2.045 0.465 ;
        RECT  1.690 -0.115 1.975 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.685 2.050 1.375 ;
        RECT  1.690 1.145 1.970 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.505 0.300 1.785 0.465 ;
        RECT  1.505 0.695 1.785 0.885 ;
        RECT  1.095 0.300 1.155 0.465 ;
        RECT  1.095 0.695 1.155 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END INVD10BWP40

MACRO INVD12BWP40
    CLASS CORE ;
    FOREIGN INVD12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.575 0.300 1.785 0.465 ;
        RECT  1.575 0.695 1.785 0.885 ;
        RECT  1.505 0.300 1.575 0.885 ;
        RECT  1.475 0.300 1.505 1.045 ;
        RECT  1.405 0.185 1.475 1.045 ;
        RECT  1.225 0.300 1.405 0.885 ;
        RECT  1.095 0.300 1.225 0.465 ;
        RECT  1.095 0.695 1.225 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.045 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.425 -0.115 2.520 0.115 ;
        RECT  2.355 -0.115 2.425 0.465 ;
        RECT  2.070 -0.115 2.355 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.145 2.520 1.375 ;
        RECT  2.350 0.685 2.430 1.375 ;
        RECT  2.070 1.145 2.350 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.645 0.300 1.785 0.465 ;
        RECT  1.645 0.695 1.785 0.885 ;
        RECT  1.095 0.300 1.155 0.465 ;
        RECT  1.095 0.695 1.155 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END INVD12BWP40

MACRO INVD14BWP40
    CLASS CORE ;
    FOREIGN INVD14BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.868000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.595 0.300 1.785 0.465 ;
        RECT  1.595 0.695 1.785 0.885 ;
        RECT  1.505 0.300 1.595 0.885 ;
        RECT  1.475 0.300 1.505 1.045 ;
        RECT  1.405 0.185 1.475 1.045 ;
        RECT  1.225 0.300 1.405 0.885 ;
        RECT  1.095 0.300 1.225 0.465 ;
        RECT  1.095 0.695 1.225 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.448000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.045 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.115 2.940 0.115 ;
        RECT  2.750 -0.115 2.840 0.465 ;
        RECT  2.450 -0.115 2.750 0.115 ;
        RECT  2.330 -0.115 2.450 0.230 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.230 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.230 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.230 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.230 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.230 ;
        RECT  0.150 -0.115 0.430 0.115 ;
        RECT  0.070 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.845 1.145 2.940 1.375 ;
        RECT  2.755 0.685 2.845 1.375 ;
        RECT  2.450 1.145 2.755 1.375 ;
        RECT  2.330 0.955 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 0.955 2.070 1.375 ;
        RECT  1.690 1.145 1.950 1.375 ;
        RECT  1.590 0.965 1.690 1.375 ;
        RECT  1.310 1.145 1.590 1.375 ;
        RECT  1.190 0.955 1.310 1.375 ;
        RECT  0.930 1.145 1.190 1.375 ;
        RECT  0.810 0.955 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.955 0.550 1.375 ;
        RECT  0.150 1.145 0.430 1.375 ;
        RECT  0.070 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.545 0.185 2.635 0.465 ;
        RECT  2.545 0.695 2.635 1.035 ;
        RECT  2.235 0.300 2.545 0.465 ;
        RECT  2.235 0.695 2.545 0.885 ;
        RECT  2.165 0.185 2.235 0.465 ;
        RECT  2.165 0.695 2.235 1.035 ;
        RECT  1.855 0.300 2.165 0.465 ;
        RECT  1.855 0.695 2.165 0.885 ;
        RECT  1.785 0.185 1.855 0.465 ;
        RECT  1.785 0.695 1.855 1.035 ;
        RECT  1.645 0.300 1.785 0.465 ;
        RECT  1.645 0.695 1.785 0.885 ;
        RECT  1.095 0.300 1.155 0.465 ;
        RECT  1.095 0.695 1.155 0.885 ;
        RECT  1.025 0.185 1.095 0.465 ;
        RECT  1.025 0.695 1.095 1.035 ;
        RECT  0.715 0.300 1.025 0.465 ;
        RECT  0.715 0.695 1.025 0.885 ;
        RECT  0.645 0.185 0.715 0.465 ;
        RECT  0.645 0.695 0.715 1.035 ;
        RECT  0.335 0.300 0.645 0.465 ;
        RECT  0.335 0.695 0.645 0.885 ;
        RECT  0.265 0.185 0.335 0.465 ;
        RECT  0.265 0.695 0.335 1.035 ;
    END
END INVD14BWP40

MACRO INVD16BWP40
    CLASS CORE ;
    FOREIGN INVD16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.575 0.300 1.765 0.465 ;
        RECT  1.575 0.695 1.765 0.885 ;
        RECT  1.505 0.300 1.575 0.885 ;
        RECT  1.455 0.300 1.505 1.045 ;
        RECT  1.385 0.185 1.455 1.045 ;
        RECT  1.225 0.300 1.385 0.885 ;
        RECT  1.075 0.300 1.225 0.465 ;
        RECT  1.075 0.695 1.225 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.512000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.050 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.465 ;
        RECT  2.810 -0.115 3.095 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.685 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.645 0.300 1.765 0.465 ;
        RECT  1.645 0.695 1.765 0.885 ;
        RECT  1.075 0.300 1.155 0.465 ;
        RECT  1.075 0.695 1.155 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END INVD16BWP40

MACRO INVD18BWP40
    CLASS CORE ;
    FOREIGN INVD18BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.080000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.575 0.300 1.765 0.465 ;
        RECT  1.575 0.695 1.765 0.885 ;
        RECT  1.505 0.300 1.575 0.885 ;
        RECT  1.455 0.300 1.505 1.045 ;
        RECT  1.385 0.185 1.455 1.045 ;
        RECT  1.225 0.300 1.385 0.885 ;
        RECT  1.075 0.300 1.225 0.465 ;
        RECT  1.075 0.695 1.225 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.576000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.050 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.585 -0.115 3.640 0.115 ;
        RECT  3.515 -0.115 3.585 0.465 ;
        RECT  3.190 -0.115 3.515 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.685 3.590 1.375 ;
        RECT  3.190 1.145 3.510 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.575 0.965 1.670 1.375 ;
        RECT  1.290 1.145 1.575 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.215 0.300 2.525 0.465 ;
        RECT  2.215 0.695 2.525 0.885 ;
        RECT  2.145 0.185 2.215 0.465 ;
        RECT  2.145 0.695 2.215 1.035 ;
        RECT  1.835 0.300 2.145 0.465 ;
        RECT  1.835 0.695 2.145 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.645 0.300 1.765 0.465 ;
        RECT  1.645 0.695 1.765 0.885 ;
        RECT  1.075 0.300 1.155 0.465 ;
        RECT  1.075 0.695 1.155 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END INVD18BWP40

MACRO INVD1BWP40
    CLASS CORE ;
    FOREIGN INVD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.112000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.185 0.385 1.045 ;
        RECT  0.280 0.185 0.315 0.425 ;
        RECT  0.290 0.710 0.315 1.045 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 -0.115 0.420 0.115 ;
        RECT  0.080 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.145 0.420 1.375 ;
        RECT  0.080 0.845 0.150 1.375 ;
        RECT  0.000 1.145 0.080 1.375 ;
        END
    END VDD
END INVD1BWP40

MACRO INVD20BWP40
    CLASS CORE ;
    FOREIGN INVD20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.208000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.275 0.300 2.525 0.465 ;
        RECT  2.275 0.695 2.525 0.885 ;
        RECT  2.215 0.300 2.275 0.885 ;
        RECT  2.135 0.185 2.215 1.045 ;
        RECT  2.125 0.185 2.135 0.885 ;
        RECT  1.925 0.300 2.125 0.885 ;
        RECT  1.835 0.300 1.925 0.465 ;
        RECT  1.835 0.695 1.925 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.640000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.620 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.465 ;
        RECT  3.570 -0.115 3.935 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.685 4.010 1.375 ;
        RECT  3.570 1.145 3.930 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.955 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.525 0.695 2.595 1.035 ;
        RECT  2.345 0.300 2.525 0.465 ;
        RECT  2.345 0.695 2.525 0.885 ;
        RECT  1.835 0.300 1.855 0.465 ;
        RECT  1.835 0.695 1.855 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END INVD20BWP40

MACRO INVD24BWP40
    CLASS CORE ;
    FOREIGN INVD24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.440000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.595 0.300 2.905 0.465 ;
        RECT  2.595 0.695 2.905 0.885 ;
        RECT  2.555 0.185 2.595 0.465 ;
        RECT  2.555 0.695 2.595 1.035 ;
        RECT  2.525 0.185 2.555 1.035 ;
        RECT  2.215 0.300 2.525 0.885 ;
        RECT  2.205 0.185 2.215 1.045 ;
        RECT  2.135 0.185 2.205 0.465 ;
        RECT  2.135 0.695 2.205 1.045 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.768000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 1.815 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 -0.115 4.760 0.115 ;
        RECT  4.600 -0.115 4.700 0.455 ;
        RECT  4.330 -0.115 4.600 0.115 ;
        RECT  4.210 -0.115 4.330 0.230 ;
        RECT  3.950 -0.115 4.210 0.115 ;
        RECT  3.830 -0.115 3.950 0.230 ;
        RECT  3.570 -0.115 3.830 0.115 ;
        RECT  3.450 -0.115 3.570 0.230 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.230 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.230 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.230 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.230 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.230 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.230 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.230 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.230 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.700 1.145 4.760 1.375 ;
        RECT  4.600 0.695 4.700 1.375 ;
        RECT  4.330 1.145 4.600 1.375 ;
        RECT  4.210 0.955 4.330 1.375 ;
        RECT  3.950 1.145 4.210 1.375 ;
        RECT  3.830 0.955 3.950 1.375 ;
        RECT  3.570 1.145 3.830 1.375 ;
        RECT  3.450 0.955 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.955 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.955 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.955 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.955 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.955 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.955 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.955 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.955 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.425 0.185 4.495 0.465 ;
        RECT  4.425 0.695 4.495 1.035 ;
        RECT  4.115 0.300 4.425 0.465 ;
        RECT  4.115 0.695 4.425 0.885 ;
        RECT  4.045 0.185 4.115 0.465 ;
        RECT  4.045 0.695 4.115 1.035 ;
        RECT  3.735 0.300 4.045 0.465 ;
        RECT  3.735 0.695 4.045 0.885 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.665 0.695 3.735 1.035 ;
        RECT  3.355 0.300 3.665 0.465 ;
        RECT  3.355 0.695 3.665 0.885 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.285 0.695 3.355 1.035 ;
        RECT  2.975 0.300 3.285 0.465 ;
        RECT  2.975 0.695 3.285 0.885 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.905 0.695 2.975 1.035 ;
        RECT  2.625 0.300 2.905 0.465 ;
        RECT  2.625 0.695 2.905 0.885 ;
        RECT  1.835 0.300 2.135 0.465 ;
        RECT  1.835 0.695 2.135 0.885 ;
        RECT  1.765 0.185 1.835 0.465 ;
        RECT  1.765 0.695 1.835 1.035 ;
        RECT  1.455 0.300 1.765 0.465 ;
        RECT  1.455 0.695 1.765 0.885 ;
        RECT  1.385 0.185 1.455 0.465 ;
        RECT  1.385 0.695 1.455 1.035 ;
        RECT  1.075 0.300 1.385 0.465 ;
        RECT  1.075 0.695 1.385 0.885 ;
        RECT  1.005 0.185 1.075 0.465 ;
        RECT  1.005 0.695 1.075 1.035 ;
        RECT  0.695 0.300 1.005 0.465 ;
        RECT  0.695 0.695 1.005 0.885 ;
        RECT  0.625 0.185 0.695 0.465 ;
        RECT  0.625 0.695 0.695 1.035 ;
        RECT  0.315 0.300 0.625 0.465 ;
        RECT  0.315 0.695 0.625 0.885 ;
        RECT  0.245 0.185 0.315 0.465 ;
        RECT  0.245 0.695 0.315 1.035 ;
    END
END INVD24BWP40

MACRO INVD2BWP40
    CLASS CORE ;
    FOREIGN INVD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.355 0.385 0.790 ;
        RECT  0.315 0.185 0.320 0.790 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.710 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.245 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.285 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.145 0.560 1.375 ;
        RECT  0.430 0.845 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END INVD2BWP40

MACRO INVD3BWP40
    CLASS CORE ;
    FOREIGN INVD3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.228000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 0.185 0.805 0.445 ;
        RECT  0.700 0.735 0.805 1.045 ;
        RECT  0.525 0.735 0.700 0.815 ;
        RECT  0.525 0.355 0.690 0.445 ;
        RECT  0.455 0.355 0.525 0.815 ;
        RECT  0.320 0.355 0.455 0.445 ;
        RECT  0.315 0.735 0.455 0.815 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.735 0.315 1.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.300 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 -0.115 0.840 0.115 ;
        RECT  0.470 -0.115 0.550 0.285 ;
        RECT  0.140 -0.115 0.470 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.145 0.840 1.375 ;
        RECT  0.450 0.910 0.570 1.375 ;
        RECT  0.140 1.145 0.450 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END INVD3BWP40

MACRO INVD4BWP40
    CLASS CORE ;
    FOREIGN INVD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.660 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.595 0.705 0.665 0.820 ;
        RECT  0.595 0.310 0.660 0.445 ;
        RECT  0.385 0.310 0.595 0.820 ;
        RECT  0.320 0.310 0.385 0.445 ;
        RECT  0.315 0.705 0.385 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.115 0.980 0.115 ;
        RECT  0.850 -0.115 0.930 0.465 ;
        RECT  0.560 -0.115 0.850 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.850 0.695 0.930 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END INVD4BWP40

MACRO INVD5BWP40
    CLASS CORE ;
    FOREIGN INVD5BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.364000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.735 0.705 1.105 0.820 ;
        RECT  0.740 0.310 1.100 0.445 ;
        RECT  0.735 0.185 0.740 0.445 ;
        RECT  0.665 0.185 0.735 1.030 ;
        RECT  0.660 0.185 0.665 0.820 ;
        RECT  0.525 0.310 0.660 0.820 ;
        RECT  0.315 0.310 0.525 0.445 ;
        RECT  0.315 0.705 0.525 0.820 ;
        RECT  0.245 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.160000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.420 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.980 -0.115 1.260 0.115 ;
        RECT  0.860 -0.115 0.980 0.240 ;
        RECT  0.560 -0.115 0.860 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.145 1.260 1.375 ;
        RECT  0.850 0.890 0.970 1.375 ;
        RECT  0.560 1.145 0.850 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.100 0.185 1.180 0.445 ;
        RECT  1.105 0.705 1.175 1.030 ;
        RECT  0.805 0.705 1.105 0.820 ;
        RECT  0.805 0.310 1.100 0.445 ;
        RECT  0.315 0.310 0.455 0.445 ;
        RECT  0.315 0.705 0.455 0.820 ;
        RECT  0.245 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END INVD5BWP40

MACRO INVD6BWP40
    CLASS CORE ;
    FOREIGN INVD6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.735 0.705 1.045 0.820 ;
        RECT  0.740 0.310 1.040 0.445 ;
        RECT  0.660 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.595 0.705 0.665 0.820 ;
        RECT  0.595 0.310 0.660 0.445 ;
        RECT  0.385 0.310 0.595 0.820 ;
        RECT  0.315 0.310 0.385 0.445 ;
        RECT  0.315 0.705 0.385 0.820 ;
        RECT  0.245 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 -0.115 1.400 0.115 ;
        RECT  1.235 -0.115 1.305 0.400 ;
        RECT  0.950 -0.115 1.235 0.115 ;
        RECT  0.830 -0.115 0.950 0.240 ;
        RECT  0.560 -0.115 0.830 0.115 ;
        RECT  0.440 -0.115 0.560 0.240 ;
        RECT  0.140 -0.115 0.440 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.145 1.400 1.375 ;
        RECT  1.235 0.725 1.305 1.375 ;
        RECT  0.960 1.145 1.235 1.375 ;
        RECT  0.830 0.890 0.960 1.375 ;
        RECT  0.560 1.145 0.830 1.375 ;
        RECT  0.440 0.890 0.560 1.375 ;
        RECT  0.140 1.145 0.440 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.185 1.120 0.445 ;
        RECT  1.045 0.705 1.115 1.030 ;
        RECT  0.735 0.705 1.045 0.820 ;
        RECT  0.740 0.310 1.040 0.445 ;
        RECT  0.665 0.185 0.740 0.445 ;
        RECT  0.665 0.705 0.735 1.030 ;
        RECT  0.245 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END INVD6BWP40

MACRO INVD8BWP40
    CLASS CORE ;
    FOREIGN INVD8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.508000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.015 0.185 1.095 0.445 ;
        RECT  1.020 0.705 1.090 1.030 ;
        RECT  0.735 0.705 1.020 0.820 ;
        RECT  0.735 0.310 1.015 0.445 ;
        RECT  0.700 0.310 0.735 0.820 ;
        RECT  0.695 0.185 0.700 0.820 ;
        RECT  0.625 0.185 0.695 1.030 ;
        RECT  0.620 0.185 0.625 0.820 ;
        RECT  0.385 0.310 0.620 0.820 ;
        RECT  0.320 0.310 0.385 0.445 ;
        RECT  0.315 0.705 0.385 0.820 ;
        RECT  0.240 0.185 0.320 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.250 0.615 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.770 0.400 ;
        RECT  1.305 -0.115 1.690 0.115 ;
        RECT  1.185 -0.115 1.305 0.240 ;
        RECT  0.910 -0.115 1.185 0.115 ;
        RECT  0.790 -0.115 0.910 0.240 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.240 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.145 1.820 1.375 ;
        RECT  1.690 0.725 1.770 1.375 ;
        RECT  1.310 1.145 1.690 1.375 ;
        RECT  1.190 0.890 1.310 1.375 ;
        RECT  0.915 1.145 1.190 1.375 ;
        RECT  0.795 0.890 0.915 1.375 ;
        RECT  0.530 1.145 0.795 1.375 ;
        RECT  0.410 0.890 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.415 0.185 1.505 0.445 ;
        RECT  1.420 0.705 1.490 1.030 ;
        RECT  1.090 0.705 1.420 0.820 ;
        RECT  1.095 0.310 1.415 0.445 ;
        RECT  1.015 0.185 1.095 0.445 ;
        RECT  1.020 0.705 1.090 1.030 ;
        RECT  0.805 0.705 1.020 0.820 ;
        RECT  0.805 0.310 1.015 0.445 ;
        RECT  0.240 0.185 0.315 0.445 ;
        RECT  0.245 0.705 0.315 1.030 ;
    END
END INVD8BWP40

MACRO IOA21D0BWP40
    CLASS CORE ;
    FOREIGN IOA21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.055625 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.210 0.945 0.790 ;
        RECT  0.820 0.210 0.875 0.285 ;
        RECT  0.725 0.720 0.875 0.790 ;
        RECT  0.655 0.720 0.725 1.025 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.425 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.560 -0.115 0.980 0.115 ;
        RECT  0.440 -0.115 0.560 0.275 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.145 0.980 1.375 ;
        RECT  0.840 0.950 0.920 1.375 ;
        RECT  0.540 1.145 0.840 1.375 ;
        RECT  0.420 0.995 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.950 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.510 0.345 0.580 0.915 ;
        RECT  0.350 0.345 0.510 0.415 ;
        RECT  0.320 0.845 0.510 0.915 ;
        RECT  0.280 0.215 0.350 0.415 ;
        RECT  0.240 0.845 0.320 1.050 ;
        RECT  0.140 0.215 0.280 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA21D0BWP40

MACRO IOA21D1BWP40
    CLASS CORE ;
    FOREIGN IOA21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.111250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.210 0.945 0.790 ;
        RECT  0.820 0.210 0.875 0.285 ;
        RECT  0.725 0.720 0.875 0.790 ;
        RECT  0.655 0.720 0.725 1.025 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.355 0.805 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.425 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.560 -0.115 0.980 0.115 ;
        RECT  0.440 -0.115 0.560 0.275 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.145 0.980 1.375 ;
        RECT  0.840 0.860 0.920 1.375 ;
        RECT  0.540 1.145 0.840 1.375 ;
        RECT  0.420 0.995 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.930 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.510 0.345 0.580 0.915 ;
        RECT  0.350 0.345 0.510 0.415 ;
        RECT  0.320 0.845 0.510 0.915 ;
        RECT  0.280 0.215 0.350 0.415 ;
        RECT  0.240 0.845 0.320 1.050 ;
        RECT  0.140 0.215 0.280 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA21D1BWP40

MACRO IOA21D2BWP40
    CLASS CORE ;
    FOREIGN IOA21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.223500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.075 0.760 1.145 1.025 ;
        RECT  0.805 0.855 1.075 0.925 ;
        RECT  0.805 0.335 0.955 0.405 ;
        RECT  0.735 0.335 0.805 0.925 ;
        RECT  0.695 0.855 0.735 0.925 ;
        RECT  0.625 0.855 0.695 1.025 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.995 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.450 0.405 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.635 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.280 -0.115 1.350 0.430 ;
        RECT  0.525 -0.115 1.280 0.115 ;
        RECT  0.410 -0.115 0.525 0.230 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.270 0.720 1.350 1.375 ;
        RECT  0.955 1.145 1.270 1.375 ;
        RECT  0.835 0.995 0.955 1.375 ;
        RECT  0.530 1.145 0.835 1.375 ;
        RECT  0.410 0.995 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.165 0.525 1.265 0.645 ;
        RECT  1.085 0.195 1.165 0.645 ;
        RECT  0.665 0.195 1.085 0.265 ;
        RECT  0.595 0.195 0.665 0.370 ;
        RECT  0.545 0.545 0.650 0.615 ;
        RECT  0.545 0.300 0.595 0.370 ;
        RECT  0.475 0.300 0.545 0.915 ;
        RECT  0.130 0.300 0.475 0.370 ;
        RECT  0.210 0.845 0.475 0.915 ;
        RECT  0.050 0.230 0.130 0.370 ;
    END
END IOA21D2BWP40

MACRO IOA21D4BWP40
    CLASS CORE ;
    FOREIGN IOA21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.375000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 0.355 2.415 1.075 ;
        RECT  2.205 0.355 2.340 0.915 ;
        RECT  1.940 0.355 2.205 0.425 ;
        RECT  2.040 0.845 2.205 0.915 ;
        RECT  1.960 0.845 2.040 1.075 ;
        RECT  1.660 0.845 1.960 0.915 ;
        RECT  1.580 0.750 1.660 1.010 ;
        RECT  1.280 0.845 1.580 0.915 ;
        RECT  1.200 0.750 1.280 1.010 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.495 2.105 0.625 ;
        RECT  1.845 0.495 1.925 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.300 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.760 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.655 -0.115 2.660 0.115 ;
        RECT  1.585 -0.115 1.655 0.285 ;
        RECT  1.275 -0.115 1.585 0.115 ;
        RECT  1.205 -0.115 1.275 0.285 ;
        RECT  0.345 -0.115 1.205 0.115 ;
        RECT  0.215 -0.115 0.345 0.220 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.145 2.660 1.375 ;
        RECT  2.530 0.720 2.605 1.375 ;
        RECT  2.230 1.145 2.530 1.375 ;
        RECT  2.150 0.985 2.230 1.375 ;
        RECT  1.850 1.145 2.150 1.375 ;
        RECT  1.770 0.985 1.850 1.375 ;
        RECT  1.470 1.145 1.770 1.375 ;
        RECT  1.390 0.985 1.470 1.375 ;
        RECT  1.090 1.145 1.390 1.375 ;
        RECT  1.015 0.795 1.090 1.375 ;
        RECT  0.715 1.145 1.015 1.375 ;
        RECT  0.605 0.900 0.715 1.375 ;
        RECT  0.335 1.145 0.605 1.375 ;
        RECT  0.225 0.900 0.335 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 0.355 2.135 0.425 ;
        RECT  2.040 0.845 2.135 0.915 ;
        RECT  1.960 0.845 2.040 1.075 ;
        RECT  1.660 0.845 1.960 0.915 ;
        RECT  1.580 0.750 1.660 1.010 ;
        RECT  1.280 0.845 1.580 0.915 ;
        RECT  1.200 0.750 1.280 1.010 ;
        RECT  2.535 0.205 2.605 0.490 ;
        RECT  1.845 0.205 2.535 0.275 ;
        RECT  1.775 0.205 1.845 0.425 ;
        RECT  1.465 0.355 1.775 0.425 ;
        RECT  0.935 0.545 1.660 0.615 ;
        RECT  1.395 0.190 1.465 0.425 ;
        RECT  1.085 0.355 1.395 0.425 ;
        RECT  1.015 0.250 1.085 0.425 ;
        RECT  0.885 0.345 0.935 0.830 ;
        RECT  0.505 0.195 0.910 0.265 ;
        RECT  0.865 0.345 0.885 1.020 ;
        RECT  0.595 0.345 0.865 0.415 ;
        RECT  0.815 0.760 0.865 1.020 ;
        RECT  0.505 0.760 0.815 0.830 ;
        RECT  0.430 0.195 0.505 0.370 ;
        RECT  0.435 0.760 0.505 1.020 ;
        RECT  0.125 0.760 0.435 0.830 ;
        RECT  0.035 0.290 0.430 0.370 ;
        RECT  0.055 0.760 0.125 1.020 ;
    END
END IOA21D4BWP40

MACRO IOA22D0BWP40
    CLASS CORE ;
    FOREIGN IOA22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.084725 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.845 1.365 1.045 ;
        RECT  0.720 0.845 1.260 0.945 ;
        RECT  0.705 0.185 0.720 0.945 ;
        RECT  0.650 0.185 0.705 1.055 ;
        RECT  0.615 0.185 0.650 0.450 ;
        RECT  0.595 0.775 0.650 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.235 0.495 1.365 0.650 ;
        RECT  1.155 0.495 1.235 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.495 1.085 0.635 ;
        RECT  0.875 0.495 0.955 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.765 ;
        RECT  0.250 0.695 0.315 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.120 0.285 ;
        RECT  0.510 -0.115 1.010 0.115 ;
        RECT  0.430 -0.115 0.510 0.270 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 1.400 1.375 ;
        RECT  0.810 1.015 0.910 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.975 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.935 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.185 1.360 0.425 ;
        RECT  0.900 0.355 1.260 0.425 ;
        RECT  0.800 0.195 0.900 0.425 ;
        RECT  0.545 0.520 0.580 0.640 ;
        RECT  0.525 0.340 0.545 0.640 ;
        RECT  0.455 0.340 0.525 0.905 ;
        RECT  0.310 0.340 0.455 0.410 ;
        RECT  0.320 0.835 0.455 0.905 ;
        RECT  0.240 0.835 0.320 1.055 ;
        RECT  0.240 0.215 0.310 0.410 ;
        RECT  0.140 0.215 0.240 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA22D0BWP40

MACRO IOA22D1BWP40
    CLASS CORE ;
    FOREIGN IOA22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.161750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.775 1.365 1.045 ;
        RECT  0.720 0.775 1.260 0.875 ;
        RECT  0.705 0.185 0.720 0.875 ;
        RECT  0.650 0.185 0.705 1.055 ;
        RECT  0.615 0.185 0.650 0.450 ;
        RECT  0.595 0.775 0.650 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.365 0.650 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.635 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.200 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.010 -0.115 1.120 0.285 ;
        RECT  0.510 -0.115 1.010 0.115 ;
        RECT  0.430 -0.115 0.510 0.285 ;
        RECT  0.000 -0.115 0.430 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 1.400 1.375 ;
        RECT  0.810 0.950 0.910 1.375 ;
        RECT  0.510 1.145 0.810 1.375 ;
        RECT  0.430 0.975 0.510 1.375 ;
        RECT  0.130 1.145 0.430 1.375 ;
        RECT  0.050 0.935 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.260 0.185 1.360 0.425 ;
        RECT  0.900 0.355 1.260 0.425 ;
        RECT  0.800 0.265 0.900 0.425 ;
        RECT  0.545 0.520 0.580 0.640 ;
        RECT  0.525 0.355 0.545 0.640 ;
        RECT  0.455 0.355 0.525 0.905 ;
        RECT  0.310 0.355 0.455 0.425 ;
        RECT  0.320 0.835 0.455 0.905 ;
        RECT  0.240 0.835 0.320 1.055 ;
        RECT  0.240 0.215 0.310 0.425 ;
        RECT  0.140 0.215 0.240 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END IOA22D1BWP40

MACRO IOA22D2BWP40
    CLASS CORE ;
    FOREIGN IOA22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.230950 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.835 1.925 1.065 ;
        RECT  1.065 0.835 1.805 0.905 ;
        RECT  0.995 0.835 1.065 1.065 ;
        RECT  0.945 0.835 0.995 0.905 ;
        RECT  0.875 0.345 0.945 0.905 ;
        RECT  0.775 0.345 0.875 0.430 ;
        RECT  0.695 0.835 0.875 0.905 ;
        RECT  0.615 0.835 0.695 0.975 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.810 0.765 ;
        RECT  1.225 0.695 1.715 0.765 ;
        RECT  1.115 0.495 1.225 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.635 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.635 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 -0.115 1.960 0.115 ;
        RECT  1.540 -0.115 1.670 0.210 ;
        RECT  1.260 -0.115 1.540 0.115 ;
        RECT  1.190 -0.115 1.260 0.240 ;
        RECT  0.130 -0.115 1.190 0.115 ;
        RECT  0.050 -0.115 0.130 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.145 1.960 1.375 ;
        RECT  1.350 1.115 1.480 1.375 ;
        RECT  0.900 1.145 1.350 1.375 ;
        RECT  0.780 1.025 0.900 1.375 ;
        RECT  0.530 1.145 0.780 1.375 ;
        RECT  0.410 0.990 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.850 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.805 0.185 1.900 0.415 ;
        RECT  1.450 0.345 1.805 0.415 ;
        RECT  1.155 0.975 1.675 1.045 ;
        RECT  1.380 0.185 1.450 0.415 ;
        RECT  1.095 0.345 1.380 0.415 ;
        RECT  1.025 0.195 1.095 0.415 ;
        RECT  0.685 0.195 1.025 0.265 ;
        RECT  0.545 0.540 0.795 0.620 ;
        RECT  0.615 0.195 0.685 0.350 ;
        RECT  0.475 0.210 0.545 0.890 ;
        RECT  0.410 0.210 0.475 0.280 ;
        RECT  0.320 0.820 0.475 0.890 ;
        RECT  0.240 0.820 0.320 1.075 ;
    END
END IOA22D2BWP40

MACRO IOA22D4BWP40
    CLASS CORE ;
    FOREIGN IOA22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.413250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.705 2.650 0.775 ;
        RECT  1.795 0.705 1.865 1.075 ;
        RECT  1.575 0.705 1.795 0.775 ;
        RECT  1.575 0.345 1.705 0.475 ;
        RECT  1.505 0.345 1.575 0.775 ;
        RECT  1.415 0.345 1.505 1.075 ;
        RECT  1.365 0.345 1.415 0.775 ;
        RECT  1.195 0.345 1.365 0.465 ;
        RECT  1.115 0.705 1.365 0.775 ;
        RECT  1.015 0.705 1.115 1.075 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.495 2.435 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.495 3.190 0.625 ;
        RECT  2.835 0.495 2.905 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.705 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 -0.115 3.640 0.115 ;
        RECT  3.285 -0.115 3.415 0.210 ;
        RECT  3.035 -0.115 3.285 0.115 ;
        RECT  2.905 -0.115 3.035 0.210 ;
        RECT  2.465 -0.115 2.905 0.115 ;
        RECT  2.345 -0.115 2.465 0.210 ;
        RECT  2.090 -0.115 2.345 0.115 ;
        RECT  1.960 -0.115 2.090 0.210 ;
        RECT  0.360 -0.115 1.960 0.115 ;
        RECT  0.280 -0.115 0.360 0.245 ;
        RECT  0.000 -0.115 0.280 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.145 3.640 1.375 ;
        RECT  3.290 1.035 3.415 1.375 ;
        RECT  3.035 1.145 3.290 1.375 ;
        RECT  2.905 1.035 3.035 1.375 ;
        RECT  1.705 1.145 2.905 1.375 ;
        RECT  1.575 0.910 1.705 1.375 ;
        RECT  1.320 1.145 1.575 1.375 ;
        RECT  1.200 0.910 1.320 1.375 ;
        RECT  0.765 1.145 1.200 1.375 ;
        RECT  0.640 0.990 0.765 1.375 ;
        RECT  0.360 1.145 0.640 1.375 ;
        RECT  0.280 0.985 0.360 1.375 ;
        RECT  0.000 1.145 0.280 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.865 0.705 2.650 0.775 ;
        RECT  1.795 0.705 1.865 1.075 ;
        RECT  1.645 0.705 1.795 0.775 ;
        RECT  1.645 0.345 1.705 0.475 ;
        RECT  1.195 0.345 1.295 0.465 ;
        RECT  1.115 0.705 1.295 0.775 ;
        RECT  1.015 0.705 1.115 1.075 ;
        RECT  3.505 0.185 3.595 0.415 ;
        RECT  3.505 0.685 3.575 1.075 ;
        RECT  3.195 0.345 3.505 0.415 ;
        RECT  3.195 0.845 3.505 0.915 ;
        RECT  3.125 0.185 3.195 0.415 ;
        RECT  3.125 0.845 3.195 1.075 ;
        RECT  2.810 0.345 3.125 0.415 ;
        RECT  2.815 0.845 3.125 0.915 ;
        RECT  2.745 0.845 2.815 1.075 ;
        RECT  2.740 0.185 2.810 0.415 ;
        RECT  2.440 0.845 2.745 0.915 ;
        RECT  2.630 0.345 2.740 0.415 ;
        RECT  2.560 0.185 2.630 0.415 ;
        RECT  2.250 0.345 2.560 0.415 ;
        RECT  2.370 0.845 2.440 1.075 ;
        RECT  2.060 0.845 2.370 0.915 ;
        RECT  2.180 0.185 2.250 0.415 ;
        RECT  1.870 0.345 2.180 0.415 ;
        RECT  1.970 0.845 2.060 1.075 ;
        RECT  1.800 0.195 1.870 0.415 ;
        RECT  1.105 0.195 1.800 0.265 ;
        RECT  0.925 0.545 1.275 0.625 ;
        RECT  1.035 0.195 1.105 0.450 ;
        RECT  0.545 0.195 0.955 0.265 ;
        RECT  0.855 0.335 0.925 1.075 ;
        RECT  0.850 0.335 0.855 0.915 ;
        RECT  0.635 0.335 0.850 0.405 ;
        RECT  0.545 0.845 0.850 0.915 ;
        RECT  0.475 0.195 0.545 0.425 ;
        RECT  0.475 0.845 0.545 1.075 ;
        RECT  0.165 0.355 0.475 0.425 ;
        RECT  0.160 0.845 0.475 0.915 ;
        RECT  0.075 0.195 0.165 0.425 ;
        RECT  0.070 0.845 0.160 1.075 ;
    END
END IOA22D4BWP40

MACRO LHCNQD0BWP40
    CLASS CORE ;
    FOREIGN LHCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.670 0.185 2.765 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 1.120 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.020800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.345 1.825 0.485 ;
        RECT  0.785 0.345 1.575 0.415 ;
        RECT  0.705 0.345 0.785 0.615 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.535 -0.115 2.800 0.115 ;
        RECT  2.455 -0.115 2.535 0.280 ;
        RECT  1.950 -0.115 2.455 0.115 ;
        RECT  1.820 -0.115 1.950 0.135 ;
        RECT  0.830 -0.115 1.820 0.115 ;
        RECT  0.720 -0.115 0.830 0.265 ;
        RECT  0.385 -0.115 0.720 0.115 ;
        RECT  0.275 -0.115 0.385 0.235 ;
        RECT  0.000 -0.115 0.275 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.540 1.145 2.800 1.375 ;
        RECT  2.460 0.945 2.540 1.375 ;
        RECT  1.940 1.145 2.460 1.375 ;
        RECT  1.820 1.140 1.940 1.375 ;
        RECT  1.050 1.145 1.820 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.350 1.145 0.930 1.375 ;
        RECT  0.260 0.980 0.350 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.520 0.405 2.590 0.760 ;
        RECT  2.330 0.405 2.520 0.475 ;
        RECT  2.330 0.690 2.520 0.760 ;
        RECT  2.135 0.545 2.410 0.620 ;
        RECT  2.250 0.185 2.330 0.475 ;
        RECT  2.250 0.690 2.330 1.050 ;
        RECT  2.055 0.185 2.135 1.060 ;
        RECT  1.790 0.990 2.055 1.060 ;
        RECT  1.905 0.205 1.975 0.920 ;
        RECT  1.275 0.205 1.905 0.275 ;
        RECT  0.730 0.850 1.905 0.920 ;
        RECT  1.650 0.990 1.790 1.075 ;
        RECT  1.260 0.705 1.670 0.780 ;
        RECT  1.270 0.990 1.440 1.075 ;
        RECT  1.260 0.490 1.310 0.580 ;
        RECT  0.490 0.990 1.270 1.060 ;
        RECT  1.190 0.490 1.260 0.780 ;
        RECT  0.650 0.695 1.190 0.780 ;
        RECT  0.630 0.695 0.650 0.920 ;
        RECT  0.560 0.185 0.630 0.920 ;
        RECT  0.420 0.305 0.490 1.060 ;
        RECT  0.380 0.305 0.420 0.910 ;
        RECT  0.190 0.305 0.380 0.375 ;
        RECT  0.175 0.840 0.380 0.910 ;
        RECT  0.070 0.210 0.190 0.375 ;
        RECT  0.090 0.840 0.175 1.040 ;
    END
END LHCNQD0BWP40

MACRO LHCNQD1BWP40
    CLASS CORE ;
    FOREIGN LHCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.670 0.185 2.765 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.035 0.495 0.175 0.630 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 1.120 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.345 1.825 0.625 ;
        RECT  0.785 0.345 1.715 0.415 ;
        RECT  0.705 0.345 0.785 0.615 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 -0.115 2.800 0.115 ;
        RECT  2.480 -0.115 2.560 0.335 ;
        RECT  1.950 -0.115 2.480 0.115 ;
        RECT  1.820 -0.115 1.950 0.135 ;
        RECT  0.835 -0.115 1.820 0.115 ;
        RECT  0.725 -0.115 0.835 0.265 ;
        RECT  0.385 -0.115 0.725 0.115 ;
        RECT  0.275 -0.115 0.385 0.235 ;
        RECT  0.000 -0.115 0.275 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.145 2.800 1.375 ;
        RECT  2.480 0.830 2.560 1.375 ;
        RECT  1.940 1.145 2.480 1.375 ;
        RECT  1.820 1.140 1.940 1.375 ;
        RECT  1.050 1.145 1.820 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.350 1.145 0.930 1.375 ;
        RECT  0.260 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.520 0.405 2.590 0.760 ;
        RECT  2.330 0.405 2.520 0.475 ;
        RECT  2.330 0.690 2.520 0.760 ;
        RECT  2.135 0.545 2.410 0.620 ;
        RECT  2.230 0.185 2.330 0.475 ;
        RECT  2.250 0.690 2.330 1.040 ;
        RECT  2.055 0.185 2.135 1.060 ;
        RECT  1.790 0.990 2.055 1.060 ;
        RECT  1.905 0.205 1.975 0.920 ;
        RECT  1.275 0.205 1.905 0.275 ;
        RECT  0.730 0.850 1.905 0.920 ;
        RECT  1.650 0.990 1.790 1.075 ;
        RECT  1.310 0.705 1.670 0.780 ;
        RECT  1.270 0.990 1.440 1.075 ;
        RECT  1.190 0.490 1.310 0.780 ;
        RECT  0.490 0.990 1.270 1.060 ;
        RECT  0.650 0.695 1.190 0.780 ;
        RECT  0.630 0.695 0.650 0.920 ;
        RECT  0.560 0.185 0.630 0.920 ;
        RECT  0.420 0.305 0.490 1.060 ;
        RECT  0.380 0.305 0.420 0.905 ;
        RECT  0.190 0.305 0.380 0.375 ;
        RECT  0.180 0.835 0.380 0.905 ;
        RECT  0.070 0.210 0.190 0.375 ;
        RECT  0.070 0.835 0.180 1.020 ;
    END
END LHCNQD1BWP40

MACRO LHCNQD2BWP40
    CLASS CORE ;
    FOREIGN LHCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.775 ;
        RECT  2.615 0.185 2.695 0.455 ;
        RECT  2.615 0.705 2.695 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 1.120 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.345 1.825 0.625 ;
        RECT  0.785 0.345 1.715 0.415 ;
        RECT  0.705 0.345 0.785 0.615 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.115 2.940 0.115 ;
        RECT  2.805 -0.115 2.885 0.290 ;
        RECT  2.500 -0.115 2.805 0.115 ;
        RECT  2.420 -0.115 2.500 0.325 ;
        RECT  1.950 -0.115 2.420 0.115 ;
        RECT  1.820 -0.115 1.950 0.135 ;
        RECT  0.835 -0.115 1.820 0.115 ;
        RECT  0.725 -0.115 0.835 0.275 ;
        RECT  0.385 -0.115 0.725 0.115 ;
        RECT  0.275 -0.115 0.385 0.235 ;
        RECT  0.000 -0.115 0.275 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.830 2.890 1.375 ;
        RECT  2.500 1.145 2.810 1.375 ;
        RECT  2.420 0.830 2.500 1.375 ;
        RECT  1.940 1.145 2.420 1.375 ;
        RECT  1.820 1.140 1.940 1.375 ;
        RECT  1.050 1.145 1.820 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.350 1.145 0.930 1.375 ;
        RECT  0.260 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.545 0.525 2.625 0.635 ;
        RECT  2.475 0.405 2.545 0.760 ;
        RECT  2.310 0.405 2.475 0.475 ;
        RECT  2.310 0.690 2.475 0.760 ;
        RECT  2.135 0.545 2.395 0.620 ;
        RECT  2.235 0.185 2.310 0.475 ;
        RECT  2.230 0.690 2.310 1.040 ;
        RECT  2.055 0.185 2.135 1.060 ;
        RECT  1.790 0.990 2.055 1.060 ;
        RECT  1.905 0.205 1.975 0.920 ;
        RECT  1.275 0.205 1.905 0.275 ;
        RECT  0.730 0.850 1.905 0.920 ;
        RECT  1.650 0.990 1.790 1.075 ;
        RECT  1.310 0.705 1.670 0.780 ;
        RECT  1.270 0.990 1.440 1.075 ;
        RECT  1.190 0.490 1.310 0.780 ;
        RECT  0.490 0.990 1.270 1.060 ;
        RECT  0.650 0.695 1.190 0.780 ;
        RECT  0.630 0.695 0.650 0.920 ;
        RECT  0.560 0.185 0.630 0.920 ;
        RECT  0.420 0.305 0.490 1.060 ;
        RECT  0.380 0.305 0.420 0.905 ;
        RECT  0.190 0.305 0.380 0.375 ;
        RECT  0.180 0.835 0.380 0.905 ;
        RECT  0.070 0.210 0.190 0.375 ;
        RECT  0.070 0.835 0.180 1.020 ;
    END
END LHCNQD2BWP40

MACRO LHCNQD4BWP40
    CLASS CORE ;
    FOREIGN LHCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 0.185 3.260 0.460 ;
        RECT  3.180 0.755 3.260 1.050 ;
        RECT  3.115 0.350 3.180 0.460 ;
        RECT  3.115 0.755 3.180 0.905 ;
        RECT  2.905 0.350 3.115 0.905 ;
        RECT  2.890 0.350 2.905 0.460 ;
        RECT  2.885 0.755 2.905 0.905 ;
        RECT  2.805 0.185 2.890 0.460 ;
        RECT  2.805 0.755 2.885 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 1.120 0.625 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.345 1.825 0.625 ;
        RECT  0.785 0.345 1.715 0.415 ;
        RECT  0.705 0.345 0.785 0.615 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.115 3.500 0.115 ;
        RECT  3.365 -0.115 3.445 0.430 ;
        RECT  3.070 -0.115 3.365 0.115 ;
        RECT  2.990 -0.115 3.070 0.275 ;
        RECT  2.690 -0.115 2.990 0.115 ;
        RECT  2.610 -0.115 2.690 0.450 ;
        RECT  2.310 -0.115 2.610 0.115 ;
        RECT  2.235 -0.115 2.310 0.435 ;
        RECT  1.950 -0.115 2.235 0.115 ;
        RECT  1.820 -0.115 1.950 0.135 ;
        RECT  0.830 -0.115 1.820 0.115 ;
        RECT  0.720 -0.115 0.830 0.265 ;
        RECT  0.385 -0.115 0.720 0.115 ;
        RECT  0.275 -0.115 0.385 0.235 ;
        RECT  0.000 -0.115 0.275 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.715 3.450 1.375 ;
        RECT  3.070 1.145 3.370 1.375 ;
        RECT  2.990 1.000 3.070 1.375 ;
        RECT  2.690 1.145 2.990 1.375 ;
        RECT  2.610 0.720 2.690 1.375 ;
        RECT  2.310 1.145 2.610 1.375 ;
        RECT  2.235 0.720 2.310 1.375 ;
        RECT  1.940 1.145 2.235 1.375 ;
        RECT  1.820 1.140 1.940 1.375 ;
        RECT  1.050 1.145 1.820 1.375 ;
        RECT  0.930 1.130 1.050 1.375 ;
        RECT  0.350 1.145 0.930 1.375 ;
        RECT  0.260 0.985 0.350 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.185 3.260 0.460 ;
        RECT  3.185 0.755 3.260 1.050 ;
        RECT  2.805 0.185 2.835 0.460 ;
        RECT  2.805 0.755 2.835 1.050 ;
        RECT  2.500 0.550 2.830 0.620 ;
        RECT  2.425 0.185 2.500 1.040 ;
        RECT  2.135 0.545 2.310 0.620 ;
        RECT  2.055 0.185 2.135 1.060 ;
        RECT  1.790 0.990 2.055 1.060 ;
        RECT  1.905 0.205 1.975 0.920 ;
        RECT  1.275 0.205 1.905 0.275 ;
        RECT  0.730 0.850 1.905 0.920 ;
        RECT  1.650 0.990 1.790 1.075 ;
        RECT  1.260 0.705 1.670 0.780 ;
        RECT  1.270 0.990 1.440 1.075 ;
        RECT  1.260 0.490 1.375 0.580 ;
        RECT  0.490 0.990 1.270 1.060 ;
        RECT  1.190 0.490 1.260 0.780 ;
        RECT  0.650 0.695 1.190 0.780 ;
        RECT  0.630 0.695 0.650 0.920 ;
        RECT  0.560 0.185 0.630 0.920 ;
        RECT  0.420 0.305 0.490 1.060 ;
        RECT  0.380 0.305 0.420 0.905 ;
        RECT  0.190 0.305 0.380 0.375 ;
        RECT  0.170 0.835 0.380 0.905 ;
        RECT  0.070 0.210 0.190 0.375 ;
        RECT  0.085 0.835 0.170 1.020 ;
    END
END LHCNQD4BWP40

MACRO LHCSNQD0BWP40
    CLASS CORE ;
    FOREIGN LHCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.620 1.590 0.765 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.185 3.185 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.630 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.995 0.495 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.365 0.635 2.495 0.930 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 -0.115 3.220 0.115 ;
        RECT  2.880 -0.115 3.000 0.210 ;
        RECT  2.580 -0.115 2.880 0.115 ;
        RECT  2.455 -0.115 2.580 0.125 ;
        RECT  1.505 -0.115 2.455 0.115 ;
        RECT  1.425 -0.115 1.505 0.260 ;
        RECT  0.710 -0.115 1.425 0.115 ;
        RECT  0.630 -0.115 0.710 0.275 ;
        RECT  0.330 -0.115 0.630 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 1.145 3.220 1.375 ;
        RECT  2.900 0.900 2.980 1.375 ;
        RECT  2.590 1.145 2.900 1.375 ;
        RECT  2.490 1.005 2.590 1.375 ;
        RECT  2.090 1.145 2.490 1.375 ;
        RECT  2.015 0.895 2.090 1.375 ;
        RECT  1.485 1.145 2.015 1.375 ;
        RECT  1.365 1.135 1.485 1.375 ;
        RECT  0.725 1.145 1.365 1.375 ;
        RECT  0.605 0.960 0.725 1.375 ;
        RECT  0.330 1.145 0.605 1.375 ;
        RECT  0.245 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.280 3.020 0.795 ;
        RECT  2.755 0.280 2.950 0.350 ;
        RECT  2.760 0.720 2.950 0.795 ;
        RECT  2.755 0.490 2.840 0.640 ;
        RECT  2.685 0.720 2.760 1.065 ;
        RECT  2.685 0.185 2.755 0.350 ;
        RECT  2.575 0.490 2.755 0.565 ;
        RECT  2.505 0.215 2.575 0.565 ;
        RECT  2.250 0.215 2.505 0.285 ;
        RECT  2.320 0.355 2.410 0.565 ;
        RECT  2.240 1.005 2.410 1.075 ;
        RECT  2.240 0.495 2.320 0.565 ;
        RECT  2.180 0.215 2.250 0.415 ;
        RECT  2.170 0.495 2.240 1.075 ;
        RECT  1.915 0.345 2.180 0.415 ;
        RECT  2.005 0.495 2.170 0.640 ;
        RECT  1.605 0.195 2.110 0.265 ;
        RECT  1.835 0.345 1.915 1.065 ;
        RECT  1.240 0.995 1.835 1.065 ;
        RECT  1.755 0.520 1.765 0.645 ;
        RECT  1.680 0.345 1.755 0.915 ;
        RECT  1.350 0.345 1.680 0.415 ;
        RECT  1.085 0.845 1.680 0.915 ;
        RECT  1.270 0.205 1.350 0.415 ;
        RECT  0.950 0.205 1.270 0.275 ;
        RECT  1.145 0.465 1.215 0.635 ;
        RECT  0.905 0.705 1.215 0.775 ;
        RECT  0.765 0.565 1.145 0.635 ;
        RECT  0.985 0.845 1.085 0.990 ;
        RECT  0.835 0.705 0.905 0.890 ;
        RECT  0.535 0.815 0.835 0.890 ;
        RECT  0.695 0.565 0.765 0.730 ;
        RECT  0.535 0.425 0.660 0.500 ;
        RECT  0.455 0.195 0.535 0.890 ;
        RECT  0.315 0.330 0.385 0.920 ;
        RECT  0.135 0.330 0.315 0.400 ;
        RECT  0.135 0.845 0.315 0.920 ;
        RECT  0.050 0.205 0.135 0.400 ;
        RECT  0.045 0.845 0.135 1.050 ;
    END
END LHCSNQD0BWP40

MACRO LHCSNQD1BWP40
    CLASS CORE ;
    FOREIGN LHCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.620 1.590 0.765 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.095 0.185 3.185 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.630 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.995 0.495 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.022800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.365 0.635 2.495 0.930 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.000 -0.115 3.220 0.115 ;
        RECT  2.875 -0.115 3.000 0.260 ;
        RECT  2.580 -0.115 2.875 0.115 ;
        RECT  2.455 -0.115 2.580 0.125 ;
        RECT  1.505 -0.115 2.455 0.115 ;
        RECT  1.425 -0.115 1.505 0.260 ;
        RECT  0.710 -0.115 1.425 0.115 ;
        RECT  0.630 -0.115 0.710 0.260 ;
        RECT  0.330 -0.115 0.630 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 1.145 3.220 1.375 ;
        RECT  2.900 0.870 2.980 1.375 ;
        RECT  2.590 1.145 2.900 1.375 ;
        RECT  2.490 1.005 2.590 1.375 ;
        RECT  2.090 1.145 2.490 1.375 ;
        RECT  2.015 0.815 2.090 1.375 ;
        RECT  1.485 1.145 2.015 1.375 ;
        RECT  1.365 1.135 1.485 1.375 ;
        RECT  0.725 1.145 1.365 1.375 ;
        RECT  0.605 0.975 0.725 1.375 ;
        RECT  0.330 1.145 0.605 1.375 ;
        RECT  0.245 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.340 3.020 0.795 ;
        RECT  2.760 0.340 2.950 0.410 ;
        RECT  2.760 0.720 2.950 0.795 ;
        RECT  2.755 0.490 2.840 0.640 ;
        RECT  2.685 0.270 2.760 0.410 ;
        RECT  2.685 0.720 2.760 1.030 ;
        RECT  2.575 0.490 2.755 0.565 ;
        RECT  2.505 0.215 2.575 0.565 ;
        RECT  2.250 0.215 2.505 0.285 ;
        RECT  2.320 0.370 2.410 0.565 ;
        RECT  2.240 1.005 2.410 1.075 ;
        RECT  2.240 0.495 2.320 0.565 ;
        RECT  2.180 0.215 2.250 0.415 ;
        RECT  2.170 0.495 2.240 1.075 ;
        RECT  1.915 0.345 2.180 0.415 ;
        RECT  2.005 0.495 2.170 0.640 ;
        RECT  1.605 0.195 2.110 0.265 ;
        RECT  1.835 0.345 1.915 1.065 ;
        RECT  1.240 0.995 1.835 1.065 ;
        RECT  1.755 0.520 1.765 0.645 ;
        RECT  1.680 0.345 1.755 0.915 ;
        RECT  1.350 0.345 1.680 0.415 ;
        RECT  1.085 0.845 1.680 0.915 ;
        RECT  1.270 0.205 1.350 0.415 ;
        RECT  0.950 0.205 1.270 0.275 ;
        RECT  1.145 0.465 1.215 0.635 ;
        RECT  0.905 0.705 1.215 0.775 ;
        RECT  0.765 0.565 1.145 0.635 ;
        RECT  0.985 0.845 1.085 1.005 ;
        RECT  0.835 0.705 0.905 0.895 ;
        RECT  0.535 0.820 0.835 0.895 ;
        RECT  0.695 0.565 0.765 0.730 ;
        RECT  0.535 0.425 0.660 0.500 ;
        RECT  0.455 0.195 0.535 0.895 ;
        RECT  0.315 0.330 0.385 0.920 ;
        RECT  0.135 0.330 0.315 0.400 ;
        RECT  0.135 0.845 0.315 0.920 ;
        RECT  0.050 0.205 0.135 0.400 ;
        RECT  0.045 0.845 0.135 1.050 ;
    END
END LHCSNQD1BWP40

MACRO LHCSNQD2BWP40
    CLASS CORE ;
    FOREIGN LHCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.635 1.585 0.765 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.355 3.185 0.775 ;
        RECT  3.025 0.185 3.115 0.455 ;
        RECT  3.025 0.705 3.115 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.990 0.495 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.022800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.635 2.515 0.905 ;
        RECT  2.340 0.650 2.415 0.905 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.310 0.300 ;
        RECT  2.950 -0.115 3.230 0.115 ;
        RECT  2.835 -0.115 2.950 0.235 ;
        RECT  2.560 -0.115 2.835 0.115 ;
        RECT  2.435 -0.115 2.560 0.125 ;
        RECT  1.500 -0.115 2.435 0.115 ;
        RECT  1.420 -0.115 1.500 0.260 ;
        RECT  0.715 -0.115 1.420 0.115 ;
        RECT  0.635 -0.115 0.715 0.260 ;
        RECT  0.330 -0.115 0.635 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.315 1.145 3.360 1.375 ;
        RECT  3.230 0.840 3.315 1.375 ;
        RECT  2.930 1.145 3.230 1.375 ;
        RECT  2.850 0.870 2.930 1.375 ;
        RECT  2.570 1.145 2.850 1.375 ;
        RECT  2.470 1.005 2.570 1.375 ;
        RECT  2.085 1.145 2.470 1.375 ;
        RECT  2.015 0.810 2.085 1.375 ;
        RECT  1.480 1.145 2.015 1.375 ;
        RECT  1.360 1.135 1.480 1.375 ;
        RECT  0.730 1.145 1.360 1.375 ;
        RECT  0.610 0.995 0.730 1.375 ;
        RECT  0.330 1.145 0.610 1.375 ;
        RECT  0.245 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.945 0.525 3.045 0.635 ;
        RECT  2.875 0.305 2.945 0.795 ;
        RECT  2.645 0.305 2.875 0.375 ;
        RECT  2.745 0.720 2.875 0.795 ;
        RECT  2.735 0.490 2.805 0.640 ;
        RECT  2.670 0.720 2.745 1.030 ;
        RECT  2.555 0.490 2.735 0.565 ;
        RECT  2.485 0.215 2.555 0.565 ;
        RECT  2.230 0.215 2.485 0.285 ;
        RECT  2.235 1.005 2.390 1.075 ;
        RECT  2.300 0.365 2.370 0.580 ;
        RECT  2.235 0.510 2.300 0.580 ;
        RECT  2.165 0.510 2.235 1.075 ;
        RECT  2.160 0.215 2.230 0.435 ;
        RECT  2.055 0.510 2.165 0.635 ;
        RECT  1.935 0.365 2.160 0.435 ;
        RECT  2.000 0.185 2.080 0.295 ;
        RECT  1.590 0.195 2.000 0.265 ;
        RECT  1.855 0.365 1.935 1.065 ;
        RECT  1.815 0.365 1.855 0.480 ;
        RECT  1.245 0.995 1.855 1.065 ;
        RECT  1.745 0.545 1.785 0.625 ;
        RECT  1.675 0.345 1.745 0.915 ;
        RECT  1.345 0.345 1.675 0.415 ;
        RECT  1.075 0.845 1.675 0.915 ;
        RECT  1.265 0.205 1.345 0.415 ;
        RECT  0.955 0.205 1.265 0.275 ;
        RECT  1.140 0.465 1.210 0.635 ;
        RECT  0.910 0.705 1.210 0.775 ;
        RECT  0.770 0.565 1.140 0.635 ;
        RECT  1.005 0.845 1.075 0.955 ;
        RECT  0.840 0.705 0.910 0.895 ;
        RECT  0.540 0.820 0.840 0.895 ;
        RECT  0.700 0.565 0.770 0.730 ;
        RECT  0.540 0.425 0.665 0.500 ;
        RECT  0.460 0.195 0.540 0.895 ;
        RECT  0.315 0.330 0.385 0.920 ;
        RECT  0.135 0.330 0.315 0.400 ;
        RECT  0.135 0.845 0.315 0.920 ;
        RECT  0.050 0.205 0.135 0.400 ;
        RECT  0.045 0.845 0.135 1.050 ;
    END
END LHCSNQD2BWP40

MACRO LHCSNQD4BWP40
    CLASS CORE ;
    FOREIGN LHCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.620 1.590 0.765 ;
        RECT  1.435 0.495 1.505 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.460 0.185 3.540 0.460 ;
        RECT  3.460 0.755 3.540 1.050 ;
        RECT  3.395 0.350 3.460 0.460 ;
        RECT  3.395 0.755 3.460 0.905 ;
        RECT  3.185 0.350 3.395 0.905 ;
        RECT  3.170 0.350 3.185 0.460 ;
        RECT  3.165 0.755 3.185 0.905 ;
        RECT  3.085 0.185 3.170 0.460 ;
        RECT  3.085 0.755 3.165 1.050 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.635 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.024000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.995 0.495 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.022800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.475 0.775 2.625 0.905 ;
        RECT  2.365 0.635 2.475 0.905 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.115 3.780 0.115 ;
        RECT  3.645 -0.115 3.725 0.440 ;
        RECT  3.350 -0.115 3.645 0.115 ;
        RECT  3.270 -0.115 3.350 0.275 ;
        RECT  2.970 -0.115 3.270 0.115 ;
        RECT  2.890 -0.115 2.970 0.265 ;
        RECT  1.505 -0.115 2.890 0.115 ;
        RECT  1.425 -0.115 1.505 0.260 ;
        RECT  0.710 -0.115 1.425 0.115 ;
        RECT  0.630 -0.115 0.710 0.260 ;
        RECT  0.330 -0.115 0.630 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.715 3.730 1.375 ;
        RECT  3.350 1.145 3.650 1.375 ;
        RECT  3.270 1.000 3.350 1.375 ;
        RECT  2.975 1.145 3.270 1.375 ;
        RECT  2.885 0.885 2.975 1.375 ;
        RECT  2.590 1.145 2.885 1.375 ;
        RECT  2.490 1.005 2.590 1.375 ;
        RECT  2.085 1.145 2.490 1.375 ;
        RECT  2.010 0.805 2.085 1.375 ;
        RECT  1.485 1.145 2.010 1.375 ;
        RECT  1.365 1.135 1.485 1.375 ;
        RECT  0.725 1.145 1.365 1.375 ;
        RECT  0.605 0.995 0.725 1.375 ;
        RECT  0.330 1.145 0.605 1.375 ;
        RECT  0.245 0.990 0.330 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.185 3.540 0.460 ;
        RECT  3.465 0.755 3.540 1.050 ;
        RECT  3.085 0.185 3.115 0.460 ;
        RECT  3.085 0.755 3.115 1.050 ;
        RECT  2.955 0.550 3.110 0.620 ;
        RECT  2.885 0.400 2.955 0.815 ;
        RECT  2.785 0.400 2.885 0.470 ;
        RECT  2.780 0.745 2.885 0.815 ;
        RECT  2.710 0.185 2.785 0.470 ;
        RECT  2.630 0.540 2.785 0.610 ;
        RECT  2.705 0.745 2.780 1.040 ;
        RECT  2.560 0.250 2.630 0.610 ;
        RECT  2.250 0.250 2.560 0.320 ;
        RECT  2.320 0.390 2.410 0.565 ;
        RECT  2.235 1.005 2.410 1.075 ;
        RECT  2.235 0.495 2.320 0.565 ;
        RECT  2.180 0.250 2.250 0.415 ;
        RECT  2.165 0.495 2.235 1.075 ;
        RECT  1.915 0.345 2.180 0.415 ;
        RECT  2.145 0.495 2.165 0.640 ;
        RECT  1.595 0.195 2.110 0.265 ;
        RECT  1.835 0.345 1.915 1.065 ;
        RECT  1.240 0.995 1.835 1.065 ;
        RECT  1.755 0.520 1.765 0.645 ;
        RECT  1.680 0.345 1.755 0.915 ;
        RECT  1.350 0.345 1.680 0.415 ;
        RECT  1.085 0.845 1.680 0.915 ;
        RECT  1.270 0.205 1.350 0.415 ;
        RECT  0.950 0.205 1.270 0.275 ;
        RECT  1.145 0.465 1.215 0.635 ;
        RECT  0.905 0.705 1.215 0.775 ;
        RECT  0.765 0.565 1.145 0.635 ;
        RECT  0.985 0.845 1.085 1.005 ;
        RECT  0.835 0.705 0.905 0.895 ;
        RECT  0.535 0.820 0.835 0.895 ;
        RECT  0.695 0.565 0.765 0.730 ;
        RECT  0.535 0.425 0.660 0.500 ;
        RECT  0.455 0.195 0.535 0.895 ;
        RECT  0.315 0.330 0.385 0.920 ;
        RECT  0.135 0.330 0.315 0.400 ;
        RECT  0.135 0.845 0.315 0.920 ;
        RECT  0.050 0.205 0.135 0.400 ;
        RECT  0.045 0.845 0.135 1.050 ;
    END
END LHCSNQD4BWP40

MACRO LHQD0BWP40
    CLASS CORE ;
    FOREIGN LHQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 0.935 ;
        RECT  1.835 0.185 1.855 0.305 ;
        RECT  1.835 0.825 1.855 0.935 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 0.570 1.785 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.115 1.960 0.115 ;
        RECT  1.650 -0.115 1.720 0.260 ;
        RECT  0.885 -0.115 1.650 0.115 ;
        RECT  0.805 -0.115 0.885 0.280 ;
        RECT  0.345 -0.115 0.805 0.115 ;
        RECT  0.215 -0.115 0.345 0.190 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.145 1.960 1.375 ;
        RECT  1.620 0.845 1.720 1.375 ;
        RECT  0.910 1.145 1.620 1.375 ;
        RECT  0.800 1.000 0.910 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 0.390 1.785 0.500 ;
        RECT  1.510 0.210 1.580 0.500 ;
        RECT  1.265 0.210 1.510 0.290 ;
        RECT  1.335 0.370 1.405 1.065 ;
        RECT  1.050 0.995 1.335 1.065 ;
        RECT  1.190 0.210 1.265 0.895 ;
        RECT  1.180 0.210 1.190 0.440 ;
        RECT  0.850 0.370 1.180 0.440 ;
        RECT  0.980 0.860 1.050 1.065 ;
        RECT  0.935 0.510 1.025 0.790 ;
        RECT  0.525 0.860 0.980 0.930 ;
        RECT  0.685 0.720 0.935 0.790 ;
        RECT  0.765 0.370 0.850 0.640 ;
        RECT  0.615 0.185 0.685 0.790 ;
        RECT  0.450 0.285 0.525 1.005 ;
        RECT  0.420 0.285 0.450 0.385 ;
        RECT  0.430 0.860 0.450 1.005 ;
        RECT  0.340 0.550 0.380 0.670 ;
        RECT  0.270 0.260 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD0BWP40

MACRO LHQD1BWP40
    CLASS CORE ;
    FOREIGN LHQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.090850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 1.045 ;
        RECT  1.835 0.185 1.855 0.305 ;
        RECT  1.835 0.695 1.855 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 0.495 1.645 0.770 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.115 1.960 0.115 ;
        RECT  1.650 -0.115 1.720 0.260 ;
        RECT  0.885 -0.115 1.650 0.115 ;
        RECT  0.805 -0.115 0.885 0.280 ;
        RECT  0.340 -0.115 0.805 0.115 ;
        RECT  0.220 -0.115 0.340 0.190 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.145 1.960 1.375 ;
        RECT  1.620 0.845 1.720 1.375 ;
        RECT  0.910 1.145 1.620 1.375 ;
        RECT  0.800 1.000 0.910 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.580 0.355 1.715 0.425 ;
        RECT  1.510 0.210 1.580 0.425 ;
        RECT  1.245 0.210 1.510 0.290 ;
        RECT  1.370 0.370 1.440 1.065 ;
        RECT  1.315 0.370 1.370 0.500 ;
        RECT  1.050 0.995 1.370 1.065 ;
        RECT  1.245 0.780 1.290 0.895 ;
        RECT  1.170 0.210 1.245 0.895 ;
        RECT  0.850 0.370 1.170 0.440 ;
        RECT  0.980 0.860 1.050 1.065 ;
        RECT  0.935 0.510 1.025 0.790 ;
        RECT  0.525 0.860 0.980 0.930 ;
        RECT  0.685 0.720 0.935 0.790 ;
        RECT  0.765 0.370 0.850 0.640 ;
        RECT  0.615 0.185 0.685 0.790 ;
        RECT  0.450 0.285 0.525 1.005 ;
        RECT  0.420 0.285 0.450 0.385 ;
        RECT  0.430 0.860 0.450 1.005 ;
        RECT  0.340 0.550 0.380 0.670 ;
        RECT  0.270 0.260 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD1BWP40

MACRO LHQD2BWP40
    CLASS CORE ;
    FOREIGN LHQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.116250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.355 1.925 0.765 ;
        RECT  1.855 0.185 1.875 1.045 ;
        RECT  1.790 0.185 1.855 0.425 ;
        RECT  1.785 0.695 1.855 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.031000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.665 1.715 0.905 ;
        RECT  1.480 0.505 1.560 0.905 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.975 -0.115 2.050 0.305 ;
        RECT  1.670 -0.115 1.975 0.115 ;
        RECT  1.600 -0.115 1.670 0.260 ;
        RECT  0.885 -0.115 1.600 0.115 ;
        RECT  0.805 -0.115 0.885 0.280 ;
        RECT  0.340 -0.115 0.805 0.115 ;
        RECT  0.215 -0.115 0.340 0.190 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.835 2.050 1.375 ;
        RECT  1.670 1.145 1.970 1.375 ;
        RECT  1.570 1.000 1.670 1.375 ;
        RECT  0.910 1.145 1.570 1.375 ;
        RECT  0.800 1.000 0.910 1.375 ;
        RECT  0.340 1.145 0.800 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 0.525 1.760 0.595 ;
        RECT  1.630 0.340 1.720 0.595 ;
        RECT  1.530 0.340 1.630 0.410 ;
        RECT  1.460 0.210 1.530 0.410 ;
        RECT  1.205 0.210 1.460 0.290 ;
        RECT  1.370 0.500 1.405 1.065 ;
        RECT  1.335 0.375 1.370 1.065 ;
        RECT  1.285 0.375 1.335 0.565 ;
        RECT  1.050 0.995 1.335 1.065 ;
        RECT  1.205 0.795 1.265 0.915 ;
        RECT  1.130 0.210 1.205 0.915 ;
        RECT  0.850 0.370 1.130 0.440 ;
        RECT  0.980 0.860 1.050 1.065 ;
        RECT  0.935 0.520 1.025 0.790 ;
        RECT  0.525 0.860 0.980 0.930 ;
        RECT  0.685 0.720 0.935 0.790 ;
        RECT  0.765 0.370 0.850 0.640 ;
        RECT  0.615 0.185 0.685 0.790 ;
        RECT  0.450 0.285 0.525 1.005 ;
        RECT  0.420 0.285 0.450 0.385 ;
        RECT  0.430 0.860 0.450 1.005 ;
        RECT  0.340 0.550 0.380 0.670 ;
        RECT  0.270 0.260 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD2BWP40

MACRO LHQD4BWP40
    CLASS CORE ;
    FOREIGN LHQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.237000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.185 2.980 0.480 ;
        RECT  2.900 0.755 2.980 1.035 ;
        RECT  2.835 0.350 2.900 0.480 ;
        RECT  2.835 0.755 2.900 0.910 ;
        RECT  2.625 0.350 2.835 0.910 ;
        RECT  2.600 0.350 2.625 0.480 ;
        RECT  2.600 0.755 2.625 0.910 ;
        RECT  2.525 0.185 2.600 0.480 ;
        RECT  2.525 0.755 2.600 1.040 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.205 0.625 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.170 0.460 ;
        RECT  2.795 -0.115 3.095 0.115 ;
        RECT  2.715 -0.115 2.795 0.275 ;
        RECT  2.405 -0.115 2.715 0.115 ;
        RECT  2.335 -0.115 2.405 0.255 ;
        RECT  2.055 -0.115 2.335 0.115 ;
        RECT  1.930 -0.115 2.055 0.140 ;
        RECT  0.885 -0.115 1.930 0.115 ;
        RECT  0.805 -0.115 0.885 0.280 ;
        RECT  0.340 -0.115 0.805 0.115 ;
        RECT  0.220 -0.115 0.340 0.190 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.720 3.170 1.375 ;
        RECT  2.790 1.145 3.090 1.375 ;
        RECT  2.715 0.985 2.790 1.375 ;
        RECT  2.410 1.145 2.715 1.375 ;
        RECT  2.330 0.785 2.410 1.375 ;
        RECT  2.025 1.145 2.330 1.375 ;
        RECT  1.955 1.005 2.025 1.375 ;
        RECT  0.900 1.145 1.955 1.375 ;
        RECT  0.790 1.000 0.900 1.375 ;
        RECT  0.340 1.145 0.790 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.185 2.980 0.480 ;
        RECT  2.905 0.755 2.980 1.035 ;
        RECT  2.525 0.185 2.555 0.480 ;
        RECT  2.525 0.755 2.555 1.040 ;
        RECT  2.425 0.550 2.555 0.640 ;
        RECT  2.355 0.350 2.425 0.640 ;
        RECT  1.485 0.350 2.355 0.420 ;
        RECT  1.565 0.210 2.240 0.280 ;
        RECT  1.560 0.845 2.240 0.915 ;
        RECT  1.365 0.995 1.870 1.065 ;
        RECT  1.560 0.570 1.660 0.765 ;
        RECT  1.340 0.570 1.560 0.640 ;
        RECT  1.415 0.195 1.485 0.420 ;
        RECT  1.170 0.195 1.415 0.265 ;
        RECT  1.290 0.720 1.365 1.065 ;
        RECT  1.240 0.345 1.340 0.640 ;
        RECT  1.170 0.720 1.290 0.790 ;
        RECT  1.040 0.995 1.220 1.065 ;
        RECT  1.100 0.195 1.170 0.790 ;
        RECT  0.830 0.720 1.100 0.790 ;
        RECT  0.970 0.860 1.040 1.065 ;
        RECT  0.935 0.360 1.005 0.640 ;
        RECT  0.525 0.860 0.970 0.930 ;
        RECT  0.680 0.360 0.935 0.430 ;
        RECT  0.760 0.510 0.830 0.790 ;
        RECT  0.680 0.195 0.710 0.265 ;
        RECT  0.610 0.195 0.680 0.790 ;
        RECT  0.590 0.195 0.610 0.265 ;
        RECT  0.450 0.295 0.525 1.005 ;
        RECT  0.420 0.295 0.450 0.395 ;
        RECT  0.430 0.860 0.450 1.005 ;
        RECT  0.340 0.550 0.380 0.670 ;
        RECT  0.270 0.260 0.340 0.920 ;
        RECT  0.055 0.260 0.270 0.380 ;
        RECT  0.130 0.850 0.270 0.920 ;
        RECT  0.050 0.850 0.130 1.060 ;
    END
END LHQD4BWP40

MACRO LHSNQD0BWP40
    CLASS CORE ;
    FOREIGN LHSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.810 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.060 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.740 2.415 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.355 0.805 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 -0.115 2.520 0.115 ;
        RECT  2.200 -0.115 2.280 0.290 ;
        RECT  1.530 -0.115 2.200 0.115 ;
        RECT  1.460 -0.115 1.530 0.260 ;
        RECT  0.745 -0.115 1.460 0.115 ;
        RECT  0.645 -0.115 0.745 0.270 ;
        RECT  0.335 -0.115 0.645 0.115 ;
        RECT  0.220 -0.115 0.335 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.200 0.975 2.280 1.375 ;
        RECT  1.910 1.145 2.200 1.375 ;
        RECT  1.830 0.980 1.910 1.375 ;
        RECT  1.540 1.145 1.830 1.375 ;
        RECT  1.440 0.990 1.540 1.375 ;
        RECT  0.730 1.145 1.440 1.375 ;
        RECT  0.660 1.000 0.730 1.375 ;
        RECT  0.310 1.145 0.660 1.375 ;
        RECT  0.220 0.990 0.310 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.525 2.345 0.635 ;
        RECT  2.050 0.205 2.120 1.050 ;
        RECT  1.980 0.205 2.050 0.275 ;
        RECT  2.000 0.980 2.050 1.050 ;
        RECT  1.895 0.345 1.970 0.910 ;
        RECT  1.885 0.185 1.895 0.910 ;
        RECT  1.825 0.185 1.885 0.415 ;
        RECT  1.720 0.840 1.885 0.910 ;
        RECT  1.480 0.340 1.825 0.415 ;
        RECT  1.640 0.840 1.720 1.060 ;
        RECT  1.450 0.645 1.615 0.715 ;
        RECT  1.360 0.340 1.480 0.440 ;
        RECT  1.380 0.540 1.450 0.920 ;
        RECT  1.245 0.540 1.380 0.610 ;
        RECT  1.050 0.850 1.380 0.920 ;
        RECT  1.095 0.690 1.260 0.780 ;
        RECT  1.175 0.185 1.245 0.610 ;
        RECT  1.060 0.185 1.175 0.265 ;
        RECT  1.015 0.335 1.095 0.780 ;
        RECT  0.970 1.005 1.040 1.075 ;
        RECT  1.010 0.335 1.015 0.465 ;
        RECT  0.530 0.695 1.015 0.780 ;
        RECT  0.900 0.850 0.970 1.075 ;
        RECT  0.380 0.850 0.900 0.920 ;
        RECT  0.460 0.185 0.530 0.780 ;
        RECT  0.310 0.315 0.380 0.920 ;
        RECT  0.145 0.315 0.310 0.390 ;
        RECT  0.125 0.850 0.310 0.920 ;
        RECT  0.055 0.200 0.145 0.390 ;
        RECT  0.055 0.850 0.125 1.000 ;
    END
END LHSNQD0BWP40

MACRO LHSNQD1BWP40
    CLASS CORE ;
    FOREIGN LHSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.495 1.805 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.060 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.740 2.415 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.255 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.495 0.945 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 -0.115 2.520 0.115 ;
        RECT  2.200 -0.115 2.280 0.455 ;
        RECT  1.530 -0.115 2.200 0.115 ;
        RECT  1.460 -0.115 1.530 0.260 ;
        RECT  0.780 -0.115 1.460 0.115 ;
        RECT  0.680 -0.115 0.780 0.425 ;
        RECT  0.370 -0.115 0.680 0.115 ;
        RECT  0.250 -0.115 0.370 0.225 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.200 0.800 2.280 1.375 ;
        RECT  1.910 1.145 2.200 1.375 ;
        RECT  1.830 0.980 1.910 1.375 ;
        RECT  1.545 1.145 1.830 1.375 ;
        RECT  1.435 0.985 1.545 1.375 ;
        RECT  0.810 1.145 1.435 1.375 ;
        RECT  0.680 1.130 0.810 1.375 ;
        RECT  0.310 1.145 0.680 1.375 ;
        RECT  0.220 0.990 0.310 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 0.525 2.345 0.635 ;
        RECT  2.050 0.205 2.120 1.050 ;
        RECT  1.970 0.205 2.050 0.275 ;
        RECT  2.000 0.980 2.050 1.050 ;
        RECT  1.885 0.345 1.970 0.910 ;
        RECT  1.325 0.345 1.885 0.415 ;
        RECT  1.720 0.840 1.885 0.910 ;
        RECT  1.640 0.840 1.720 1.030 ;
        RECT  1.410 0.535 1.620 0.615 ;
        RECT  1.340 0.535 1.410 0.915 ;
        RECT  1.240 0.535 1.340 0.605 ;
        RECT  1.040 0.845 1.340 0.915 ;
        RECT  1.090 0.675 1.265 0.775 ;
        RECT  1.170 0.195 1.240 0.605 ;
        RECT  1.160 0.195 1.170 0.265 ;
        RECT  1.040 0.185 1.160 0.265 ;
        RECT  1.020 0.335 1.090 0.775 ;
        RECT  0.915 0.990 1.085 1.075 ;
        RECT  0.960 0.335 1.020 0.415 ;
        RECT  0.620 0.695 1.020 0.775 ;
        RECT  0.450 0.990 0.915 1.060 ;
        RECT  0.610 0.695 0.620 0.900 ;
        RECT  0.520 0.185 0.610 0.900 ;
        RECT  0.380 0.315 0.450 1.060 ;
        RECT  0.145 0.315 0.380 0.390 ;
        RECT  0.145 0.850 0.380 0.920 ;
        RECT  0.035 0.200 0.145 0.390 ;
        RECT  0.035 0.850 0.145 1.025 ;
    END
END LHSNQD1BWP40

MACRO LHSNQD2BWP40
    CLASS CORE ;
    FOREIGN LHSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.495 1.785 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 0.355 2.485 0.770 ;
        RECT  2.415 0.185 2.440 1.060 ;
        RECT  2.345 0.185 2.415 0.460 ;
        RECT  2.345 0.700 2.415 1.060 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.355 0.805 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.615 -0.115 2.660 0.115 ;
        RECT  2.525 -0.115 2.615 0.275 ;
        RECT  2.240 -0.115 2.525 0.115 ;
        RECT  2.160 -0.115 2.240 0.450 ;
        RECT  1.480 -0.115 2.160 0.115 ;
        RECT  1.410 -0.115 1.480 0.265 ;
        RECT  0.725 -0.115 1.410 0.115 ;
        RECT  0.625 -0.115 0.725 0.270 ;
        RECT  0.340 -0.115 0.625 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.535 0.820 2.610 1.375 ;
        RECT  2.240 1.145 2.535 1.375 ;
        RECT  2.160 0.800 2.240 1.375 ;
        RECT  1.860 1.145 2.160 1.375 ;
        RECT  1.780 0.985 1.860 1.375 ;
        RECT  1.495 1.145 1.780 1.375 ;
        RECT  1.380 0.995 1.495 1.375 ;
        RECT  0.720 1.145 1.380 1.375 ;
        RECT  0.625 1.000 0.720 1.375 ;
        RECT  0.310 1.145 0.625 1.375 ;
        RECT  0.220 0.990 0.310 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.080 0.545 2.345 0.615 ;
        RECT  2.010 0.205 2.080 1.065 ;
        RECT  1.935 0.205 2.010 0.275 ;
        RECT  1.950 0.995 2.010 1.065 ;
        RECT  1.855 0.345 1.925 0.915 ;
        RECT  1.845 0.345 1.855 0.415 ;
        RECT  1.670 0.845 1.855 0.915 ;
        RECT  1.775 0.185 1.845 0.415 ;
        RECT  1.275 0.345 1.775 0.415 ;
        RECT  1.590 0.845 1.670 1.055 ;
        RECT  1.365 0.530 1.570 0.615 ;
        RECT  1.295 0.530 1.365 0.915 ;
        RECT  1.195 0.530 1.295 0.600 ;
        RECT  1.010 0.845 1.295 0.915 ;
        RECT  1.015 0.680 1.225 0.765 ;
        RECT  1.125 0.185 1.195 0.600 ;
        RECT  1.010 0.185 1.125 0.265 ;
        RECT  1.015 0.350 1.055 0.420 ;
        RECT  0.920 0.990 1.030 1.075 ;
        RECT  0.930 0.350 1.015 0.765 ;
        RECT  0.565 0.695 0.930 0.765 ;
        RECT  0.850 0.850 0.920 1.075 ;
        RECT  0.385 0.850 0.850 0.920 ;
        RECT  0.535 0.695 0.565 0.780 ;
        RECT  0.465 0.185 0.535 0.780 ;
        RECT  0.315 0.315 0.385 0.920 ;
        RECT  0.125 0.315 0.315 0.390 ;
        RECT  0.130 0.850 0.315 0.920 ;
        RECT  0.055 0.850 0.130 0.995 ;
        RECT  0.055 0.200 0.125 0.390 ;
    END
END LHSNQD2BWP40

MACRO LHSNQD4BWP40
    CLASS CORE ;
    FOREIGN LHSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.495 1.925 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.190 2.980 0.465 ;
        RECT  2.900 0.715 2.980 0.995 ;
        RECT  2.835 0.345 2.900 0.465 ;
        RECT  2.835 0.715 2.900 0.860 ;
        RECT  2.625 0.345 2.835 0.860 ;
        RECT  2.605 0.345 2.625 0.465 ;
        RECT  2.600 0.715 2.625 0.860 ;
        RECT  2.520 0.185 2.605 0.465 ;
        RECT  2.520 0.715 2.600 0.995 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.630 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.345 0.805 0.625 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.445 ;
        RECT  2.785 -0.115 3.095 0.115 ;
        RECT  2.710 -0.115 2.785 0.275 ;
        RECT  2.415 -0.115 2.710 0.115 ;
        RECT  2.325 -0.115 2.415 0.470 ;
        RECT  2.025 -0.115 2.325 0.115 ;
        RECT  1.955 -0.115 2.025 0.275 ;
        RECT  1.470 -0.115 1.955 0.115 ;
        RECT  1.400 -0.115 1.470 0.265 ;
        RECT  0.720 -0.115 1.400 0.115 ;
        RECT  0.620 -0.115 0.720 0.270 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 1.145 3.220 1.375 ;
        RECT  3.090 0.720 3.165 1.375 ;
        RECT  2.785 1.145 3.090 1.375 ;
        RECT  2.710 1.005 2.785 1.375 ;
        RECT  2.410 1.145 2.710 1.375 ;
        RECT  2.330 0.725 2.410 1.375 ;
        RECT  2.025 1.145 2.330 1.375 ;
        RECT  1.955 0.935 2.025 1.375 ;
        RECT  1.845 1.145 1.955 1.375 ;
        RECT  1.775 0.935 1.845 1.375 ;
        RECT  1.485 1.145 1.775 1.375 ;
        RECT  1.375 0.995 1.485 1.375 ;
        RECT  0.715 1.145 1.375 1.375 ;
        RECT  0.630 1.030 0.715 1.375 ;
        RECT  0.345 1.145 0.630 1.375 ;
        RECT  0.220 1.020 0.345 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.190 2.980 0.465 ;
        RECT  2.905 0.715 2.980 0.995 ;
        RECT  2.520 0.185 2.555 0.465 ;
        RECT  2.520 0.715 2.555 0.995 ;
        RECT  2.215 0.545 2.550 0.615 ;
        RECT  2.145 0.185 2.215 1.050 ;
        RECT  1.995 0.345 2.065 0.850 ;
        RECT  1.265 0.345 1.995 0.415 ;
        RECT  1.660 0.780 1.995 0.850 ;
        RECT  1.580 0.780 1.660 1.060 ;
        RECT  1.360 0.530 1.560 0.615 ;
        RECT  1.290 0.530 1.360 0.915 ;
        RECT  1.185 0.530 1.290 0.600 ;
        RECT  1.000 0.845 1.290 0.915 ;
        RECT  1.005 0.680 1.220 0.765 ;
        RECT  1.115 0.185 1.185 0.600 ;
        RECT  1.000 0.185 1.115 0.265 ;
        RECT  1.005 0.350 1.045 0.430 ;
        RECT  0.910 0.990 1.025 1.075 ;
        RECT  0.935 0.350 1.005 0.765 ;
        RECT  0.550 0.695 0.935 0.765 ;
        RECT  0.840 0.875 0.910 1.075 ;
        RECT  0.385 0.875 0.840 0.950 ;
        RECT  0.530 0.695 0.550 0.780 ;
        RECT  0.460 0.185 0.530 0.780 ;
        RECT  0.315 0.315 0.385 0.950 ;
        RECT  0.125 0.315 0.315 0.390 ;
        RECT  0.130 0.880 0.315 0.950 ;
        RECT  0.055 0.880 0.130 0.990 ;
        RECT  0.055 0.200 0.125 0.390 ;
    END
END LHSNQD4BWP40

MACRO LNCNQD0BWP40
    CLASS CORE ;
    FOREIGN LNCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.765 1.045 ;
        RECT  2.670 0.185 2.695 0.465 ;
        RECT  2.670 0.705 2.695 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.350 0.460 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.640 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.020800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.350 1.830 0.485 ;
        RECT  0.805 0.350 1.575 0.420 ;
        RECT  0.715 0.350 0.805 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 -0.115 2.800 0.115 ;
        RECT  2.460 -0.115 2.580 0.250 ;
        RECT  1.975 -0.115 2.460 0.115 ;
        RECT  1.855 -0.115 1.975 0.140 ;
        RECT  0.820 -0.115 1.855 0.115 ;
        RECT  0.700 -0.115 0.820 0.255 ;
        RECT  0.365 -0.115 0.700 0.115 ;
        RECT  0.285 -0.115 0.365 0.240 ;
        RECT  0.000 -0.115 0.285 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.555 1.145 2.800 1.375 ;
        RECT  2.485 0.955 2.555 1.375 ;
        RECT  1.975 1.145 2.485 1.375 ;
        RECT  1.855 1.140 1.975 1.375 ;
        RECT  1.045 1.145 1.855 1.375 ;
        RECT  0.925 1.130 1.045 1.375 ;
        RECT  0.385 1.145 0.925 1.375 ;
        RECT  0.265 1.135 0.385 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.575 0.520 2.625 0.640 ;
        RECT  2.505 0.345 2.575 0.825 ;
        RECT  2.365 0.345 2.505 0.425 ;
        RECT  2.370 0.745 2.505 0.825 ;
        RECT  2.290 0.745 2.370 1.040 ;
        RECT  2.295 0.185 2.365 0.425 ;
        RECT  2.180 0.520 2.335 0.640 ;
        RECT  2.100 0.185 2.180 1.060 ;
        RECT  1.825 0.990 2.100 1.060 ;
        RECT  1.935 0.210 2.005 0.920 ;
        RECT  1.255 0.210 1.935 0.280 ;
        RECT  0.705 0.850 1.935 0.920 ;
        RECT  1.675 0.990 1.825 1.075 ;
        RECT  1.325 0.710 1.695 0.780 ;
        RECT  1.235 0.990 1.445 1.075 ;
        RECT  1.205 0.490 1.325 0.780 ;
        RECT  0.105 0.990 1.235 1.060 ;
        RECT  0.610 0.710 1.205 0.780 ;
        RECT  0.540 0.195 0.610 0.780 ;
        RECT  0.245 0.710 0.540 0.780 ;
        RECT  0.175 0.520 0.245 0.780 ;
        RECT  0.105 0.195 0.160 0.270 ;
        RECT  0.035 0.195 0.105 1.060 ;
    END
END LNCNQD0BWP40

MACRO LNCNQD1BWP40
    CLASS CORE ;
    FOREIGN LNCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.087400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.185 2.765 1.045 ;
        RECT  2.670 0.185 2.695 0.465 ;
        RECT  2.670 0.705 2.695 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.350 0.460 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.640 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.350 1.830 0.625 ;
        RECT  0.805 0.350 1.715 0.420 ;
        RECT  0.715 0.350 0.805 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.580 -0.115 2.800 0.115 ;
        RECT  2.460 -0.115 2.580 0.250 ;
        RECT  1.975 -0.115 2.460 0.115 ;
        RECT  1.855 -0.115 1.975 0.140 ;
        RECT  0.820 -0.115 1.855 0.115 ;
        RECT  0.700 -0.115 0.820 0.255 ;
        RECT  0.365 -0.115 0.700 0.115 ;
        RECT  0.285 -0.115 0.365 0.270 ;
        RECT  0.000 -0.115 0.285 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.555 1.145 2.800 1.375 ;
        RECT  2.485 0.910 2.555 1.375 ;
        RECT  1.975 1.145 2.485 1.375 ;
        RECT  1.855 1.140 1.975 1.375 ;
        RECT  1.045 1.145 1.855 1.375 ;
        RECT  0.925 1.130 1.045 1.375 ;
        RECT  0.385 1.145 0.925 1.375 ;
        RECT  0.265 1.135 0.385 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.575 0.520 2.625 0.640 ;
        RECT  2.505 0.345 2.575 0.825 ;
        RECT  2.370 0.345 2.505 0.445 ;
        RECT  2.370 0.745 2.505 0.825 ;
        RECT  2.180 0.540 2.380 0.615 ;
        RECT  2.295 0.195 2.370 0.445 ;
        RECT  2.290 0.745 2.370 1.010 ;
        RECT  2.100 0.185 2.180 1.060 ;
        RECT  1.825 0.990 2.100 1.060 ;
        RECT  1.935 0.210 2.005 0.920 ;
        RECT  1.255 0.210 1.935 0.280 ;
        RECT  0.705 0.850 1.935 0.920 ;
        RECT  1.675 0.990 1.825 1.075 ;
        RECT  1.325 0.710 1.695 0.780 ;
        RECT  1.235 0.990 1.445 1.075 ;
        RECT  1.205 0.490 1.325 0.780 ;
        RECT  0.105 0.990 1.235 1.060 ;
        RECT  0.610 0.710 1.205 0.780 ;
        RECT  0.540 0.195 0.610 0.910 ;
        RECT  0.245 0.745 0.540 0.815 ;
        RECT  0.175 0.520 0.245 0.815 ;
        RECT  0.105 0.195 0.160 0.270 ;
        RECT  0.035 0.195 0.105 1.060 ;
    END
END LNCNQD1BWP40

MACRO LNCNQD2BWP40
    CLASS CORE ;
    FOREIGN LNCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.114000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 0.355 2.765 0.775 ;
        RECT  2.695 0.185 2.720 1.045 ;
        RECT  2.620 0.185 2.695 0.465 ;
        RECT  2.620 0.705 2.695 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.350 0.460 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.640 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.350 1.805 0.625 ;
        RECT  0.805 0.350 1.715 0.420 ;
        RECT  0.715 0.350 0.805 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.885 0.255 ;
        RECT  2.530 -0.115 2.810 0.115 ;
        RECT  2.410 -0.115 2.530 0.250 ;
        RECT  1.950 -0.115 2.410 0.115 ;
        RECT  1.830 -0.115 1.950 0.140 ;
        RECT  0.820 -0.115 1.830 0.115 ;
        RECT  0.700 -0.115 0.820 0.270 ;
        RECT  0.365 -0.115 0.700 0.115 ;
        RECT  0.285 -0.115 0.365 0.270 ;
        RECT  0.000 -0.115 0.285 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.815 0.825 2.890 1.375 ;
        RECT  2.505 1.145 2.815 1.375 ;
        RECT  2.435 0.955 2.505 1.375 ;
        RECT  1.950 1.145 2.435 1.375 ;
        RECT  1.830 1.140 1.950 1.375 ;
        RECT  1.045 1.145 1.830 1.375 ;
        RECT  0.925 1.130 1.045 1.375 ;
        RECT  0.385 1.145 0.925 1.375 ;
        RECT  0.265 1.135 0.385 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.525 0.520 2.575 0.640 ;
        RECT  2.455 0.365 2.525 0.825 ;
        RECT  2.315 0.365 2.455 0.445 ;
        RECT  2.315 0.745 2.455 0.825 ;
        RECT  2.145 0.540 2.345 0.615 ;
        RECT  2.245 0.185 2.315 0.445 ;
        RECT  2.245 0.745 2.315 1.055 ;
        RECT  2.065 0.185 2.145 1.060 ;
        RECT  1.800 0.990 2.065 1.060 ;
        RECT  1.910 0.210 1.980 0.920 ;
        RECT  1.230 0.210 1.910 0.280 ;
        RECT  0.705 0.850 1.910 0.920 ;
        RECT  1.650 0.990 1.800 1.075 ;
        RECT  1.300 0.710 1.670 0.780 ;
        RECT  1.210 0.990 1.420 1.075 ;
        RECT  1.180 0.490 1.300 0.780 ;
        RECT  0.105 0.990 1.210 1.060 ;
        RECT  0.610 0.710 1.180 0.780 ;
        RECT  0.540 0.195 0.610 0.920 ;
        RECT  0.245 0.850 0.540 0.920 ;
        RECT  0.175 0.520 0.245 0.920 ;
        RECT  0.105 0.195 0.160 0.270 ;
        RECT  0.035 0.195 0.105 1.060 ;
    END
END LNCNQD2BWP40

MACRO LNCNQD4BWP40
    CLASS CORE ;
    FOREIGN LNCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.228000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 0.185 3.260 0.460 ;
        RECT  3.180 0.755 3.260 1.050 ;
        RECT  3.115 0.350 3.180 0.460 ;
        RECT  3.115 0.755 3.180 0.905 ;
        RECT  2.905 0.350 3.115 0.905 ;
        RECT  2.890 0.350 2.905 0.460 ;
        RECT  2.885 0.755 2.905 0.905 ;
        RECT  2.805 0.185 2.890 0.460 ;
        RECT  2.805 0.755 2.885 1.050 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.350 0.460 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.640 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.025800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.350 1.795 0.625 ;
        RECT  0.805 0.350 1.715 0.420 ;
        RECT  0.715 0.350 0.805 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.115 3.500 0.115 ;
        RECT  3.365 -0.115 3.445 0.435 ;
        RECT  3.070 -0.115 3.365 0.115 ;
        RECT  2.990 -0.115 3.070 0.275 ;
        RECT  2.690 -0.115 2.990 0.115 ;
        RECT  2.610 -0.115 2.690 0.435 ;
        RECT  2.310 -0.115 2.610 0.115 ;
        RECT  2.235 -0.115 2.310 0.435 ;
        RECT  1.940 -0.115 2.235 0.115 ;
        RECT  1.820 -0.115 1.940 0.140 ;
        RECT  0.820 -0.115 1.820 0.115 ;
        RECT  0.700 -0.115 0.820 0.255 ;
        RECT  0.365 -0.115 0.700 0.115 ;
        RECT  0.285 -0.115 0.365 0.240 ;
        RECT  0.000 -0.115 0.285 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.725 3.450 1.375 ;
        RECT  3.070 1.145 3.370 1.375 ;
        RECT  2.990 1.000 3.070 1.375 ;
        RECT  2.690 1.145 2.990 1.375 ;
        RECT  2.610 0.725 2.690 1.375 ;
        RECT  2.310 1.145 2.610 1.375 ;
        RECT  2.235 0.815 2.310 1.375 ;
        RECT  1.940 1.145 2.235 1.375 ;
        RECT  1.820 1.140 1.940 1.375 ;
        RECT  1.045 1.145 1.820 1.375 ;
        RECT  0.925 1.130 1.045 1.375 ;
        RECT  0.385 1.145 0.925 1.375 ;
        RECT  0.265 1.135 0.385 1.375 ;
        RECT  0.000 1.145 0.265 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.185 3.260 0.460 ;
        RECT  3.185 0.755 3.260 1.050 ;
        RECT  2.805 0.185 2.835 0.460 ;
        RECT  2.805 0.755 2.835 1.050 ;
        RECT  2.500 0.550 2.830 0.620 ;
        RECT  2.425 0.185 2.500 1.040 ;
        RECT  2.135 0.545 2.265 0.620 ;
        RECT  2.055 0.185 2.135 1.060 ;
        RECT  1.790 0.990 2.055 1.060 ;
        RECT  1.900 0.210 1.970 0.920 ;
        RECT  1.230 0.210 1.900 0.280 ;
        RECT  0.705 0.850 1.900 0.920 ;
        RECT  1.640 0.990 1.790 1.075 ;
        RECT  1.315 0.710 1.660 0.780 ;
        RECT  1.200 0.990 1.410 1.075 ;
        RECT  1.170 0.490 1.315 0.780 ;
        RECT  0.105 0.990 1.200 1.060 ;
        RECT  0.610 0.710 1.170 0.780 ;
        RECT  0.540 0.195 0.610 0.780 ;
        RECT  0.245 0.710 0.540 0.780 ;
        RECT  0.175 0.520 0.245 0.780 ;
        RECT  0.105 0.195 0.160 0.270 ;
        RECT  0.035 0.195 0.105 1.060 ;
    END
END LNCNQD4BWP40

MACRO LNCSNQD0BWP40
    CLASS CORE ;
    FOREIGN LNCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.535 1.610 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.054000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.185 1.060 ;
        RECT  3.090 0.185 3.115 0.465 ;
        RECT  3.090 0.740 3.115 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.355 0.980 0.515 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.485 0.765 ;
        RECT  2.340 0.555 2.415 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 -0.115 3.220 0.115 ;
        RECT  2.860 -0.115 2.980 0.235 ;
        RECT  2.510 -0.115 2.860 0.115 ;
        RECT  2.440 -0.115 2.510 0.405 ;
        RECT  1.495 -0.115 2.440 0.115 ;
        RECT  1.425 -0.115 1.495 0.250 ;
        RECT  0.695 -0.115 1.425 0.115 ;
        RECT  0.605 -0.115 0.695 0.260 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.955 1.145 3.220 1.375 ;
        RECT  2.885 0.985 2.955 1.375 ;
        RECT  2.540 1.145 2.885 1.375 ;
        RECT  2.420 1.135 2.540 1.375 ;
        RECT  2.120 1.145 2.420 1.375 ;
        RECT  2.000 1.130 2.120 1.375 ;
        RECT  1.530 1.145 2.000 1.375 ;
        RECT  1.410 1.135 1.530 1.375 ;
        RECT  0.685 1.145 1.410 1.375 ;
        RECT  0.615 0.800 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.980 0.520 3.025 0.645 ;
        RECT  2.910 0.305 2.980 0.795 ;
        RECT  2.735 0.305 2.910 0.375 ;
        RECT  2.765 0.720 2.910 0.795 ;
        RECT  2.625 0.520 2.835 0.640 ;
        RECT  2.695 0.720 2.765 1.030 ;
        RECT  2.665 0.200 2.735 0.375 ;
        RECT  2.555 0.520 2.625 1.055 ;
        RECT  1.935 0.980 2.555 1.055 ;
        RECT  2.095 0.840 2.330 0.910 ;
        RECT  2.095 0.360 2.325 0.430 ;
        RECT  1.630 0.205 2.140 0.275 ;
        RECT  2.025 0.360 2.095 0.910 ;
        RECT  1.865 0.345 1.935 1.055 ;
        RECT  1.825 0.345 1.865 0.445 ;
        RECT  1.380 0.985 1.865 1.055 ;
        RECT  1.750 0.535 1.795 0.655 ;
        RECT  1.680 0.345 1.750 0.915 ;
        RECT  1.330 0.345 1.680 0.415 ;
        RECT  0.980 0.845 1.680 0.915 ;
        RECT  1.255 0.985 1.380 1.070 ;
        RECT  1.250 0.205 1.330 0.415 ;
        RECT  0.980 0.205 1.250 0.275 ;
        RECT  1.075 0.410 1.165 0.665 ;
        RECT  0.530 0.595 1.075 0.665 ;
        RECT  0.460 0.190 0.530 1.035 ;
        RECT  0.435 0.190 0.460 0.335 ;
        RECT  0.440 0.915 0.460 1.035 ;
        RECT  0.345 0.520 0.380 0.640 ;
        RECT  0.275 0.325 0.345 0.960 ;
        RECT  0.150 0.325 0.275 0.405 ;
        RECT  0.145 0.890 0.275 0.960 ;
        RECT  0.035 0.215 0.150 0.405 ;
        RECT  0.035 0.890 0.145 1.040 ;
    END
END LNCSNQD0BWP40

MACRO LNCSNQD1BWP40
    CLASS CORE ;
    FOREIGN LNCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.535 1.610 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.108000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.185 3.185 1.060 ;
        RECT  3.090 0.185 3.115 0.465 ;
        RECT  3.090 0.740 3.115 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.355 0.980 0.515 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.265 0.555 2.485 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 -0.115 3.220 0.115 ;
        RECT  2.860 -0.115 2.980 0.235 ;
        RECT  2.510 -0.115 2.860 0.115 ;
        RECT  2.440 -0.115 2.510 0.405 ;
        RECT  1.495 -0.115 2.440 0.115 ;
        RECT  1.425 -0.115 1.495 0.250 ;
        RECT  0.695 -0.115 1.425 0.115 ;
        RECT  0.605 -0.115 0.695 0.260 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.955 1.145 3.220 1.375 ;
        RECT  2.885 0.875 2.955 1.375 ;
        RECT  2.540 1.145 2.885 1.375 ;
        RECT  2.420 1.135 2.540 1.375 ;
        RECT  2.120 1.145 2.420 1.375 ;
        RECT  2.000 1.130 2.120 1.375 ;
        RECT  1.530 1.145 2.000 1.375 ;
        RECT  1.410 1.135 1.530 1.375 ;
        RECT  0.685 1.145 1.410 1.375 ;
        RECT  0.615 0.800 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.980 0.520 3.025 0.645 ;
        RECT  2.910 0.330 2.980 0.795 ;
        RECT  2.745 0.330 2.910 0.440 ;
        RECT  2.765 0.720 2.910 0.795 ;
        RECT  2.625 0.520 2.835 0.640 ;
        RECT  2.695 0.720 2.765 1.030 ;
        RECT  2.660 0.190 2.745 0.440 ;
        RECT  2.555 0.520 2.625 1.055 ;
        RECT  1.935 0.980 2.555 1.055 ;
        RECT  2.120 0.840 2.330 0.910 ;
        RECT  2.120 0.395 2.325 0.465 ;
        RECT  1.630 0.205 2.140 0.275 ;
        RECT  2.050 0.395 2.120 0.910 ;
        RECT  1.865 0.345 1.935 1.055 ;
        RECT  1.830 0.345 1.865 0.445 ;
        RECT  1.380 0.985 1.865 1.055 ;
        RECT  1.750 0.535 1.795 0.655 ;
        RECT  1.680 0.345 1.750 0.915 ;
        RECT  1.330 0.345 1.680 0.415 ;
        RECT  0.980 0.845 1.680 0.915 ;
        RECT  1.255 0.985 1.380 1.070 ;
        RECT  1.250 0.205 1.330 0.415 ;
        RECT  0.980 0.205 1.250 0.275 ;
        RECT  1.075 0.410 1.165 0.665 ;
        RECT  0.530 0.595 1.075 0.665 ;
        RECT  0.460 0.190 0.530 1.035 ;
        RECT  0.435 0.190 0.460 0.335 ;
        RECT  0.440 0.915 0.460 1.035 ;
        RECT  0.345 0.520 0.380 0.640 ;
        RECT  0.275 0.325 0.345 0.960 ;
        RECT  0.150 0.325 0.275 0.405 ;
        RECT  0.145 0.890 0.275 0.960 ;
        RECT  0.035 0.215 0.150 0.405 ;
        RECT  0.035 0.890 0.145 1.040 ;
    END
END LNCSNQD1BWP40

MACRO LNCSNQD2BWP40
    CLASS CORE ;
    FOREIGN LNCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.545 1.580 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 0.355 3.185 0.795 ;
        RECT  3.120 0.355 3.130 1.060 ;
        RECT  3.115 0.185 3.120 1.060 ;
        RECT  3.040 0.185 3.115 0.455 ;
        RECT  3.040 0.715 3.115 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.355 0.965 0.515 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.555 2.415 0.765 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 -0.115 3.360 0.115 ;
        RECT  3.230 -0.115 3.305 0.255 ;
        RECT  2.950 -0.115 3.230 0.115 ;
        RECT  2.830 -0.115 2.950 0.235 ;
        RECT  2.480 -0.115 2.830 0.115 ;
        RECT  2.410 -0.115 2.480 0.435 ;
        RECT  1.475 -0.115 2.410 0.115 ;
        RECT  1.405 -0.115 1.475 0.310 ;
        RECT  0.695 -0.115 1.405 0.115 ;
        RECT  0.605 -0.115 0.695 0.275 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.305 1.145 3.360 1.375 ;
        RECT  3.230 0.865 3.305 1.375 ;
        RECT  2.925 1.145 3.230 1.375 ;
        RECT  2.855 0.865 2.925 1.375 ;
        RECT  2.510 1.145 2.855 1.375 ;
        RECT  2.390 1.135 2.510 1.375 ;
        RECT  2.090 1.145 2.390 1.375 ;
        RECT  1.970 1.130 2.090 1.375 ;
        RECT  1.510 1.145 1.970 1.375 ;
        RECT  1.390 1.135 1.510 1.375 ;
        RECT  0.685 1.145 1.390 1.375 ;
        RECT  0.615 0.800 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.950 0.525 3.045 0.635 ;
        RECT  2.880 0.305 2.950 0.795 ;
        RECT  2.600 0.305 2.880 0.375 ;
        RECT  2.735 0.720 2.880 0.795 ;
        RECT  2.595 0.520 2.805 0.640 ;
        RECT  2.665 0.720 2.735 1.030 ;
        RECT  2.525 0.520 2.595 1.055 ;
        RECT  1.900 0.985 2.525 1.055 ;
        RECT  2.040 0.835 2.300 0.905 ;
        RECT  2.040 0.395 2.295 0.465 ;
        RECT  1.600 0.205 2.110 0.275 ;
        RECT  1.970 0.395 2.040 0.905 ;
        RECT  1.830 0.345 1.900 1.055 ;
        RECT  1.800 0.345 1.830 0.445 ;
        RECT  1.360 0.985 1.830 1.055 ;
        RECT  1.720 0.530 1.760 0.655 ;
        RECT  1.650 0.395 1.720 0.915 ;
        RECT  1.310 0.395 1.650 0.465 ;
        RECT  0.960 0.845 1.650 0.915 ;
        RECT  1.235 0.985 1.360 1.070 ;
        RECT  1.230 0.205 1.310 0.465 ;
        RECT  0.960 0.205 1.230 0.275 ;
        RECT  1.055 0.410 1.145 0.665 ;
        RECT  0.530 0.595 1.055 0.665 ;
        RECT  0.460 0.190 0.530 1.035 ;
        RECT  0.435 0.190 0.460 0.335 ;
        RECT  0.440 0.915 0.460 1.035 ;
        RECT  0.345 0.520 0.380 0.640 ;
        RECT  0.275 0.325 0.345 0.960 ;
        RECT  0.150 0.325 0.275 0.405 ;
        RECT  0.145 0.890 0.275 0.960 ;
        RECT  0.035 0.215 0.150 0.405 ;
        RECT  0.035 0.890 0.145 1.040 ;
    END
END LNCSNQD2BWP40

MACRO LNCSNQD4BWP40
    CLASS CORE ;
    FOREIGN LNCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.545 1.580 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.460 0.185 3.540 0.460 ;
        RECT  3.460 0.755 3.540 1.050 ;
        RECT  3.395 0.350 3.460 0.460 ;
        RECT  3.395 0.755 3.460 0.905 ;
        RECT  3.185 0.350 3.395 0.905 ;
        RECT  3.170 0.350 3.185 0.460 ;
        RECT  3.165 0.755 3.185 0.905 ;
        RECT  3.085 0.185 3.170 0.460 ;
        RECT  3.085 0.755 3.165 1.050 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.355 0.965 0.515 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 0.770 2.625 0.910 ;
        RECT  2.365 0.635 2.490 0.910 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.115 3.780 0.115 ;
        RECT  3.645 -0.115 3.725 0.465 ;
        RECT  3.350 -0.115 3.645 0.115 ;
        RECT  3.270 -0.115 3.350 0.275 ;
        RECT  2.970 -0.115 3.270 0.115 ;
        RECT  2.890 -0.115 2.970 0.320 ;
        RECT  2.580 -0.115 2.890 0.115 ;
        RECT  2.455 -0.115 2.580 0.125 ;
        RECT  1.475 -0.115 2.455 0.115 ;
        RECT  1.405 -0.115 1.475 0.250 ;
        RECT  0.695 -0.115 1.405 0.115 ;
        RECT  0.605 -0.115 0.695 0.275 ;
        RECT  0.340 -0.115 0.605 0.115 ;
        RECT  0.220 -0.115 0.340 0.225 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.720 3.730 1.375 ;
        RECT  3.350 1.145 3.650 1.375 ;
        RECT  3.270 1.000 3.350 1.375 ;
        RECT  2.975 1.145 3.270 1.375 ;
        RECT  2.885 0.885 2.975 1.375 ;
        RECT  2.590 1.145 2.885 1.375 ;
        RECT  2.490 1.005 2.590 1.375 ;
        RECT  2.160 1.145 2.490 1.375 ;
        RECT  2.040 1.130 2.160 1.375 ;
        RECT  1.510 1.145 2.040 1.375 ;
        RECT  1.390 1.135 1.510 1.375 ;
        RECT  0.685 1.145 1.390 1.375 ;
        RECT  0.615 0.800 0.685 1.375 ;
        RECT  0.340 1.145 0.615 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.465 0.185 3.540 0.460 ;
        RECT  3.465 0.755 3.540 1.050 ;
        RECT  3.085 0.185 3.115 0.460 ;
        RECT  3.085 0.755 3.115 1.050 ;
        RECT  2.955 0.550 3.110 0.620 ;
        RECT  2.885 0.400 2.955 0.815 ;
        RECT  2.785 0.400 2.885 0.470 ;
        RECT  2.780 0.745 2.885 0.815 ;
        RECT  2.710 0.185 2.785 0.470 ;
        RECT  2.630 0.540 2.785 0.610 ;
        RECT  2.705 0.745 2.780 1.040 ;
        RECT  2.560 0.215 2.630 0.610 ;
        RECT  2.250 0.215 2.560 0.285 ;
        RECT  2.320 0.370 2.410 0.565 ;
        RECT  2.085 0.980 2.410 1.050 ;
        RECT  2.085 0.495 2.320 0.565 ;
        RECT  2.180 0.215 2.250 0.415 ;
        RECT  1.900 0.345 2.180 0.415 ;
        RECT  1.600 0.195 2.110 0.265 ;
        RECT  2.015 0.495 2.085 1.050 ;
        RECT  1.830 0.345 1.900 1.055 ;
        RECT  1.360 0.985 1.830 1.055 ;
        RECT  1.720 0.530 1.760 0.655 ;
        RECT  1.650 0.345 1.720 0.915 ;
        RECT  1.310 0.345 1.650 0.415 ;
        RECT  0.960 0.845 1.650 0.915 ;
        RECT  1.235 0.985 1.360 1.070 ;
        RECT  1.230 0.205 1.310 0.415 ;
        RECT  0.960 0.205 1.230 0.275 ;
        RECT  1.055 0.410 1.145 0.665 ;
        RECT  0.530 0.595 1.055 0.665 ;
        RECT  0.460 0.190 0.530 1.035 ;
        RECT  0.435 0.190 0.460 0.335 ;
        RECT  0.440 0.915 0.460 1.035 ;
        RECT  0.345 0.520 0.380 0.640 ;
        RECT  0.275 0.325 0.345 0.960 ;
        RECT  0.150 0.325 0.275 0.405 ;
        RECT  0.145 0.890 0.275 0.960 ;
        RECT  0.035 0.215 0.150 0.405 ;
        RECT  0.035 0.890 0.145 1.040 ;
    END
END LNCSNQD4BWP40

MACRO LNQD0BWP40
    CLASS CORE ;
    FOREIGN LNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 1.045 ;
        RECT  1.835 0.185 1.855 0.305 ;
        RECT  1.835 0.745 1.855 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.500 0.495 1.575 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.115 1.960 0.115 ;
        RECT  1.610 -0.115 1.735 0.235 ;
        RECT  0.930 -0.115 1.610 0.115 ;
        RECT  0.810 -0.115 0.930 0.290 ;
        RECT  0.340 -0.115 0.810 0.115 ;
        RECT  0.220 -0.115 0.340 0.240 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.145 1.960 1.375 ;
        RECT  1.635 0.895 1.715 1.375 ;
        RECT  0.930 1.145 1.635 1.375 ;
        RECT  0.810 1.025 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.540 0.355 1.715 0.425 ;
        RECT  1.470 0.200 1.540 0.425 ;
        RECT  1.435 0.685 1.505 1.065 ;
        RECT  1.240 0.200 1.470 0.270 ;
        RECT  1.400 0.685 1.435 0.755 ;
        RECT  1.090 0.995 1.435 1.065 ;
        RECT  1.330 0.370 1.400 0.755 ;
        RECT  1.240 0.840 1.355 0.910 ;
        RECT  1.160 0.200 1.240 0.910 ;
        RECT  0.855 0.720 1.160 0.790 ;
        RECT  1.020 0.885 1.090 1.065 ;
        RECT  0.970 0.365 1.060 0.640 ;
        RECT  0.340 0.885 1.020 0.955 ;
        RECT  0.710 0.365 0.970 0.435 ;
        RECT  0.780 0.520 0.855 0.790 ;
        RECT  0.640 0.210 0.710 0.815 ;
        RECT  0.620 0.210 0.640 0.350 ;
        RECT  0.600 0.715 0.640 0.815 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.205 0.525 0.815 ;
        RECT  0.420 0.205 0.455 0.305 ;
        RECT  0.425 0.695 0.455 0.815 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.320 0.340 0.955 ;
        RECT  0.145 0.320 0.270 0.390 ;
        RECT  0.145 0.885 0.270 0.955 ;
        RECT  0.035 0.195 0.145 0.390 ;
        RECT  0.035 0.885 0.145 1.040 ;
    END
END LNQD0BWP40

MACRO LNQD1BWP40
    CLASS CORE ;
    FOREIGN LNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.185 1.925 1.045 ;
        RECT  1.835 0.185 1.855 0.305 ;
        RECT  1.835 0.745 1.855 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.765 ;
        RECT  1.500 0.495 1.575 0.615 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.115 1.960 0.115 ;
        RECT  1.610 -0.115 1.735 0.275 ;
        RECT  0.930 -0.115 1.610 0.115 ;
        RECT  0.810 -0.115 0.930 0.290 ;
        RECT  0.340 -0.115 0.810 0.115 ;
        RECT  0.220 -0.115 0.340 0.240 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.145 1.960 1.375 ;
        RECT  1.635 0.850 1.715 1.375 ;
        RECT  0.930 1.145 1.635 1.375 ;
        RECT  0.810 1.025 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.355 1.785 0.640 ;
        RECT  1.540 0.355 1.715 0.425 ;
        RECT  1.470 0.200 1.540 0.425 ;
        RECT  1.435 0.685 1.505 1.065 ;
        RECT  1.240 0.200 1.470 0.270 ;
        RECT  1.400 0.685 1.435 0.755 ;
        RECT  1.090 0.995 1.435 1.065 ;
        RECT  1.330 0.370 1.400 0.755 ;
        RECT  1.240 0.840 1.355 0.910 ;
        RECT  1.160 0.200 1.240 0.910 ;
        RECT  0.855 0.720 1.160 0.790 ;
        RECT  1.020 0.885 1.090 1.065 ;
        RECT  0.970 0.365 1.060 0.640 ;
        RECT  0.340 0.885 1.020 0.955 ;
        RECT  0.710 0.365 0.970 0.435 ;
        RECT  0.780 0.520 0.855 0.790 ;
        RECT  0.640 0.210 0.710 0.815 ;
        RECT  0.620 0.210 0.640 0.350 ;
        RECT  0.600 0.715 0.640 0.815 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.195 0.525 0.815 ;
        RECT  0.420 0.195 0.455 0.295 ;
        RECT  0.425 0.695 0.455 0.815 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.320 0.340 0.955 ;
        RECT  0.145 0.320 0.270 0.390 ;
        RECT  0.145 0.885 0.270 0.955 ;
        RECT  0.035 0.195 0.145 0.390 ;
        RECT  0.035 0.885 0.145 1.015 ;
    END
END LNQD1BWP40

MACRO LNQD2BWP40
    CLASS CORE ;
    FOREIGN LNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.117750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.355 1.925 0.765 ;
        RECT  1.860 0.355 1.875 1.045 ;
        RECT  1.855 0.185 1.860 1.045 ;
        RECT  1.790 0.185 1.855 0.425 ;
        RECT  1.785 0.685 1.855 1.045 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.031400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.665 1.675 0.905 ;
        RECT  1.495 0.515 1.580 0.905 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.975 -0.115 2.050 0.255 ;
        RECT  1.665 -0.115 1.975 0.115 ;
        RECT  1.595 -0.115 1.665 0.255 ;
        RECT  0.895 -0.115 1.595 0.115 ;
        RECT  0.785 -0.115 0.895 0.290 ;
        RECT  0.340 -0.115 0.785 0.115 ;
        RECT  0.220 -0.115 0.340 0.240 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.145 2.100 1.375 ;
        RECT  1.970 0.850 2.050 1.375 ;
        RECT  1.670 1.145 1.970 1.375 ;
        RECT  1.590 0.985 1.670 1.375 ;
        RECT  0.900 1.145 1.590 1.375 ;
        RECT  0.780 1.025 0.900 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.720 0.505 1.785 0.595 ;
        RECT  1.650 0.355 1.720 0.595 ;
        RECT  1.525 0.355 1.650 0.425 ;
        RECT  1.455 0.200 1.525 0.425 ;
        RECT  1.190 0.200 1.455 0.270 ;
        RECT  1.370 0.660 1.425 1.065 ;
        RECT  1.355 0.370 1.370 1.065 ;
        RECT  1.300 0.370 1.355 0.730 ;
        RECT  1.040 0.995 1.355 1.065 ;
        RECT  1.190 0.805 1.285 0.920 ;
        RECT  1.110 0.200 1.190 0.920 ;
        RECT  0.850 0.720 1.110 0.790 ;
        RECT  0.970 0.885 1.040 1.065 ;
        RECT  0.950 0.365 1.030 0.640 ;
        RECT  0.340 0.885 0.970 0.955 ;
        RECT  0.710 0.365 0.950 0.435 ;
        RECT  0.780 0.520 0.850 0.790 ;
        RECT  0.640 0.210 0.710 0.815 ;
        RECT  0.620 0.210 0.640 0.350 ;
        RECT  0.600 0.715 0.640 0.815 ;
        RECT  0.525 0.520 0.570 0.640 ;
        RECT  0.455 0.195 0.525 0.815 ;
        RECT  0.420 0.195 0.455 0.295 ;
        RECT  0.425 0.695 0.455 0.815 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.320 0.340 0.955 ;
        RECT  0.145 0.320 0.270 0.390 ;
        RECT  0.145 0.885 0.270 0.955 ;
        RECT  0.035 0.195 0.145 0.390 ;
        RECT  0.035 0.885 0.145 1.035 ;
    END
END LNQD2BWP40

MACRO LNQD4BWP40
    CLASS CORE ;
    FOREIGN LNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.185 2.980 0.480 ;
        RECT  2.900 0.755 2.980 1.035 ;
        RECT  2.835 0.350 2.900 0.480 ;
        RECT  2.835 0.755 2.900 0.910 ;
        RECT  2.625 0.350 2.835 0.910 ;
        RECT  2.600 0.350 2.625 0.480 ;
        RECT  2.600 0.755 2.625 0.910 ;
        RECT  2.525 0.185 2.600 0.480 ;
        RECT  2.525 0.755 2.600 1.040 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.205 0.625 ;
        RECT  1.995 0.495 2.065 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.170 0.465 ;
        RECT  2.795 -0.115 3.095 0.115 ;
        RECT  2.715 -0.115 2.795 0.275 ;
        RECT  2.405 -0.115 2.715 0.115 ;
        RECT  2.335 -0.115 2.405 0.255 ;
        RECT  2.055 -0.115 2.335 0.115 ;
        RECT  1.930 -0.115 2.055 0.140 ;
        RECT  0.895 -0.115 1.930 0.115 ;
        RECT  0.785 -0.115 0.895 0.260 ;
        RECT  0.340 -0.115 0.785 0.115 ;
        RECT  0.220 -0.115 0.340 0.240 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.720 3.170 1.375 ;
        RECT  2.790 1.145 3.090 1.375 ;
        RECT  2.715 0.985 2.790 1.375 ;
        RECT  2.410 1.145 2.715 1.375 ;
        RECT  2.330 0.755 2.410 1.375 ;
        RECT  2.025 1.145 2.330 1.375 ;
        RECT  1.955 1.005 2.025 1.375 ;
        RECT  0.900 1.145 1.955 1.375 ;
        RECT  0.780 1.030 0.900 1.375 ;
        RECT  0.340 1.145 0.780 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.185 2.980 0.480 ;
        RECT  2.905 0.755 2.980 1.035 ;
        RECT  2.525 0.185 2.555 0.480 ;
        RECT  2.525 0.755 2.555 1.040 ;
        RECT  2.425 0.550 2.555 0.640 ;
        RECT  2.355 0.350 2.425 0.640 ;
        RECT  1.485 0.350 2.355 0.420 ;
        RECT  1.565 0.210 2.240 0.280 ;
        RECT  2.135 0.845 2.235 1.075 ;
        RECT  1.560 0.845 2.135 0.915 ;
        RECT  1.465 0.995 1.870 1.065 ;
        RECT  1.570 0.535 1.675 0.765 ;
        RECT  1.340 0.535 1.570 0.605 ;
        RECT  1.415 0.195 1.485 0.420 ;
        RECT  1.390 0.720 1.465 1.065 ;
        RECT  1.170 0.195 1.415 0.265 ;
        RECT  1.285 0.720 1.390 0.790 ;
        RECT  1.240 0.345 1.340 0.605 ;
        RECT  1.215 0.720 1.285 0.835 ;
        RECT  1.040 0.995 1.220 1.065 ;
        RECT  1.170 0.720 1.215 0.790 ;
        RECT  1.100 0.195 1.170 0.790 ;
        RECT  0.850 0.720 1.100 0.790 ;
        RECT  0.970 0.890 1.040 1.065 ;
        RECT  0.950 0.365 1.020 0.610 ;
        RECT  0.340 0.890 0.970 0.960 ;
        RECT  0.710 0.365 0.950 0.435 ;
        RECT  0.780 0.520 0.850 0.790 ;
        RECT  0.640 0.195 0.710 0.815 ;
        RECT  0.590 0.195 0.640 0.265 ;
        RECT  0.600 0.715 0.640 0.815 ;
        RECT  0.520 0.520 0.570 0.640 ;
        RECT  0.450 0.205 0.520 0.815 ;
        RECT  0.420 0.205 0.450 0.305 ;
        RECT  0.425 0.695 0.450 0.815 ;
        RECT  0.340 0.520 0.380 0.640 ;
        RECT  0.270 0.320 0.340 0.960 ;
        RECT  0.145 0.320 0.270 0.390 ;
        RECT  0.145 0.885 0.270 0.960 ;
        RECT  0.035 0.195 0.145 0.390 ;
        RECT  0.035 0.885 0.145 1.035 ;
    END
END LNQD4BWP40

MACRO LNSNQD0BWP40
    CLASS CORE ;
    FOREIGN LNSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.495 1.925 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.070725 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.060 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.740 2.415 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.290 0.145 ;
        RECT  1.510 -0.115 2.170 0.115 ;
        RECT  1.430 -0.115 1.510 0.290 ;
        RECT  0.695 -0.115 1.430 0.115 ;
        RECT  0.615 -0.115 0.695 0.260 ;
        RECT  0.330 -0.115 0.615 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.160 1.005 2.280 1.375 ;
        RECT  1.885 1.145 2.160 1.375 ;
        RECT  1.815 0.855 1.885 1.375 ;
        RECT  1.560 1.145 1.815 1.375 ;
        RECT  1.440 1.135 1.560 1.375 ;
        RECT  0.740 1.145 1.440 1.375 ;
        RECT  0.620 1.130 0.740 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.240 1.135 0.355 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.300 0.520 2.345 0.640 ;
        RECT  2.230 0.215 2.300 0.930 ;
        RECT  1.970 0.215 2.230 0.285 ;
        RECT  1.980 0.860 2.230 0.930 ;
        RECT  2.005 0.355 2.075 0.785 ;
        RECT  1.885 0.355 2.005 0.425 ;
        RECT  1.695 0.715 2.005 0.785 ;
        RECT  1.815 0.190 1.885 0.425 ;
        RECT  1.625 0.715 1.695 1.065 ;
        RECT  1.300 0.990 1.625 1.065 ;
        RECT  1.540 0.520 1.575 0.640 ;
        RECT  1.470 0.390 1.540 0.900 ;
        RECT  1.270 0.390 1.470 0.460 ;
        RECT  1.000 0.830 1.470 0.900 ;
        RECT  1.200 0.185 1.270 0.460 ;
        RECT  1.120 0.690 1.260 0.760 ;
        RECT  1.015 0.185 1.200 0.255 ;
        RECT  1.050 0.355 1.120 0.760 ;
        RECT  0.515 0.355 1.050 0.425 ;
        RECT  0.875 0.970 1.015 1.075 ;
        RECT  0.105 0.970 0.875 1.040 ;
        RECT  0.300 0.805 0.520 0.875 ;
        RECT  0.405 0.205 0.515 0.425 ;
        RECT  0.300 0.355 0.405 0.425 ;
        RECT  0.230 0.355 0.300 0.875 ;
        RECT  0.105 0.195 0.150 0.275 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END LNSNQD0BWP40

MACRO LNSNQD1BWP40
    CLASS CORE ;
    FOREIGN LNSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.026000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.495 1.925 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.087400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.185 2.485 1.060 ;
        RECT  2.395 0.185 2.415 0.465 ;
        RECT  2.395 0.740 2.415 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.640 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.290 -0.115 2.520 0.115 ;
        RECT  2.170 -0.115 2.290 0.145 ;
        RECT  1.510 -0.115 2.170 0.115 ;
        RECT  1.430 -0.115 1.510 0.290 ;
        RECT  0.695 -0.115 1.430 0.115 ;
        RECT  0.615 -0.115 0.695 0.260 ;
        RECT  0.330 -0.115 0.615 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.145 2.520 1.375 ;
        RECT  2.160 1.005 2.280 1.375 ;
        RECT  1.885 1.145 2.160 1.375 ;
        RECT  1.815 0.865 1.885 1.375 ;
        RECT  1.560 1.145 1.815 1.375 ;
        RECT  1.440 1.135 1.560 1.375 ;
        RECT  0.740 1.145 1.440 1.375 ;
        RECT  0.620 1.130 0.740 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.240 1.135 0.355 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.300 0.520 2.345 0.640 ;
        RECT  2.230 0.215 2.300 0.930 ;
        RECT  1.970 0.215 2.230 0.285 ;
        RECT  1.980 0.860 2.230 0.930 ;
        RECT  2.005 0.355 2.075 0.785 ;
        RECT  1.790 0.355 2.005 0.425 ;
        RECT  1.695 0.715 2.005 0.785 ;
        RECT  1.625 0.715 1.695 1.055 ;
        RECT  1.300 0.980 1.625 1.055 ;
        RECT  1.540 0.520 1.575 0.640 ;
        RECT  1.470 0.390 1.540 0.900 ;
        RECT  1.270 0.390 1.470 0.460 ;
        RECT  1.000 0.830 1.470 0.900 ;
        RECT  1.200 0.185 1.270 0.460 ;
        RECT  1.120 0.675 1.240 0.745 ;
        RECT  1.015 0.185 1.200 0.255 ;
        RECT  1.050 0.345 1.120 0.745 ;
        RECT  0.515 0.345 1.050 0.415 ;
        RECT  0.875 0.970 1.015 1.075 ;
        RECT  0.105 0.970 0.875 1.040 ;
        RECT  0.300 0.805 0.520 0.875 ;
        RECT  0.405 0.205 0.515 0.415 ;
        RECT  0.300 0.345 0.405 0.415 ;
        RECT  0.230 0.345 0.300 0.875 ;
        RECT  0.105 0.195 0.150 0.275 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END LNSNQD1BWP40

MACRO LNSNQD2BWP40
    CLASS CORE ;
    FOREIGN LNSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.026000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.495 1.925 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.114000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.355 2.485 0.780 ;
        RECT  2.415 0.185 2.435 1.060 ;
        RECT  2.345 0.185 2.415 0.455 ;
        RECT  2.345 0.710 2.415 1.060 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.635 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.605 -0.115 2.660 0.115 ;
        RECT  2.535 -0.115 2.605 0.295 ;
        RECT  2.250 -0.115 2.535 0.115 ;
        RECT  2.130 -0.115 2.250 0.145 ;
        RECT  1.480 -0.115 2.130 0.115 ;
        RECT  1.400 -0.115 1.480 0.290 ;
        RECT  0.695 -0.115 1.400 0.115 ;
        RECT  0.615 -0.115 0.695 0.260 ;
        RECT  0.330 -0.115 0.615 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.615 1.145 2.660 1.375 ;
        RECT  2.530 0.835 2.615 1.375 ;
        RECT  2.250 1.145 2.530 1.375 ;
        RECT  2.130 1.005 2.250 1.375 ;
        RECT  1.855 1.145 2.130 1.375 ;
        RECT  1.785 0.865 1.855 1.375 ;
        RECT  1.530 1.145 1.785 1.375 ;
        RECT  1.410 1.135 1.530 1.375 ;
        RECT  0.740 1.145 1.410 1.375 ;
        RECT  0.620 1.130 0.740 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.240 1.135 0.355 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.250 0.525 2.345 0.635 ;
        RECT  2.180 0.215 2.250 0.930 ;
        RECT  1.940 0.215 2.180 0.285 ;
        RECT  1.950 0.860 2.180 0.930 ;
        RECT  1.995 0.355 2.065 0.785 ;
        RECT  1.710 0.355 1.995 0.425 ;
        RECT  1.665 0.715 1.995 0.785 ;
        RECT  1.595 0.715 1.665 1.055 ;
        RECT  1.270 0.980 1.595 1.055 ;
        RECT  1.510 0.520 1.545 0.640 ;
        RECT  1.440 0.390 1.510 0.900 ;
        RECT  1.260 0.390 1.440 0.460 ;
        RECT  0.990 0.830 1.440 0.900 ;
        RECT  1.190 0.185 1.260 0.460 ;
        RECT  1.110 0.675 1.230 0.745 ;
        RECT  0.995 0.185 1.190 0.255 ;
        RECT  1.040 0.345 1.110 0.745 ;
        RECT  0.515 0.345 1.040 0.415 ;
        RECT  0.865 0.970 1.005 1.075 ;
        RECT  0.105 0.970 0.865 1.040 ;
        RECT  0.300 0.805 0.520 0.875 ;
        RECT  0.405 0.205 0.515 0.415 ;
        RECT  0.300 0.345 0.405 0.415 ;
        RECT  0.230 0.345 0.300 0.875 ;
        RECT  0.105 0.195 0.150 0.275 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END LNSNQD2BWP40

MACRO LNSNQD4BWP40
    CLASS CORE ;
    FOREIGN LNSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SDN
        ANTENNAGATEAREA 0.026000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.495 1.925 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.228000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.190 2.980 0.465 ;
        RECT  2.900 0.715 2.980 0.995 ;
        RECT  2.835 0.345 2.900 0.465 ;
        RECT  2.835 0.715 2.900 0.860 ;
        RECT  2.625 0.345 2.835 0.860 ;
        RECT  2.605 0.345 2.625 0.465 ;
        RECT  2.600 0.715 2.625 0.860 ;
        RECT  2.520 0.185 2.605 0.465 ;
        RECT  2.520 0.715 2.600 0.995 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.640 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.635 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 -0.115 3.220 0.115 ;
        RECT  3.095 -0.115 3.165 0.445 ;
        RECT  2.785 -0.115 3.095 0.115 ;
        RECT  2.710 -0.115 2.785 0.275 ;
        RECT  2.415 -0.115 2.710 0.115 ;
        RECT  2.325 -0.115 2.415 0.470 ;
        RECT  2.025 -0.115 2.325 0.115 ;
        RECT  1.955 -0.115 2.025 0.280 ;
        RECT  1.470 -0.115 1.955 0.115 ;
        RECT  1.390 -0.115 1.470 0.290 ;
        RECT  0.695 -0.115 1.390 0.115 ;
        RECT  0.615 -0.115 0.695 0.260 ;
        RECT  0.330 -0.115 0.615 0.115 ;
        RECT  0.230 -0.115 0.330 0.250 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.165 1.145 3.220 1.375 ;
        RECT  3.090 0.720 3.165 1.375 ;
        RECT  2.785 1.145 3.090 1.375 ;
        RECT  2.710 1.005 2.785 1.375 ;
        RECT  2.410 1.145 2.710 1.375 ;
        RECT  2.330 0.805 2.410 1.375 ;
        RECT  2.025 1.145 2.330 1.375 ;
        RECT  1.955 0.845 2.025 1.375 ;
        RECT  1.845 1.145 1.955 1.375 ;
        RECT  1.775 0.845 1.845 1.375 ;
        RECT  1.520 1.145 1.775 1.375 ;
        RECT  1.400 1.135 1.520 1.375 ;
        RECT  0.740 1.145 1.400 1.375 ;
        RECT  0.620 1.130 0.740 1.375 ;
        RECT  0.355 1.145 0.620 1.375 ;
        RECT  0.240 1.135 0.355 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.905 0.190 2.980 0.465 ;
        RECT  2.905 0.715 2.980 0.995 ;
        RECT  2.520 0.185 2.555 0.465 ;
        RECT  2.520 0.715 2.555 0.995 ;
        RECT  2.215 0.545 2.550 0.615 ;
        RECT  2.145 0.185 2.215 1.050 ;
        RECT  1.995 0.355 2.065 0.775 ;
        RECT  1.740 0.355 1.995 0.425 ;
        RECT  1.655 0.705 1.995 0.775 ;
        RECT  1.585 0.705 1.655 1.055 ;
        RECT  1.260 0.980 1.585 1.055 ;
        RECT  1.500 0.520 1.535 0.640 ;
        RECT  1.430 0.390 1.500 0.900 ;
        RECT  1.250 0.390 1.430 0.460 ;
        RECT  0.980 0.830 1.430 0.900 ;
        RECT  1.180 0.185 1.250 0.460 ;
        RECT  1.100 0.675 1.220 0.745 ;
        RECT  0.985 0.185 1.180 0.255 ;
        RECT  1.030 0.345 1.100 0.745 ;
        RECT  0.515 0.345 1.030 0.415 ;
        RECT  0.855 0.970 0.995 1.075 ;
        RECT  0.105 0.970 0.855 1.040 ;
        RECT  0.300 0.805 0.520 0.875 ;
        RECT  0.405 0.205 0.515 0.415 ;
        RECT  0.300 0.345 0.405 0.415 ;
        RECT  0.230 0.345 0.300 0.875 ;
        RECT  0.105 0.195 0.150 0.275 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END LNSNQD4BWP40

MACRO MAOI222D0BWP40
    CLASS CORE ;
    FOREIGN MAOI222D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.124000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.795 ;
        RECT  0.920 0.355 1.155 0.425 ;
        RECT  1.015 0.725 1.155 0.795 ;
        RECT  0.945 0.725 1.015 0.925 ;
        RECT  0.130 0.855 0.945 0.925 ;
        RECT  0.105 0.855 0.130 1.055 ;
        RECT  0.105 0.215 0.125 0.375 ;
        RECT  0.035 0.215 0.105 1.055 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.635 0.805 0.785 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.645 ;
        RECT  0.445 0.495 0.875 0.565 ;
        RECT  0.410 0.495 0.445 0.765 ;
        RECT  0.315 0.355 0.410 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 -0.115 1.260 0.115 ;
        RECT  0.500 -0.115 0.575 0.415 ;
        RECT  0.000 -0.115 0.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.145 1.260 1.375 ;
        RECT  0.510 0.995 0.590 1.375 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.120 0.185 1.220 0.285 ;
        RECT  1.130 0.895 1.210 1.065 ;
        RECT  0.680 0.995 1.130 1.065 ;
        RECT  0.800 0.205 1.120 0.275 ;
        RECT  0.720 0.205 0.800 0.425 ;
    END
END MAOI222D0BWP40

MACRO MAOI222D1BWP40
    CLASS CORE ;
    FOREIGN MAOI222D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.204925 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.225 0.795 ;
        RECT  0.920 0.355 1.155 0.425 ;
        RECT  1.015 0.725 1.155 0.795 ;
        RECT  0.945 0.725 1.015 0.925 ;
        RECT  0.130 0.855 0.945 0.925 ;
        RECT  0.105 0.855 0.130 1.055 ;
        RECT  0.105 0.215 0.125 0.375 ;
        RECT  0.035 0.215 0.105 1.055 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.022200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.635 0.805 0.785 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.047800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.955 0.645 ;
        RECT  0.445 0.495 0.875 0.565 ;
        RECT  0.410 0.495 0.445 0.765 ;
        RECT  0.315 0.355 0.410 0.765 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.445 0.245 0.765 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 -0.115 1.260 0.115 ;
        RECT  0.500 -0.115 0.570 0.400 ;
        RECT  0.000 -0.115 0.500 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.145 1.260 1.375 ;
        RECT  0.510 0.995 0.590 1.375 ;
        RECT  0.000 1.145 0.510 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.120 0.185 1.220 0.285 ;
        RECT  1.130 0.895 1.210 1.065 ;
        RECT  0.680 0.995 1.130 1.065 ;
        RECT  0.800 0.205 1.120 0.275 ;
        RECT  0.720 0.205 0.800 0.425 ;
    END
END MAOI222D1BWP40

MACRO MAOI222D2BWP40
    CLASS CORE ;
    FOREIGN MAOI222D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.403675 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.635 2.485 1.065 ;
        RECT  2.225 0.855 2.380 0.925 ;
        RECT  2.135 0.355 2.225 0.925 ;
        RECT  1.710 0.355 2.135 0.425 ;
        RECT  0.115 0.855 2.135 0.925 ;
        RECT  0.115 0.335 0.590 0.425 ;
        RECT  0.035 0.335 0.115 0.925 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.042800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.635 1.550 0.785 ;
        RECT  1.015 0.635 1.295 0.725 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.095600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.495 1.925 0.625 ;
        RECT  0.845 0.495 1.690 0.565 ;
        RECT  0.775 0.495 0.845 0.785 ;
        RECT  0.265 0.710 0.775 0.785 ;
        RECT  0.185 0.515 0.265 0.785 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.355 0.495 0.685 0.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 -0.115 2.520 0.115 ;
        RECT  1.315 -0.115 1.435 0.275 ;
        RECT  1.000 -0.115 1.315 0.115 ;
        RECT  0.880 -0.115 1.000 0.380 ;
        RECT  0.150 -0.115 0.880 0.115 ;
        RECT  0.035 -0.115 0.150 0.265 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.420 1.145 2.520 1.375 ;
        RECT  1.295 1.135 1.420 1.375 ;
        RECT  0.995 1.145 1.295 1.375 ;
        RECT  0.915 0.995 0.995 1.375 ;
        RECT  0.150 1.145 0.915 1.375 ;
        RECT  0.045 0.995 0.150 1.375 ;
        RECT  0.000 1.145 0.045 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.205 2.425 0.485 ;
        RECT  1.620 0.205 2.345 0.275 ;
        RECT  1.085 0.995 2.220 1.065 ;
        RECT  1.540 0.205 1.620 0.425 ;
        RECT  1.085 0.355 1.540 0.425 ;
        RECT  0.245 0.995 0.770 1.065 ;
        RECT  0.240 0.195 0.755 0.265 ;
    END
END MAOI222D2BWP40

MACRO MAOI222D4BWP40
    CLASS CORE ;
    FOREIGN MAOI222D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.695700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.330 0.725 4.420 1.025 ;
        RECT  4.235 0.725 4.330 0.795 ;
        RECT  4.030 0.355 4.235 0.795 ;
        RECT  4.025 0.355 4.030 0.925 ;
        RECT  2.985 0.355 4.025 0.425 ;
        RECT  3.960 0.725 4.025 0.925 ;
        RECT  0.115 0.855 3.960 0.925 ;
        RECT  0.115 0.335 1.470 0.425 ;
        RECT  0.035 0.335 0.115 0.925 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.085600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.635 2.785 0.785 ;
        RECT  1.860 0.635 2.415 0.725 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.191200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.930 0.495 3.300 0.625 ;
        RECT  1.715 0.495 2.930 0.565 ;
        RECT  1.575 0.495 1.715 0.640 ;
        RECT  0.945 0.495 1.575 0.565 ;
        RECT  0.875 0.495 0.945 0.785 ;
        RECT  0.265 0.710 0.875 0.785 ;
        RECT  0.185 0.515 0.265 0.785 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.355 0.495 0.685 0.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.670 -0.115 4.480 0.115 ;
        RECT  2.545 -0.115 2.670 0.275 ;
        RECT  2.290 -0.115 2.545 0.115 ;
        RECT  2.165 -0.115 2.290 0.275 ;
        RECT  1.845 -0.115 2.165 0.115 ;
        RECT  1.765 -0.115 1.845 0.400 ;
        RECT  1.000 -0.115 1.765 0.115 ;
        RECT  0.880 -0.115 1.000 0.265 ;
        RECT  0.150 -0.115 0.880 0.115 ;
        RECT  0.050 -0.115 0.150 0.265 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.145 4.480 1.375 ;
        RECT  2.570 1.135 2.695 1.375 ;
        RECT  2.270 1.145 2.570 1.375 ;
        RECT  2.145 1.135 2.270 1.375 ;
        RECT  1.840 1.145 2.145 1.375 ;
        RECT  1.760 0.995 1.840 1.375 ;
        RECT  0.995 1.145 1.760 1.375 ;
        RECT  0.915 0.995 0.995 1.375 ;
        RECT  0.150 1.145 0.915 1.375 ;
        RECT  0.045 0.995 0.150 1.375 ;
        RECT  0.000 1.145 0.045 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.330 0.725 4.420 1.025 ;
        RECT  4.305 0.725 4.330 0.795 ;
        RECT  2.985 0.355 3.955 0.425 ;
        RECT  0.115 0.855 3.955 0.925 ;
        RECT  0.115 0.335 1.470 0.425 ;
        RECT  0.035 0.335 0.115 0.925 ;
        RECT  2.895 0.205 4.435 0.275 ;
        RECT  1.935 0.995 4.245 1.065 ;
        RECT  2.815 0.205 2.895 0.425 ;
        RECT  1.935 0.355 2.815 0.425 ;
    END
END MAOI222D4BWP40

MACRO MAOI22D0BWP40
    CLASS CORE ;
    FOREIGN MAOI22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.079350 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 0.905 ;
        RECT  0.595 0.195 0.875 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.155 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.150 -0.115 1.260 0.115 ;
        RECT  1.070 -0.115 1.150 0.305 ;
        RECT  0.540 -0.115 1.070 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.145 1.260 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.985 1.180 1.055 ;
        RECT  0.525 0.520 0.610 0.650 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.220 0.215 0.455 0.285 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.020 ;
    END
END MAOI22D0BWP40

MACRO MAOI22D1BWP40
    CLASS CORE ;
    FOREIGN MAOI22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.138100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 0.905 ;
        RECT  0.595 0.195 0.875 0.275 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.150 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 0.805 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.150 -0.115 1.260 0.115 ;
        RECT  1.070 -0.115 1.150 0.420 ;
        RECT  0.540 -0.115 1.070 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.320 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.145 1.260 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.985 1.175 1.055 ;
        RECT  0.525 0.520 0.610 0.650 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.220 0.215 0.455 0.285 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.020 ;
    END
END MAOI22D1BWP40

MACRO MAOI22D2BWP40
    CLASS CORE ;
    FOREIGN MAOI22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.297800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.730 1.925 1.045 ;
        RECT  0.945 0.730 1.840 0.800 ;
        RECT  0.945 0.335 1.340 0.415 ;
        RECT  0.875 0.335 0.945 0.800 ;
        RECT  0.595 0.335 0.875 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.495 1.925 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.495 1.420 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.115 1.960 0.115 ;
        RECT  1.595 -0.115 1.725 0.215 ;
        RECT  0.940 -0.115 1.595 0.115 ;
        RECT  0.820 -0.115 0.940 0.135 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 1.960 1.375 ;
        RECT  0.830 1.010 0.930 1.375 ;
        RECT  0.530 1.145 0.830 1.375 ;
        RECT  0.430 0.995 0.530 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.495 0.335 1.910 0.415 ;
        RECT  0.620 0.870 1.720 0.940 ;
        RECT  1.425 0.195 1.495 0.415 ;
        RECT  1.000 0.195 1.425 0.265 ;
        RECT  0.525 0.520 0.670 0.650 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.220 0.215 0.455 0.285 ;
        RECT  0.130 0.845 0.455 0.915 ;
        RECT  0.050 0.845 0.130 1.020 ;
    END
END MAOI22D2BWP40

MACRO MAOI22D4BWP40
    CLASS CORE ;
    FOREIGN MAOI22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.514500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.730 3.605 1.045 ;
        RECT  1.995 0.730 3.515 0.800 ;
        RECT  1.995 0.335 2.660 0.415 ;
        RECT  1.785 0.335 1.995 0.800 ;
        RECT  1.285 0.335 1.785 0.415 ;
        RECT  1.200 0.230 1.285 0.415 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.495 0.980 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.325 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.495 3.325 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.085 0.495 2.495 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.425 -0.115 3.640 0.115 ;
        RECT  3.295 -0.115 3.425 0.215 ;
        RECT  3.035 -0.115 3.295 0.115 ;
        RECT  2.905 -0.115 3.035 0.215 ;
        RECT  1.890 -0.115 2.905 0.115 ;
        RECT  1.770 -0.115 1.890 0.135 ;
        RECT  1.490 -0.115 1.770 0.115 ;
        RECT  1.370 -0.115 1.490 0.250 ;
        RECT  1.110 -0.115 1.370 0.115 ;
        RECT  0.980 -0.115 1.110 0.250 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.580 -0.115 0.720 0.255 ;
        RECT  0.320 -0.115 0.580 0.115 ;
        RECT  0.240 -0.115 0.320 0.255 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.145 3.640 1.375 ;
        RECT  1.780 1.010 1.880 1.375 ;
        RECT  1.505 1.145 1.780 1.375 ;
        RECT  1.365 1.015 1.505 1.375 ;
        RECT  1.110 1.145 1.365 1.375 ;
        RECT  0.970 1.015 1.110 1.375 ;
        RECT  0.720 1.145 0.970 1.375 ;
        RECT  0.580 1.015 0.720 1.375 ;
        RECT  0.000 1.145 0.580 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.515 0.730 3.605 1.045 ;
        RECT  2.065 0.730 3.515 0.800 ;
        RECT  2.065 0.335 2.660 0.415 ;
        RECT  1.285 0.335 1.715 0.415 ;
        RECT  1.200 0.230 1.285 0.415 ;
        RECT  3.510 0.235 3.590 0.415 ;
        RECT  2.815 0.335 3.510 0.415 ;
        RECT  1.170 0.870 3.420 0.940 ;
        RECT  2.745 0.195 2.815 0.415 ;
        RECT  1.935 0.195 2.745 0.265 ;
        RECT  1.130 0.520 1.650 0.650 ;
        RECT  1.060 0.340 1.130 0.770 ;
        RECT  0.035 0.340 1.060 0.410 ;
        RECT  0.345 0.700 1.060 0.770 ;
        RECT  0.035 0.865 0.935 0.935 ;
        RECT  0.220 0.700 0.345 0.785 ;
    END
END MAOI22D4BWP40

MACRO MOAI22D0BWP40
    CLASS CORE ;
    FOREIGN MOAI22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.085250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.960 ;
        RECT  0.745 0.880 0.875 0.960 ;
        RECT  0.665 0.880 0.745 1.020 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.155 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.540 -0.115 1.260 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.145 1.260 1.375 ;
        RECT  1.070 0.960 1.150 1.375 ;
        RECT  0.515 1.145 1.070 1.375 ;
        RECT  0.445 0.975 0.515 1.375 ;
        RECT  0.130 1.145 0.445 1.375 ;
        RECT  0.050 0.940 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.640 0.205 1.170 0.275 ;
        RECT  0.525 0.520 0.610 0.640 ;
        RECT  0.455 0.205 0.525 0.885 ;
        RECT  0.035 0.205 0.455 0.275 ;
        RECT  0.320 0.815 0.455 0.885 ;
        RECT  0.240 0.815 0.320 1.075 ;
    END
END MOAI22D0BWP40

MACRO MOAI22D1BWP40
    CLASS CORE ;
    FOREIGN MOAI22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.140500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 0.945 0.960 ;
        RECT  0.745 0.880 0.875 0.960 ;
        RECT  0.665 0.880 0.745 1.020 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.355 0.385 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.355 1.225 0.640 ;
        RECT  1.015 0.495 1.150 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.540 -0.115 1.260 0.115 ;
        RECT  0.420 -0.115 0.540 0.135 ;
        RECT  0.000 -0.115 0.420 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.145 1.260 1.375 ;
        RECT  1.070 0.805 1.160 1.375 ;
        RECT  0.515 1.145 1.070 1.375 ;
        RECT  0.445 0.975 0.515 1.375 ;
        RECT  0.130 1.145 0.445 1.375 ;
        RECT  0.050 0.940 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.205 1.180 0.275 ;
        RECT  0.525 0.520 0.610 0.640 ;
        RECT  0.455 0.205 0.525 0.885 ;
        RECT  0.130 0.205 0.455 0.275 ;
        RECT  0.320 0.815 0.455 0.885 ;
        RECT  0.240 0.815 0.320 1.075 ;
        RECT  0.050 0.205 0.130 0.330 ;
    END
END MOAI22D1BWP40

MACRO MOAI22D2BWP40
    CLASS CORE ;
    FOREIGN MOAI22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.287800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 0.215 1.895 0.425 ;
        RECT  0.945 0.355 1.810 0.425 ;
        RECT  0.945 0.845 1.340 0.915 ;
        RECT  0.875 0.355 0.945 0.915 ;
        RECT  0.595 0.845 0.875 0.915 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 0.495 0.385 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 1.925 0.765 ;
        RECT  1.655 0.495 1.855 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.495 1.375 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.115 1.960 0.115 ;
        RECT  0.815 -0.115 0.945 0.145 ;
        RECT  0.520 -0.115 0.815 0.115 ;
        RECT  0.440 -0.115 0.520 0.260 ;
        RECT  0.000 -0.115 0.440 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 1.145 1.960 1.375 ;
        RECT  1.595 1.045 1.725 1.375 ;
        RECT  0.935 1.145 1.595 1.375 ;
        RECT  0.820 1.005 0.935 1.375 ;
        RECT  0.540 1.145 0.820 1.375 ;
        RECT  0.420 1.125 0.540 1.375 ;
        RECT  0.130 1.145 0.420 1.375 ;
        RECT  0.050 0.975 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.495 0.845 1.910 0.925 ;
        RECT  0.620 0.215 1.720 0.285 ;
        RECT  1.425 0.845 1.495 1.065 ;
        RECT  1.005 0.995 1.425 1.065 ;
        RECT  0.525 0.510 0.670 0.640 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.035 0.345 0.455 0.415 ;
        RECT  0.220 0.975 0.455 1.045 ;
    END
END MOAI22D2BWP40

MACRO MOAI22D4BWP40
    CLASS CORE ;
    FOREIGN MOAI22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.511500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.270 3.605 0.420 ;
        RECT  1.995 0.350 3.515 0.420 ;
        RECT  1.995 0.765 2.660 0.845 ;
        RECT  1.785 0.350 1.995 0.845 ;
        RECT  1.285 0.765 1.785 0.845 ;
        RECT  1.200 0.765 1.285 1.030 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.725 0.495 0.875 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.310 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 0.495 3.325 0.765 ;
        RECT  3.095 0.495 3.255 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.085 0.495 2.495 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.895 -0.115 3.640 0.115 ;
        RECT  1.765 -0.115 1.895 0.140 ;
        RECT  1.515 -0.115 1.765 0.115 ;
        RECT  1.370 -0.115 1.515 0.140 ;
        RECT  1.100 -0.115 1.370 0.115 ;
        RECT  0.980 -0.115 1.100 0.230 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.580 -0.115 0.720 0.140 ;
        RECT  0.000 -0.115 0.580 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.425 1.145 3.640 1.375 ;
        RECT  3.295 1.045 3.425 1.375 ;
        RECT  3.035 1.145 3.295 1.375 ;
        RECT  2.905 1.045 3.035 1.375 ;
        RECT  1.885 1.145 2.905 1.375 ;
        RECT  1.770 1.005 1.885 1.375 ;
        RECT  1.490 1.145 1.770 1.375 ;
        RECT  1.370 1.010 1.490 1.375 ;
        RECT  1.110 1.145 1.370 1.375 ;
        RECT  0.980 1.010 1.110 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.580 1.005 0.720 1.375 ;
        RECT  0.320 1.145 0.580 1.375 ;
        RECT  0.240 1.005 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.515 0.270 3.605 0.420 ;
        RECT  2.065 0.350 3.515 0.420 ;
        RECT  2.065 0.765 2.660 0.845 ;
        RECT  1.285 0.765 1.715 0.845 ;
        RECT  1.200 0.765 1.285 1.030 ;
        RECT  3.510 0.845 3.590 1.040 ;
        RECT  2.815 0.845 3.510 0.925 ;
        RECT  1.180 0.210 3.420 0.280 ;
        RECT  2.745 0.845 2.815 1.040 ;
        RECT  1.955 0.970 2.745 1.040 ;
        RECT  1.130 0.510 1.650 0.640 ;
        RECT  1.060 0.350 1.130 0.920 ;
        RECT  0.210 0.350 1.060 0.420 ;
        RECT  0.140 0.850 1.060 0.920 ;
        RECT  0.035 0.210 0.900 0.280 ;
        RECT  0.050 0.850 0.140 1.010 ;
    END
END MOAI22D4BWP40

MACRO MUX2D0BWP40
    CLASS CORE ;
    FOREIGN MUX2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.074000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.215 1.505 1.030 ;
        RECT  1.310 0.215 1.425 0.315 ;
        RECT  1.355 0.930 1.425 1.030 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.420 0.790 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.540 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.540 1.375 ;
        RECT  1.120 1.000 1.220 1.375 ;
        RECT  0.340 1.145 1.120 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.205 0.515 1.285 0.925 ;
        RECT  0.790 0.850 1.205 0.925 ;
        RECT  0.940 0.195 1.040 0.275 ;
        RECT  0.940 0.710 1.040 0.780 ;
        RECT  0.860 0.195 0.940 0.780 ;
        RECT  0.770 0.995 0.940 1.075 ;
        RECT  0.690 0.335 0.790 0.925 ;
        RECT  0.580 0.995 0.770 1.065 ;
        RECT  0.510 0.315 0.580 0.800 ;
        RECT  0.510 0.870 0.580 1.065 ;
        RECT  0.125 0.870 0.510 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D0BWP40

MACRO MUX2D1BWP40
    CLASS CORE ;
    FOREIGN MUX2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.148000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.205 1.505 1.065 ;
        RECT  1.390 0.205 1.425 0.470 ;
        RECT  1.400 0.665 1.425 1.065 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.420 0.790 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.115 1.540 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.145 1.540 1.375 ;
        RECT  1.120 1.000 1.220 1.375 ;
        RECT  0.340 1.145 1.120 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.205 0.515 1.285 0.925 ;
        RECT  0.790 0.850 1.205 0.925 ;
        RECT  0.940 0.195 1.040 0.275 ;
        RECT  0.940 0.710 1.040 0.780 ;
        RECT  0.860 0.195 0.940 0.780 ;
        RECT  0.770 0.995 0.910 1.075 ;
        RECT  0.690 0.335 0.790 0.925 ;
        RECT  0.580 0.995 0.770 1.065 ;
        RECT  0.510 0.315 0.580 0.800 ;
        RECT  0.510 0.870 0.580 1.065 ;
        RECT  0.125 0.870 0.510 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D1BWP40

MACRO MUX2D2BWP40
    CLASS CORE ;
    FOREIGN MUX2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.385 1.925 0.775 ;
        RECT  1.715 0.385 1.850 0.465 ;
        RECT  1.725 0.695 1.850 0.775 ;
        RECT  1.645 0.695 1.725 1.060 ;
        RECT  1.645 0.200 1.715 0.465 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.036800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.840 -0.115 1.910 0.275 ;
        RECT  1.540 -0.115 1.840 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.250 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.840 0.965 1.910 1.375 ;
        RECT  1.540 1.145 1.840 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.565 0.545 1.750 0.615 ;
        RECT  1.490 0.545 1.565 0.925 ;
        RECT  1.085 0.850 1.490 0.925 ;
        RECT  1.225 0.195 1.360 0.275 ;
        RECT  1.225 0.710 1.350 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.155 0.195 1.225 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.010 0.310 1.085 0.925 ;
        RECT  0.830 0.320 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.320 0.830 0.390 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.320 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D2BWP40

MACRO MUX2D3BWP40
    CLASS CORE ;
    FOREIGN MUX2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.205 2.160 0.480 ;
        RECT  2.075 0.750 2.145 1.055 ;
        RECT  1.995 0.750 2.075 0.830 ;
        RECT  1.995 0.345 2.070 0.480 ;
        RECT  1.785 0.345 1.995 0.830 ;
        RECT  1.750 0.345 1.785 0.470 ;
        RECT  1.745 0.750 1.785 0.830 ;
        RECT  1.645 0.215 1.750 0.470 ;
        RECT  1.670 0.750 1.745 1.055 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.036800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.965 -0.115 2.240 0.115 ;
        RECT  1.855 -0.115 1.965 0.265 ;
        RECT  1.540 -0.115 1.855 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.250 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.955 1.145 2.240 1.375 ;
        RECT  1.865 0.965 1.955 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.070 0.205 2.160 0.480 ;
        RECT  2.075 0.750 2.145 1.055 ;
        RECT  2.065 0.750 2.075 0.830 ;
        RECT  2.065 0.345 2.070 0.480 ;
        RECT  1.645 0.215 1.715 0.470 ;
        RECT  1.670 0.750 1.715 1.055 ;
        RECT  1.600 0.545 1.705 0.615 ;
        RECT  1.520 0.545 1.600 0.925 ;
        RECT  1.085 0.850 1.520 0.925 ;
        RECT  1.225 0.195 1.360 0.275 ;
        RECT  1.225 0.710 1.360 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.155 0.195 1.225 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.010 0.280 1.085 0.925 ;
        RECT  0.830 0.320 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.320 0.830 0.390 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.320 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D3BWP40

MACRO MUX2D4BWP40
    CLASS CORE ;
    FOREIGN MUX2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.215 2.570 0.465 ;
        RECT  2.480 0.785 2.550 1.060 ;
        RECT  2.415 0.785 2.480 0.905 ;
        RECT  2.415 0.355 2.470 0.465 ;
        RECT  2.205 0.355 2.415 0.905 ;
        RECT  2.170 0.355 2.205 0.465 ;
        RECT  2.160 0.785 2.205 0.905 ;
        RECT  2.070 0.215 2.170 0.465 ;
        RECT  2.090 0.785 2.160 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.063200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.355 1.540 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.055200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 0.510 0.835 0.610 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.680 -0.115 2.750 0.455 ;
        RECT  2.385 -0.115 2.680 0.115 ;
        RECT  2.275 -0.115 2.385 0.265 ;
        RECT  1.970 -0.115 2.275 0.115 ;
        RECT  1.900 -0.115 1.970 0.425 ;
        RECT  1.610 -0.115 1.900 0.115 ;
        RECT  1.510 -0.115 1.610 0.275 ;
        RECT  0.780 -0.115 1.510 0.115 ;
        RECT  0.660 -0.115 0.780 0.295 ;
        RECT  0.370 -0.115 0.660 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.680 0.720 2.750 1.375 ;
        RECT  2.385 1.145 2.680 1.375 ;
        RECT  2.275 0.985 2.385 1.375 ;
        RECT  1.990 1.145 2.275 1.375 ;
        RECT  1.865 0.995 1.990 1.375 ;
        RECT  1.610 1.145 1.865 1.375 ;
        RECT  1.510 1.000 1.610 1.375 ;
        RECT  0.780 1.145 1.510 1.375 ;
        RECT  0.660 1.010 0.780 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.215 2.570 0.465 ;
        RECT  2.485 0.785 2.550 1.060 ;
        RECT  2.070 0.215 2.135 0.465 ;
        RECT  2.090 0.785 2.135 1.060 ;
        RECT  2.020 0.545 2.125 0.625 ;
        RECT  1.940 0.545 2.020 0.925 ;
        RECT  1.180 0.850 1.940 0.925 ;
        RECT  1.795 0.670 1.820 0.780 ;
        RECT  1.705 0.195 1.795 0.780 ;
        RECT  1.330 0.710 1.705 0.780 ;
        RECT  1.330 0.195 1.430 0.275 ;
        RECT  1.250 0.195 1.330 0.780 ;
        RECT  1.160 0.995 1.330 1.075 ;
        RECT  1.080 0.335 1.180 0.925 ;
        RECT  0.970 0.995 1.160 1.065 ;
        RECT  0.940 0.365 1.010 0.800 ;
        RECT  0.900 0.870 0.970 1.065 ;
        RECT  0.465 0.365 0.940 0.440 ;
        RECT  0.470 0.710 0.940 0.800 ;
        RECT  0.125 0.870 0.900 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D4BWP40

MACRO MUX2D6BWP40
    CLASS CORE ;
    FOREIGN MUX2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.215 2.970 0.465 ;
        RECT  2.880 0.770 2.950 1.060 ;
        RECT  2.695 0.770 2.880 0.905 ;
        RECT  2.695 0.355 2.870 0.465 ;
        RECT  2.570 0.355 2.695 0.905 ;
        RECT  2.560 0.215 2.570 0.905 ;
        RECT  2.485 0.215 2.560 1.060 ;
        RECT  2.470 0.215 2.485 0.465 ;
        RECT  2.480 0.770 2.485 1.060 ;
        RECT  2.160 0.770 2.480 0.905 ;
        RECT  2.170 0.355 2.470 0.465 ;
        RECT  2.070 0.215 2.170 0.465 ;
        RECT  2.090 0.770 2.160 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.063200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.355 1.535 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.055200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 0.495 0.845 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 -0.115 3.220 0.115 ;
        RECT  3.080 -0.115 3.150 0.465 ;
        RECT  2.750 -0.115 3.080 0.115 ;
        RECT  2.680 -0.115 2.750 0.265 ;
        RECT  2.385 -0.115 2.680 0.115 ;
        RECT  2.275 -0.115 2.385 0.265 ;
        RECT  1.970 -0.115 2.275 0.115 ;
        RECT  1.900 -0.115 1.970 0.430 ;
        RECT  1.610 -0.115 1.900 0.115 ;
        RECT  1.510 -0.115 1.610 0.275 ;
        RECT  0.780 -0.115 1.510 0.115 ;
        RECT  0.660 -0.115 0.780 0.280 ;
        RECT  0.370 -0.115 0.660 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.145 3.220 1.375 ;
        RECT  3.080 0.730 3.150 1.375 ;
        RECT  2.750 1.145 3.080 1.375 ;
        RECT  2.680 0.985 2.750 1.375 ;
        RECT  2.385 1.145 2.680 1.375 ;
        RECT  2.275 0.985 2.385 1.375 ;
        RECT  1.990 1.145 2.275 1.375 ;
        RECT  1.865 0.995 1.990 1.375 ;
        RECT  1.610 1.145 1.865 1.375 ;
        RECT  1.510 1.000 1.610 1.375 ;
        RECT  0.780 1.145 1.510 1.375 ;
        RECT  0.660 1.010 0.780 1.375 ;
        RECT  0.340 1.145 0.660 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.870 0.215 2.970 0.465 ;
        RECT  2.880 0.770 2.950 1.060 ;
        RECT  2.765 0.770 2.880 0.905 ;
        RECT  2.765 0.355 2.870 0.465 ;
        RECT  2.170 0.355 2.415 0.465 ;
        RECT  2.160 0.770 2.415 0.905 ;
        RECT  2.070 0.215 2.170 0.465 ;
        RECT  2.090 0.770 2.160 1.060 ;
        RECT  2.020 0.545 2.405 0.625 ;
        RECT  1.940 0.545 2.020 0.925 ;
        RECT  1.180 0.850 1.940 0.925 ;
        RECT  1.795 0.670 1.820 0.780 ;
        RECT  1.710 0.195 1.795 0.780 ;
        RECT  1.330 0.710 1.710 0.780 ;
        RECT  1.330 0.195 1.430 0.275 ;
        RECT  1.250 0.195 1.330 0.780 ;
        RECT  1.160 0.995 1.330 1.075 ;
        RECT  1.080 0.335 1.180 0.925 ;
        RECT  0.970 0.995 1.160 1.065 ;
        RECT  0.940 0.350 1.010 0.800 ;
        RECT  0.900 0.870 0.970 1.065 ;
        RECT  0.465 0.350 0.940 0.425 ;
        RECT  0.470 0.710 0.940 0.800 ;
        RECT  0.125 0.870 0.900 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D6BWP40

MACRO MUX2D8BWP40
    CLASS CORE ;
    FOREIGN MUX2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.710 0.215 4.810 0.465 ;
        RECT  4.720 0.770 4.790 1.060 ;
        RECT  4.400 0.770 4.720 0.905 ;
        RECT  4.410 0.355 4.710 0.465 ;
        RECT  4.310 0.215 4.410 0.465 ;
        RECT  4.330 0.770 4.400 1.060 ;
        RECT  4.235 0.770 4.330 0.905 ;
        RECT  4.235 0.355 4.310 0.465 ;
        RECT  4.030 0.355 4.235 0.905 ;
        RECT  4.025 0.215 4.030 0.905 ;
        RECT  3.930 0.215 4.025 0.465 ;
        RECT  4.010 0.770 4.025 0.905 ;
        RECT  3.940 0.770 4.010 1.060 ;
        RECT  3.620 0.770 3.940 0.905 ;
        RECT  3.630 0.355 3.930 0.465 ;
        RECT  3.530 0.215 3.630 0.465 ;
        RECT  3.550 0.770 3.620 1.060 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.280 0.765 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.094800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.495 3.075 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.099200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.495 1.515 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.920 -0.115 4.990 0.450 ;
        RECT  4.625 -0.115 4.920 0.115 ;
        RECT  4.515 -0.115 4.625 0.265 ;
        RECT  4.210 -0.115 4.515 0.115 ;
        RECT  4.140 -0.115 4.210 0.265 ;
        RECT  3.845 -0.115 4.140 0.115 ;
        RECT  3.735 -0.115 3.845 0.265 ;
        RECT  3.440 -0.115 3.735 0.115 ;
        RECT  3.340 -0.115 3.440 0.385 ;
        RECT  3.045 -0.115 3.340 0.115 ;
        RECT  2.945 -0.115 3.045 0.265 ;
        RECT  1.495 -0.115 2.945 0.115 ;
        RECT  1.375 -0.115 1.495 0.280 ;
        RECT  1.115 -0.115 1.375 0.115 ;
        RECT  0.995 -0.115 1.115 0.280 ;
        RECT  0.725 -0.115 0.995 0.115 ;
        RECT  0.605 -0.115 0.725 0.280 ;
        RECT  0.345 -0.115 0.605 0.115 ;
        RECT  0.225 -0.115 0.345 0.300 ;
        RECT  0.000 -0.115 0.225 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.920 0.720 4.990 1.375 ;
        RECT  4.625 1.145 4.920 1.375 ;
        RECT  4.515 0.985 4.625 1.375 ;
        RECT  4.230 1.145 4.515 1.375 ;
        RECT  4.105 0.995 4.230 1.375 ;
        RECT  3.845 1.145 4.105 1.375 ;
        RECT  3.735 0.985 3.845 1.375 ;
        RECT  3.440 1.145 3.735 1.375 ;
        RECT  3.340 1.000 3.440 1.375 ;
        RECT  3.045 1.145 3.340 1.375 ;
        RECT  2.945 1.000 3.045 1.375 ;
        RECT  1.495 1.145 2.945 1.375 ;
        RECT  1.375 1.010 1.495 1.375 ;
        RECT  1.065 1.145 1.375 1.375 ;
        RECT  0.945 1.010 1.065 1.375 ;
        RECT  0.555 1.145 0.945 1.375 ;
        RECT  0.435 1.010 0.555 1.375 ;
        RECT  0.340 1.145 0.435 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.710 0.215 4.810 0.465 ;
        RECT  4.720 0.770 4.790 1.060 ;
        RECT  4.400 0.770 4.720 0.905 ;
        RECT  4.410 0.355 4.710 0.465 ;
        RECT  4.310 0.215 4.410 0.465 ;
        RECT  4.330 0.770 4.400 1.060 ;
        RECT  4.305 0.770 4.330 0.905 ;
        RECT  4.305 0.355 4.310 0.465 ;
        RECT  3.930 0.215 3.955 0.465 ;
        RECT  3.940 0.770 3.955 1.060 ;
        RECT  3.620 0.770 3.940 0.905 ;
        RECT  3.630 0.355 3.930 0.465 ;
        RECT  3.530 0.215 3.630 0.465 ;
        RECT  3.550 0.770 3.620 1.060 ;
        RECT  3.480 0.545 3.915 0.625 ;
        RECT  3.400 0.545 3.480 0.925 ;
        RECT  2.240 0.855 3.400 0.925 ;
        RECT  3.230 0.670 3.255 0.780 ;
        RECT  3.145 0.345 3.230 0.780 ;
        RECT  2.370 0.345 3.145 0.415 ;
        RECT  2.325 0.710 3.145 0.780 ;
        RECT  2.240 0.195 2.690 0.265 ;
        RECT  1.685 0.995 2.415 1.065 ;
        RECT  2.170 0.195 2.240 0.925 ;
        RECT  1.765 0.195 2.170 0.265 ;
        RECT  1.765 0.855 2.170 0.925 ;
        RECT  2.010 0.350 2.080 0.785 ;
        RECT  0.410 0.350 2.010 0.425 ;
        RECT  0.675 0.710 2.010 0.785 ;
        RECT  1.615 0.870 1.685 1.065 ;
        RECT  0.125 0.870 1.615 0.940 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2D8BWP40

MACRO MUX2ND0BWP40
    CLASS CORE ;
    FOREIGN MUX2ND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.062000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.215 1.925 1.045 ;
        RECT  1.760 0.215 1.855 0.315 ;
        RECT  1.740 0.945 1.855 1.045 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.355 0.430 0.625 ;
        RECT  0.315 0.355 0.415 0.780 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 -0.115 1.960 0.115 ;
        RECT  1.570 -0.115 1.650 0.315 ;
        RECT  1.260 -0.115 1.570 0.115 ;
        RECT  1.160 -0.115 1.260 0.285 ;
        RECT  0.370 -0.115 1.160 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.145 1.960 1.375 ;
        RECT  1.575 0.925 1.645 1.375 ;
        RECT  1.250 1.145 1.575 1.375 ;
        RECT  1.170 0.980 1.250 1.375 ;
        RECT  0.340 1.145 1.170 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.605 0.395 1.675 0.845 ;
        RECT  1.465 0.395 1.605 0.465 ;
        RECT  1.465 0.775 1.605 0.845 ;
        RECT  1.395 0.210 1.465 0.465 ;
        RECT  1.395 0.775 1.465 0.915 ;
        RECT  1.275 0.545 1.400 0.620 ;
        RECT  1.205 0.545 1.275 0.910 ;
        RECT  0.780 0.840 1.205 0.910 ;
        RECT  0.940 0.700 1.070 0.770 ;
        RECT  0.940 0.205 1.060 0.275 ;
        RECT  0.790 0.995 0.960 1.075 ;
        RECT  0.860 0.205 0.940 0.770 ;
        RECT  0.580 0.995 0.790 1.065 ;
        RECT  0.700 0.325 0.780 0.910 ;
        RECT  0.530 0.335 0.600 0.780 ;
        RECT  0.510 0.850 0.580 1.065 ;
        RECT  0.500 0.335 0.530 0.455 ;
        RECT  0.485 0.685 0.530 0.780 ;
        RECT  0.125 0.850 0.510 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND0BWP40

MACRO MUX2ND1BWP40
    CLASS CORE ;
    FOREIGN MUX2ND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.148000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.195 1.925 1.065 ;
        RECT  1.790 0.195 1.855 0.460 ;
        RECT  1.820 0.665 1.855 1.065 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.355 0.430 0.625 ;
        RECT  0.315 0.355 0.415 0.780 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 -0.115 1.960 0.115 ;
        RECT  1.570 -0.115 1.650 0.315 ;
        RECT  1.260 -0.115 1.570 0.115 ;
        RECT  1.160 -0.115 1.260 0.275 ;
        RECT  0.370 -0.115 1.160 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.145 1.960 1.375 ;
        RECT  1.575 0.925 1.645 1.375 ;
        RECT  1.250 1.145 1.575 1.375 ;
        RECT  1.170 0.980 1.250 1.375 ;
        RECT  0.340 1.145 1.170 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.605 0.395 1.675 0.845 ;
        RECT  1.465 0.395 1.605 0.465 ;
        RECT  1.465 0.775 1.605 0.845 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        RECT  1.275 0.545 1.380 0.620 ;
        RECT  1.205 0.545 1.275 0.910 ;
        RECT  0.780 0.840 1.205 0.910 ;
        RECT  0.940 0.700 1.070 0.770 ;
        RECT  0.940 0.205 1.060 0.275 ;
        RECT  0.790 0.995 0.960 1.075 ;
        RECT  0.860 0.205 0.940 0.770 ;
        RECT  0.580 0.995 0.790 1.065 ;
        RECT  0.700 0.325 0.780 0.910 ;
        RECT  0.530 0.335 0.600 0.780 ;
        RECT  0.510 0.850 0.580 1.065 ;
        RECT  0.500 0.335 0.530 0.455 ;
        RECT  0.485 0.685 0.530 0.780 ;
        RECT  0.125 0.850 0.510 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND1BWP40

MACRO MUX2ND2BWP40
    CLASS CORE ;
    FOREIGN MUX2ND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.335 1.925 0.895 ;
        RECT  1.760 0.195 1.855 0.470 ;
        RECT  1.850 0.760 1.855 0.895 ;
        RECT  1.770 0.760 1.850 1.065 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.355 0.430 0.625 ;
        RECT  0.315 0.355 0.415 0.780 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.115 2.100 0.115 ;
        RECT  1.945 -0.115 2.055 0.250 ;
        RECT  1.650 -0.115 1.945 0.115 ;
        RECT  1.570 -0.115 1.650 0.315 ;
        RECT  1.260 -0.115 1.570 0.115 ;
        RECT  1.160 -0.115 1.260 0.275 ;
        RECT  0.370 -0.115 1.160 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 1.145 2.100 1.375 ;
        RECT  1.945 0.995 2.055 1.375 ;
        RECT  1.665 1.145 1.945 1.375 ;
        RECT  1.575 0.925 1.665 1.375 ;
        RECT  1.250 1.145 1.575 1.375 ;
        RECT  1.170 0.980 1.250 1.375 ;
        RECT  0.340 1.145 1.170 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.605 0.395 1.675 0.845 ;
        RECT  1.465 0.395 1.605 0.465 ;
        RECT  1.465 0.775 1.605 0.845 ;
        RECT  1.395 0.185 1.465 0.465 ;
        RECT  1.395 0.775 1.465 1.055 ;
        RECT  1.275 0.545 1.400 0.620 ;
        RECT  1.205 0.545 1.275 0.910 ;
        RECT  0.780 0.840 1.205 0.910 ;
        RECT  0.940 0.700 1.070 0.770 ;
        RECT  0.940 0.205 1.060 0.275 ;
        RECT  0.790 0.995 0.960 1.075 ;
        RECT  0.860 0.205 0.940 0.770 ;
        RECT  0.580 0.995 0.790 1.065 ;
        RECT  0.700 0.325 0.780 0.910 ;
        RECT  0.530 0.335 0.600 0.780 ;
        RECT  0.510 0.850 0.580 1.065 ;
        RECT  0.500 0.335 0.530 0.455 ;
        RECT  0.485 0.685 0.530 0.780 ;
        RECT  0.125 0.850 0.510 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND2BWP40

MACRO MUX2ND3BWP40
    CLASS CORE ;
    FOREIGN MUX2ND3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.224000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.110 0.195 2.205 0.470 ;
        RECT  2.105 0.760 2.205 1.060 ;
        RECT  1.955 0.335 2.110 0.470 ;
        RECT  1.955 0.760 2.105 0.875 ;
        RECT  1.830 0.335 1.955 0.875 ;
        RECT  1.805 0.335 1.830 0.470 ;
        RECT  1.800 0.760 1.830 0.875 ;
        RECT  1.715 0.195 1.805 0.470 ;
        RECT  1.715 0.760 1.800 1.060 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.355 1.115 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.415 0.355 0.430 0.625 ;
        RECT  0.315 0.355 0.415 0.780 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.115 2.240 0.115 ;
        RECT  1.890 -0.115 2.000 0.250 ;
        RECT  1.605 -0.115 1.890 0.115 ;
        RECT  1.525 -0.115 1.605 0.315 ;
        RECT  1.250 -0.115 1.525 0.115 ;
        RECT  1.150 -0.115 1.250 0.285 ;
        RECT  0.370 -0.115 1.150 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.145 2.240 1.375 ;
        RECT  1.890 0.995 2.000 1.375 ;
        RECT  1.600 1.145 1.890 1.375 ;
        RECT  1.530 0.925 1.600 1.375 ;
        RECT  1.230 1.145 1.530 1.375 ;
        RECT  1.150 0.980 1.230 1.375 ;
        RECT  0.340 1.145 1.150 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.560 0.395 1.630 0.845 ;
        RECT  1.420 0.395 1.560 0.465 ;
        RECT  1.420 0.775 1.560 0.845 ;
        RECT  1.350 0.185 1.420 0.465 ;
        RECT  1.350 0.775 1.420 1.055 ;
        RECT  1.275 0.545 1.355 0.620 ;
        RECT  1.205 0.545 1.275 0.910 ;
        RECT  0.780 0.840 1.205 0.910 ;
        RECT  0.940 0.700 1.070 0.770 ;
        RECT  0.940 0.205 1.060 0.275 ;
        RECT  0.790 0.995 0.960 1.075 ;
        RECT  0.860 0.205 0.940 0.770 ;
        RECT  0.580 0.995 0.790 1.065 ;
        RECT  0.700 0.325 0.780 0.910 ;
        RECT  0.530 0.335 0.600 0.780 ;
        RECT  0.510 0.850 0.580 1.065 ;
        RECT  0.500 0.335 0.530 0.455 ;
        RECT  0.485 0.685 0.530 0.780 ;
        RECT  0.125 0.850 0.510 0.920 ;
        RECT  0.105 0.215 0.140 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.215 0.105 1.030 ;
    END
END MUX2ND3BWP40

MACRO MUX2ND4BWP40
    CLASS CORE ;
    FOREIGN MUX2ND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.185 2.560 0.445 ;
        RECT  2.485 0.705 2.555 1.030 ;
        RECT  2.415 0.705 2.485 0.820 ;
        RECT  2.415 0.310 2.480 0.445 ;
        RECT  2.205 0.310 2.415 0.820 ;
        RECT  2.140 0.310 2.205 0.445 ;
        RECT  2.135 0.705 2.205 0.820 ;
        RECT  2.060 0.185 2.140 0.445 ;
        RECT  2.065 0.705 2.135 1.030 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.037200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.465 ;
        RECT  2.380 -0.115 2.670 0.115 ;
        RECT  2.260 -0.115 2.380 0.240 ;
        RECT  1.950 -0.115 2.260 0.115 ;
        RECT  1.880 -0.115 1.950 0.270 ;
        RECT  1.540 -0.115 1.880 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.250 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.695 2.750 1.375 ;
        RECT  2.380 1.145 2.670 1.375 ;
        RECT  2.260 0.890 2.380 1.375 ;
        RECT  1.950 1.145 2.260 1.375 ;
        RECT  1.880 0.965 1.950 1.375 ;
        RECT  1.540 1.145 1.880 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.185 2.560 0.445 ;
        RECT  2.485 0.705 2.555 1.030 ;
        RECT  2.060 0.185 2.135 0.445 ;
        RECT  2.065 0.705 2.135 1.030 ;
        RECT  1.965 0.545 2.110 0.615 ;
        RECT  1.890 0.385 1.965 0.805 ;
        RECT  1.720 0.385 1.890 0.465 ;
        RECT  1.735 0.725 1.890 0.805 ;
        RECT  1.580 0.545 1.745 0.615 ;
        RECT  1.650 0.725 1.735 1.060 ;
        RECT  1.645 0.195 1.720 0.465 ;
        RECT  1.500 0.545 1.580 0.925 ;
        RECT  1.080 0.850 1.500 0.925 ;
        RECT  1.220 0.195 1.360 0.275 ;
        RECT  1.220 0.710 1.360 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.150 0.195 1.220 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.010 0.255 1.080 0.925 ;
        RECT  0.830 0.320 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.320 0.830 0.390 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.320 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2ND4BWP40

MACRO MUX2ND6BWP40
    CLASS CORE ;
    FOREIGN MUX2ND6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.860 0.185 2.940 0.445 ;
        RECT  2.865 0.705 2.935 1.030 ;
        RECT  2.555 0.705 2.865 0.820 ;
        RECT  2.560 0.310 2.860 0.445 ;
        RECT  2.555 0.185 2.560 0.445 ;
        RECT  2.485 0.185 2.555 1.030 ;
        RECT  2.480 0.185 2.485 0.820 ;
        RECT  2.345 0.310 2.480 0.820 ;
        RECT  2.140 0.310 2.345 0.445 ;
        RECT  2.135 0.705 2.345 0.820 ;
        RECT  2.060 0.185 2.140 0.445 ;
        RECT  2.065 0.705 2.135 1.030 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.037200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 -0.115 3.220 0.115 ;
        RECT  3.030 -0.115 3.150 0.240 ;
        RECT  2.770 -0.115 3.030 0.115 ;
        RECT  2.650 -0.115 2.770 0.240 ;
        RECT  2.380 -0.115 2.650 0.115 ;
        RECT  2.260 -0.115 2.380 0.240 ;
        RECT  1.970 -0.115 2.260 0.115 ;
        RECT  1.850 -0.115 1.970 0.255 ;
        RECT  1.540 -0.115 1.850 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.260 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.145 3.220 1.375 ;
        RECT  3.030 0.750 3.150 1.375 ;
        RECT  2.770 1.145 3.030 1.375 ;
        RECT  2.650 0.890 2.770 1.375 ;
        RECT  2.380 1.145 2.650 1.375 ;
        RECT  2.260 0.890 2.380 1.375 ;
        RECT  1.950 1.145 2.260 1.375 ;
        RECT  1.865 1.005 1.950 1.375 ;
        RECT  1.540 1.145 1.865 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.860 0.185 2.940 0.445 ;
        RECT  2.865 0.705 2.935 1.030 ;
        RECT  2.625 0.705 2.865 0.820 ;
        RECT  2.625 0.310 2.860 0.445 ;
        RECT  2.140 0.310 2.275 0.445 ;
        RECT  2.135 0.705 2.275 0.820 ;
        RECT  2.060 0.185 2.140 0.445 ;
        RECT  2.065 0.705 2.135 1.030 ;
        RECT  1.965 0.545 2.265 0.615 ;
        RECT  1.885 0.375 1.965 0.830 ;
        RECT  1.720 0.375 1.885 0.455 ;
        RECT  1.730 0.750 1.885 0.830 ;
        RECT  1.580 0.545 1.730 0.615 ;
        RECT  1.650 0.750 1.730 1.060 ;
        RECT  1.640 0.195 1.720 0.455 ;
        RECT  1.500 0.545 1.580 0.925 ;
        RECT  1.085 0.850 1.500 0.925 ;
        RECT  1.225 0.195 1.360 0.275 ;
        RECT  1.225 0.710 1.360 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.155 0.195 1.225 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.010 0.310 1.085 0.925 ;
        RECT  0.830 0.330 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.330 0.830 0.400 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.330 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2ND6BWP40

MACRO MUX2ND8BWP40
    CLASS CORE ;
    FOREIGN MUX2ND8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.585 0.185 3.675 0.445 ;
        RECT  3.590 0.705 3.660 1.030 ;
        RECT  3.280 0.705 3.590 0.820 ;
        RECT  3.285 0.310 3.585 0.445 ;
        RECT  3.205 0.185 3.285 0.445 ;
        RECT  3.210 0.705 3.280 1.030 ;
        RECT  3.115 0.705 3.210 0.820 ;
        RECT  3.115 0.310 3.205 0.445 ;
        RECT  2.905 0.310 3.115 0.820 ;
        RECT  2.825 0.185 2.905 0.445 ;
        RECT  2.830 0.705 2.905 1.045 ;
        RECT  2.520 0.705 2.830 0.820 ;
        RECT  2.525 0.310 2.825 0.445 ;
        RECT  2.445 0.185 2.525 0.445 ;
        RECT  2.450 0.705 2.520 1.030 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.395 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.037200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.470 0.685 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.795 -0.115 3.870 0.455 ;
        RECT  3.495 -0.115 3.795 0.115 ;
        RECT  3.375 -0.115 3.495 0.240 ;
        RECT  3.115 -0.115 3.375 0.115 ;
        RECT  2.995 -0.115 3.115 0.240 ;
        RECT  2.735 -0.115 2.995 0.115 ;
        RECT  2.615 -0.115 2.735 0.240 ;
        RECT  2.345 -0.115 2.615 0.115 ;
        RECT  2.245 -0.115 2.345 0.415 ;
        RECT  1.970 -0.115 2.245 0.115 ;
        RECT  1.885 -0.115 1.970 0.295 ;
        RECT  1.540 -0.115 1.885 0.115 ;
        RECT  1.440 -0.115 1.540 0.275 ;
        RECT  0.710 -0.115 1.440 0.115 ;
        RECT  0.590 -0.115 0.710 0.250 ;
        RECT  0.340 -0.115 0.590 0.115 ;
        RECT  0.220 -0.115 0.340 0.300 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.145 3.920 1.375 ;
        RECT  3.785 0.720 3.880 1.375 ;
        RECT  3.500 1.145 3.785 1.375 ;
        RECT  3.375 0.890 3.500 1.375 ;
        RECT  3.120 1.145 3.375 1.375 ;
        RECT  2.995 0.890 3.120 1.375 ;
        RECT  2.735 1.145 2.995 1.375 ;
        RECT  2.615 0.890 2.735 1.375 ;
        RECT  2.345 1.145 2.615 1.375 ;
        RECT  2.245 0.730 2.345 1.375 ;
        RECT  1.950 1.145 2.245 1.375 ;
        RECT  1.880 0.965 1.950 1.375 ;
        RECT  1.540 1.145 1.880 1.375 ;
        RECT  1.440 1.000 1.540 1.375 ;
        RECT  0.710 1.145 1.440 1.375 ;
        RECT  0.590 1.010 0.710 1.375 ;
        RECT  0.340 1.145 0.590 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.585 0.185 3.675 0.445 ;
        RECT  3.590 0.705 3.660 1.030 ;
        RECT  3.280 0.705 3.590 0.820 ;
        RECT  3.285 0.310 3.585 0.445 ;
        RECT  3.205 0.185 3.285 0.445 ;
        RECT  3.210 0.705 3.280 1.030 ;
        RECT  3.185 0.705 3.210 0.820 ;
        RECT  3.185 0.310 3.205 0.445 ;
        RECT  2.825 0.185 2.835 0.445 ;
        RECT  2.830 0.705 2.835 1.045 ;
        RECT  2.520 0.705 2.830 0.820 ;
        RECT  2.525 0.310 2.825 0.445 ;
        RECT  2.445 0.185 2.525 0.445 ;
        RECT  2.450 0.705 2.520 1.030 ;
        RECT  2.160 0.545 2.725 0.615 ;
        RECT  2.150 0.545 2.160 1.060 ;
        RECT  2.080 0.195 2.150 1.060 ;
        RECT  2.075 0.375 2.080 1.060 ;
        RECT  2.045 0.375 2.075 0.835 ;
        RECT  1.740 0.375 2.045 0.455 ;
        RECT  1.750 0.755 2.045 0.835 ;
        RECT  1.600 0.545 1.890 0.615 ;
        RECT  1.670 0.755 1.750 1.060 ;
        RECT  1.660 0.195 1.740 0.455 ;
        RECT  1.520 0.545 1.600 0.925 ;
        RECT  1.085 0.850 1.520 0.925 ;
        RECT  1.225 0.195 1.360 0.275 ;
        RECT  1.225 0.710 1.360 0.780 ;
        RECT  1.090 0.995 1.260 1.075 ;
        RECT  1.155 0.195 1.225 0.780 ;
        RECT  0.900 0.995 1.090 1.065 ;
        RECT  1.015 0.315 1.085 0.925 ;
        RECT  0.830 0.320 0.900 0.800 ;
        RECT  0.830 0.870 0.900 1.065 ;
        RECT  0.500 0.320 0.830 0.390 ;
        RECT  0.125 0.870 0.830 0.940 ;
        RECT  0.420 0.320 0.500 0.800 ;
        RECT  0.405 0.700 0.420 0.800 ;
        RECT  0.105 0.215 0.125 0.335 ;
        RECT  0.105 0.870 0.125 1.040 ;
        RECT  0.035 0.215 0.105 1.040 ;
    END
END MUX2ND8BWP40

MACRO MUX3D0BWP40
    CLASS CORE ;
    FOREIGN MUX3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.052500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.215 2.485 1.045 ;
        RECT  2.390 0.215 2.415 0.420 ;
        RECT  2.335 0.970 2.415 1.045 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.260 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.090 0.775 2.205 0.905 ;
        RECT  1.990 0.495 2.090 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.355 1.085 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.015600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.440 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.260 0.135 ;
        RECT  1.220 -0.115 2.140 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.140 1.005 2.260 1.375 ;
        RECT  1.230 1.145 2.140 1.375 ;
        RECT  1.110 1.115 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.295 0.520 2.315 0.640 ;
        RECT  2.225 0.205 2.295 0.640 ;
        RECT  1.780 0.205 2.225 0.275 ;
        RECT  1.920 0.350 2.030 0.420 ;
        RECT  1.920 0.985 2.030 1.065 ;
        RECT  1.850 0.350 1.920 1.065 ;
        RECT  1.710 0.205 1.780 1.045 ;
        RECT  1.560 0.320 1.630 1.045 ;
        RECT  1.520 0.320 1.560 0.480 ;
        RECT  1.135 0.975 1.560 1.045 ;
        RECT  1.450 0.570 1.490 0.690 ;
        RECT  1.380 0.230 1.450 0.905 ;
        RECT  1.310 0.230 1.380 0.300 ;
        RECT  1.280 0.835 1.380 0.905 ;
        RECT  1.045 0.845 1.135 1.045 ;
        RECT  0.780 0.845 1.045 0.915 ;
        RECT  0.920 0.705 1.030 0.775 ;
        RECT  0.920 0.195 1.015 0.275 ;
        RECT  0.770 0.985 0.940 1.075 ;
        RECT  0.850 0.195 0.920 0.775 ;
        RECT  0.700 0.325 0.780 0.915 ;
        RECT  0.550 0.985 0.770 1.055 ;
        RECT  0.650 0.835 0.700 0.915 ;
        RECT  0.520 0.325 0.600 0.770 ;
        RECT  0.480 0.850 0.550 1.055 ;
        RECT  0.480 0.700 0.520 0.770 ;
        RECT  0.125 0.850 0.480 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D0BWP40

MACRO MUX3D1BWP40
    CLASS CORE ;
    FOREIGN MUX3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.097500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.195 2.485 1.065 ;
        RECT  2.380 0.195 2.415 0.465 ;
        RECT  2.380 0.675 2.415 1.065 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.260 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.100 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.029800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.355 1.085 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.440 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.260 0.135 ;
        RECT  1.220 -0.115 2.140 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.145 2.520 1.375 ;
        RECT  2.170 0.700 2.240 1.375 ;
        RECT  1.230 1.145 2.170 1.375 ;
        RECT  1.110 1.115 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 0.520 2.335 0.615 ;
        RECT  2.210 0.205 2.280 0.615 ;
        RECT  1.780 0.205 2.210 0.275 ;
        RECT  1.920 0.350 2.030 0.420 ;
        RECT  1.920 0.985 2.030 1.065 ;
        RECT  1.850 0.350 1.920 1.065 ;
        RECT  1.710 0.205 1.780 1.045 ;
        RECT  1.560 0.320 1.630 1.045 ;
        RECT  1.520 0.320 1.560 0.480 ;
        RECT  1.135 0.975 1.560 1.045 ;
        RECT  1.450 0.570 1.490 0.690 ;
        RECT  1.380 0.230 1.450 0.905 ;
        RECT  1.310 0.230 1.380 0.300 ;
        RECT  1.280 0.835 1.380 0.905 ;
        RECT  1.045 0.845 1.135 1.045 ;
        RECT  0.780 0.845 1.045 0.915 ;
        RECT  0.920 0.705 1.030 0.775 ;
        RECT  0.920 0.195 1.015 0.275 ;
        RECT  0.770 0.985 0.940 1.075 ;
        RECT  0.850 0.195 0.920 0.775 ;
        RECT  0.700 0.325 0.780 0.915 ;
        RECT  0.550 0.985 0.770 1.055 ;
        RECT  0.650 0.835 0.700 0.915 ;
        RECT  0.520 0.325 0.600 0.770 ;
        RECT  0.480 0.850 0.550 1.055 ;
        RECT  0.480 0.700 0.520 0.770 ;
        RECT  0.125 0.850 0.480 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D1BWP40

MACRO MUX3D2BWP40
    CLASS CORE ;
    FOREIGN MUX3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.330 3.045 0.770 ;
        RECT  2.840 0.330 2.955 0.455 ;
        RECT  2.860 0.695 2.955 0.770 ;
        RECT  2.740 0.695 2.860 1.065 ;
        RECT  2.760 0.195 2.840 0.455 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.680 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.495 2.485 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.029800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.355 1.505 0.625 ;
        RECT  1.385 0.505 1.410 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.036400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.355 0.820 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 -0.115 3.080 0.115 ;
        RECT  2.930 -0.115 3.045 0.255 ;
        RECT  2.640 -0.115 2.930 0.115 ;
        RECT  2.520 -0.115 2.640 0.135 ;
        RECT  1.600 -0.115 2.520 0.115 ;
        RECT  1.500 -0.115 1.600 0.275 ;
        RECT  0.770 -0.115 1.500 0.115 ;
        RECT  0.650 -0.115 0.770 0.280 ;
        RECT  0.370 -0.115 0.650 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.945 0.850 3.030 1.375 ;
        RECT  2.635 1.145 2.945 1.375 ;
        RECT  2.565 0.735 2.635 1.375 ;
        RECT  1.610 1.145 2.565 1.375 ;
        RECT  1.490 1.115 1.610 1.375 ;
        RECT  0.770 1.145 1.490 1.375 ;
        RECT  0.650 0.990 0.770 1.375 ;
        RECT  0.340 1.145 0.650 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.675 0.545 2.850 0.615 ;
        RECT  2.605 0.205 2.675 0.615 ;
        RECT  2.160 0.205 2.605 0.275 ;
        RECT  2.300 0.350 2.410 0.420 ;
        RECT  2.300 0.985 2.410 1.065 ;
        RECT  2.230 0.350 2.300 1.065 ;
        RECT  2.090 0.205 2.160 1.045 ;
        RECT  1.940 0.320 2.010 1.045 ;
        RECT  1.900 0.320 1.940 0.480 ;
        RECT  1.515 0.975 1.940 1.045 ;
        RECT  1.830 0.570 1.870 0.690 ;
        RECT  1.760 0.200 1.830 0.905 ;
        RECT  1.690 0.200 1.760 0.270 ;
        RECT  1.660 0.835 1.760 0.905 ;
        RECT  1.425 0.845 1.515 1.045 ;
        RECT  1.160 0.845 1.425 0.915 ;
        RECT  1.300 0.705 1.410 0.775 ;
        RECT  1.300 0.195 1.395 0.275 ;
        RECT  1.150 0.985 1.320 1.075 ;
        RECT  1.230 0.195 1.300 0.775 ;
        RECT  1.080 0.325 1.160 0.915 ;
        RECT  0.930 0.985 1.150 1.055 ;
        RECT  1.030 0.835 1.080 0.915 ;
        RECT  0.900 0.325 0.980 0.770 ;
        RECT  0.860 0.850 0.930 1.055 ;
        RECT  0.515 0.700 0.900 0.770 ;
        RECT  0.125 0.850 0.860 0.920 ;
        RECT  0.515 0.340 0.545 0.470 ;
        RECT  0.445 0.340 0.515 0.770 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D2BWP40

MACRO MUX3D4BWP40
    CLASS CORE ;
    FOREIGN MUX3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.260 0.720 4.360 1.010 ;
        RECT  4.235 0.195 4.355 0.475 ;
        RECT  4.235 0.720 4.260 0.820 ;
        RECT  4.025 0.365 4.235 0.820 ;
        RECT  3.965 0.365 4.025 0.455 ;
        RECT  3.955 0.715 4.025 0.820 ;
        RECT  3.865 0.195 3.965 0.455 ;
        RECT  3.870 0.715 3.955 1.010 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.415 2.490 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.465 0.765 ;
        RECT  3.195 0.495 3.395 0.630 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.059600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.505 2.275 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.061200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.785 0.500 1.240 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.535 -0.115 4.620 0.115 ;
        RECT  4.445 -0.115 4.535 0.450 ;
        RECT  4.165 -0.115 4.445 0.115 ;
        RECT  4.050 -0.115 4.165 0.285 ;
        RECT  3.790 -0.115 4.050 0.115 ;
        RECT  3.670 -0.115 3.790 0.135 ;
        RECT  3.420 -0.115 3.670 0.115 ;
        RECT  3.300 -0.115 3.420 0.135 ;
        RECT  2.410 -0.115 3.300 0.115 ;
        RECT  2.310 -0.115 2.410 0.275 ;
        RECT  1.980 -0.115 2.310 0.115 ;
        RECT  1.880 -0.115 1.980 0.275 ;
        RECT  1.190 -0.115 1.880 0.115 ;
        RECT  1.070 -0.115 1.190 0.280 ;
        RECT  0.770 -0.115 1.070 0.115 ;
        RECT  0.650 -0.115 0.770 0.280 ;
        RECT  0.370 -0.115 0.650 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.575 1.145 4.620 1.375 ;
        RECT  4.485 0.715 4.575 1.375 ;
        RECT  4.170 1.145 4.485 1.375 ;
        RECT  4.050 0.965 4.170 1.375 ;
        RECT  3.780 1.145 4.050 1.375 ;
        RECT  3.690 0.790 3.780 1.375 ;
        RECT  3.400 1.145 3.690 1.375 ;
        RECT  3.320 1.005 3.400 1.375 ;
        RECT  2.420 1.145 3.320 1.375 ;
        RECT  2.300 1.115 2.420 1.375 ;
        RECT  1.990 1.145 2.300 1.375 ;
        RECT  1.870 1.005 1.990 1.375 ;
        RECT  1.120 1.145 1.870 1.375 ;
        RECT  1.000 0.990 1.120 1.375 ;
        RECT  0.570 1.145 1.000 1.375 ;
        RECT  0.450 0.990 0.570 1.375 ;
        RECT  0.340 1.145 0.450 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.720 4.360 1.010 ;
        RECT  4.305 0.195 4.355 0.475 ;
        RECT  3.865 0.195 3.955 0.455 ;
        RECT  3.870 0.715 3.955 1.010 ;
        RECT  3.795 0.545 3.925 0.615 ;
        RECT  3.725 0.205 3.795 0.615 ;
        RECT  2.970 0.205 3.725 0.275 ;
        RECT  3.110 0.350 3.620 0.420 ;
        RECT  3.505 0.845 3.590 1.025 ;
        RECT  3.110 0.845 3.505 0.925 ;
        RECT  3.040 0.350 3.110 0.925 ;
        RECT  2.900 0.205 2.970 1.045 ;
        RECT  2.750 0.320 2.820 1.045 ;
        RECT  2.710 0.320 2.750 0.480 ;
        RECT  2.325 0.975 2.750 1.045 ;
        RECT  2.640 0.570 2.680 0.690 ;
        RECT  2.570 0.230 2.640 0.905 ;
        RECT  2.500 0.230 2.570 0.300 ;
        RECT  2.470 0.835 2.570 0.905 ;
        RECT  2.215 0.845 2.325 1.045 ;
        RECT  1.580 0.845 2.215 0.915 ;
        RECT  1.860 0.705 2.200 0.775 ;
        RECT  2.120 0.195 2.185 0.275 ;
        RECT  2.050 0.195 2.120 0.425 ;
        RECT  1.810 0.350 2.050 0.425 ;
        RECT  1.785 0.660 1.860 0.775 ;
        RECT  1.785 0.230 1.810 0.425 ;
        RECT  1.705 0.230 1.785 0.775 ;
        RECT  1.570 0.985 1.740 1.075 ;
        RECT  1.500 0.325 1.580 0.915 ;
        RECT  1.350 0.985 1.570 1.055 ;
        RECT  1.450 0.835 1.500 0.915 ;
        RECT  1.320 0.325 1.400 0.770 ;
        RECT  1.280 0.850 1.350 1.055 ;
        RECT  0.575 0.350 1.320 0.430 ;
        RECT  0.635 0.700 1.320 0.770 ;
        RECT  0.125 0.850 1.280 0.920 ;
        RECT  0.445 0.350 0.575 0.470 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3D4BWP40

MACRO MUX3ND0BWP40
    CLASS CORE ;
    FOREIGN MUX3ND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.058000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.675 0.185 2.765 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.355 1.275 0.655 ;
        RECT  1.155 0.355 1.230 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.440 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.100 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.355 1.085 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.015600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.440 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.115 2.800 0.115 ;
        RECT  2.450 -0.115 2.530 0.300 ;
        RECT  2.170 -0.115 2.450 0.115 ;
        RECT  2.070 -0.115 2.170 0.275 ;
        RECT  1.210 -0.115 2.070 0.115 ;
        RECT  1.110 -0.115 1.210 0.285 ;
        RECT  0.370 -0.115 1.110 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.145 2.800 1.375 ;
        RECT  2.430 1.005 2.550 1.375 ;
        RECT  2.180 1.145 2.430 1.375 ;
        RECT  2.060 1.030 2.180 1.375 ;
        RECT  1.230 1.145 2.060 1.375 ;
        RECT  1.110 1.115 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.380 2.565 0.930 ;
        RECT  2.350 0.380 2.490 0.450 ;
        RECT  2.345 0.860 2.490 0.930 ;
        RECT  2.250 0.235 2.350 0.450 ;
        RECT  2.275 0.860 2.345 1.020 ;
        RECT  2.220 0.520 2.290 0.780 ;
        RECT  2.190 0.710 2.220 0.780 ;
        RECT  2.120 0.710 2.190 0.960 ;
        RECT  1.790 0.890 2.120 0.960 ;
        RECT  1.915 0.750 2.010 0.820 ;
        RECT  1.915 0.205 1.990 0.275 ;
        RECT  1.845 0.205 1.915 0.820 ;
        RECT  1.770 0.890 1.790 1.045 ;
        RECT  1.700 0.285 1.770 1.045 ;
        RECT  1.560 0.320 1.630 1.045 ;
        RECT  1.500 0.320 1.560 0.480 ;
        RECT  1.135 0.975 1.560 1.045 ;
        RECT  1.430 0.570 1.490 0.690 ;
        RECT  1.360 0.210 1.430 0.905 ;
        RECT  1.290 0.210 1.360 0.280 ;
        RECT  1.310 0.835 1.360 0.905 ;
        RECT  1.045 0.845 1.135 1.045 ;
        RECT  0.780 0.845 1.045 0.915 ;
        RECT  0.920 0.705 1.030 0.775 ;
        RECT  0.920 0.195 1.015 0.275 ;
        RECT  0.770 0.985 0.940 1.075 ;
        RECT  0.850 0.195 0.920 0.775 ;
        RECT  0.700 0.325 0.780 0.915 ;
        RECT  0.550 0.985 0.770 1.055 ;
        RECT  0.650 0.835 0.700 0.915 ;
        RECT  0.520 0.325 0.600 0.770 ;
        RECT  0.480 0.850 0.550 1.055 ;
        RECT  0.480 0.700 0.520 0.770 ;
        RECT  0.125 0.850 0.480 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND0BWP40

MACRO MUX3ND1BWP40
    CLASS CORE ;
    FOREIGN MUX3ND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.116000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.675 0.185 2.765 1.065 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.355 1.275 0.655 ;
        RECT  1.155 0.355 1.230 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.440 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.355 2.100 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.030600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.355 1.085 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.440 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.530 -0.115 2.800 0.115 ;
        RECT  2.450 -0.115 2.530 0.300 ;
        RECT  2.170 -0.115 2.450 0.115 ;
        RECT  2.070 -0.115 2.170 0.275 ;
        RECT  1.210 -0.115 2.070 0.115 ;
        RECT  1.110 -0.115 1.210 0.275 ;
        RECT  0.370 -0.115 1.110 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.145 2.800 1.375 ;
        RECT  2.430 1.005 2.550 1.375 ;
        RECT  2.180 1.145 2.430 1.375 ;
        RECT  2.060 1.030 2.180 1.375 ;
        RECT  1.230 1.145 2.060 1.375 ;
        RECT  1.110 1.115 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.490 0.380 2.565 0.930 ;
        RECT  2.350 0.380 2.490 0.450 ;
        RECT  2.345 0.860 2.490 0.930 ;
        RECT  2.250 0.190 2.350 0.450 ;
        RECT  2.275 0.860 2.345 1.020 ;
        RECT  2.190 0.520 2.280 0.780 ;
        RECT  2.120 0.710 2.190 0.960 ;
        RECT  1.790 0.890 2.120 0.960 ;
        RECT  1.915 0.750 2.010 0.820 ;
        RECT  1.915 0.210 1.990 0.280 ;
        RECT  1.845 0.210 1.915 0.820 ;
        RECT  1.770 0.890 1.790 1.045 ;
        RECT  1.700 0.285 1.770 1.045 ;
        RECT  1.560 0.320 1.630 1.045 ;
        RECT  1.500 0.320 1.560 0.480 ;
        RECT  1.135 0.975 1.560 1.045 ;
        RECT  1.430 0.570 1.490 0.690 ;
        RECT  1.360 0.205 1.430 0.905 ;
        RECT  1.280 0.205 1.360 0.275 ;
        RECT  1.310 0.835 1.360 0.905 ;
        RECT  1.045 0.845 1.135 1.045 ;
        RECT  0.780 0.845 1.045 0.915 ;
        RECT  0.920 0.705 1.030 0.775 ;
        RECT  0.920 0.195 1.015 0.275 ;
        RECT  0.770 0.985 0.940 1.075 ;
        RECT  0.850 0.195 0.920 0.775 ;
        RECT  0.700 0.325 0.780 0.915 ;
        RECT  0.550 0.985 0.770 1.055 ;
        RECT  0.650 0.835 0.700 0.915 ;
        RECT  0.520 0.325 0.600 0.770 ;
        RECT  0.480 0.850 0.550 1.055 ;
        RECT  0.480 0.700 0.520 0.770 ;
        RECT  0.125 0.850 0.480 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND1BWP40

MACRO MUX3ND2BWP40
    CLASS CORE ;
    FOREIGN MUX3ND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.355 2.905 0.815 ;
        RECT  2.835 0.185 2.840 0.815 ;
        RECT  2.760 0.185 2.835 0.445 ;
        RECT  2.765 0.735 2.835 1.035 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.260 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.495 2.090 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.030200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.355 1.085 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.440 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.285 ;
        RECT  2.660 -0.115 2.950 0.115 ;
        RECT  2.560 -0.115 2.660 0.415 ;
        RECT  2.260 -0.115 2.560 0.115 ;
        RECT  2.140 -0.115 2.260 0.135 ;
        RECT  1.220 -0.115 2.140 0.115 ;
        RECT  1.120 -0.115 1.220 0.275 ;
        RECT  0.370 -0.115 1.120 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.910 3.030 1.375 ;
        RECT  2.660 1.145 2.950 1.375 ;
        RECT  2.560 0.845 2.660 1.375 ;
        RECT  2.240 1.145 2.560 1.375 ;
        RECT  2.160 0.730 2.240 1.375 ;
        RECT  1.230 1.145 2.160 1.375 ;
        RECT  1.110 1.115 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.485 0.545 2.765 0.615 ;
        RECT  2.415 0.195 2.485 1.060 ;
        RECT  2.380 0.195 2.415 0.450 ;
        RECT  2.380 0.760 2.415 1.060 ;
        RECT  2.295 0.525 2.345 0.640 ;
        RECT  2.225 0.205 2.295 0.640 ;
        RECT  1.780 0.205 2.225 0.275 ;
        RECT  1.920 0.350 2.030 0.420 ;
        RECT  1.920 0.985 2.030 1.065 ;
        RECT  1.850 0.350 1.920 1.065 ;
        RECT  1.710 0.205 1.780 1.045 ;
        RECT  1.560 0.320 1.630 1.045 ;
        RECT  1.520 0.320 1.560 0.480 ;
        RECT  1.135 0.975 1.560 1.045 ;
        RECT  1.450 0.570 1.490 0.690 ;
        RECT  1.380 0.230 1.450 0.905 ;
        RECT  1.310 0.230 1.380 0.300 ;
        RECT  1.280 0.835 1.380 0.905 ;
        RECT  1.045 0.845 1.135 1.045 ;
        RECT  0.780 0.845 1.045 0.915 ;
        RECT  0.920 0.705 1.030 0.775 ;
        RECT  0.920 0.195 1.015 0.275 ;
        RECT  0.770 0.985 0.940 1.075 ;
        RECT  0.850 0.195 0.920 0.775 ;
        RECT  0.700 0.325 0.780 0.915 ;
        RECT  0.550 0.985 0.770 1.055 ;
        RECT  0.650 0.835 0.700 0.915 ;
        RECT  0.520 0.325 0.600 0.770 ;
        RECT  0.480 0.850 0.550 1.055 ;
        RECT  0.480 0.700 0.520 0.770 ;
        RECT  0.125 0.850 0.480 0.920 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND2BWP40

MACRO MUX3ND4BWP40
    CLASS CORE ;
    FOREIGN MUX3ND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.600 0.185 3.680 0.445 ;
        RECT  3.605 0.705 3.675 1.030 ;
        RECT  3.535 0.705 3.605 0.820 ;
        RECT  3.535 0.310 3.600 0.445 ;
        RECT  3.325 0.310 3.535 0.820 ;
        RECT  3.260 0.310 3.325 0.445 ;
        RECT  3.255 0.705 3.325 0.820 ;
        RECT  3.180 0.185 3.260 0.445 ;
        RECT  3.165 0.705 3.255 1.030 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.355 1.680 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.450 0.245 0.770 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.495 2.485 0.905 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.029800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.355 1.505 0.625 ;
        RECT  1.385 0.505 1.410 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.036400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.355 0.820 0.630 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 -0.115 3.920 0.115 ;
        RECT  3.790 -0.115 3.870 0.465 ;
        RECT  3.500 -0.115 3.790 0.115 ;
        RECT  3.380 -0.115 3.500 0.240 ;
        RECT  3.045 -0.115 3.380 0.115 ;
        RECT  2.930 -0.115 3.045 0.285 ;
        RECT  2.640 -0.115 2.930 0.115 ;
        RECT  2.520 -0.115 2.640 0.135 ;
        RECT  1.600 -0.115 2.520 0.115 ;
        RECT  1.500 -0.115 1.600 0.275 ;
        RECT  0.770 -0.115 1.500 0.115 ;
        RECT  0.650 -0.115 0.770 0.280 ;
        RECT  0.370 -0.115 0.650 0.115 ;
        RECT  0.250 -0.115 0.370 0.275 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.145 3.920 1.375 ;
        RECT  3.790 0.695 3.870 1.375 ;
        RECT  3.500 1.145 3.790 1.375 ;
        RECT  3.380 0.890 3.500 1.375 ;
        RECT  3.030 1.145 3.380 1.375 ;
        RECT  2.945 0.875 3.030 1.375 ;
        RECT  2.640 1.145 2.945 1.375 ;
        RECT  2.555 0.730 2.640 1.375 ;
        RECT  1.610 1.145 2.555 1.375 ;
        RECT  1.490 1.115 1.610 1.375 ;
        RECT  0.770 1.145 1.490 1.375 ;
        RECT  0.650 0.990 0.770 1.375 ;
        RECT  0.340 1.145 0.650 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.185 3.680 0.445 ;
        RECT  3.605 0.705 3.675 1.030 ;
        RECT  3.180 0.185 3.255 0.445 ;
        RECT  3.165 0.705 3.255 1.030 ;
        RECT  3.045 0.545 3.245 0.615 ;
        RECT  2.955 0.355 3.045 0.795 ;
        RECT  2.845 0.355 2.955 0.455 ;
        RECT  2.860 0.695 2.955 0.795 ;
        RECT  2.740 0.695 2.860 1.065 ;
        RECT  2.675 0.545 2.850 0.615 ;
        RECT  2.760 0.195 2.845 0.455 ;
        RECT  2.605 0.205 2.675 0.615 ;
        RECT  2.160 0.205 2.605 0.275 ;
        RECT  2.300 0.350 2.410 0.420 ;
        RECT  2.300 0.985 2.410 1.065 ;
        RECT  2.230 0.350 2.300 1.065 ;
        RECT  2.090 0.205 2.160 1.045 ;
        RECT  1.940 0.320 2.010 1.045 ;
        RECT  1.900 0.320 1.940 0.480 ;
        RECT  1.515 0.975 1.940 1.045 ;
        RECT  1.830 0.570 1.870 0.690 ;
        RECT  1.760 0.200 1.830 0.905 ;
        RECT  1.690 0.200 1.760 0.270 ;
        RECT  1.660 0.835 1.760 0.905 ;
        RECT  1.425 0.845 1.515 1.045 ;
        RECT  1.160 0.845 1.425 0.915 ;
        RECT  1.300 0.705 1.410 0.775 ;
        RECT  1.300 0.195 1.395 0.275 ;
        RECT  1.150 0.985 1.320 1.075 ;
        RECT  1.230 0.195 1.300 0.775 ;
        RECT  1.080 0.325 1.160 0.915 ;
        RECT  0.930 0.985 1.150 1.055 ;
        RECT  1.030 0.835 1.080 0.915 ;
        RECT  0.900 0.325 0.980 0.770 ;
        RECT  0.860 0.850 0.930 1.055 ;
        RECT  0.515 0.700 0.900 0.770 ;
        RECT  0.125 0.850 0.860 0.920 ;
        RECT  0.515 0.340 0.545 0.470 ;
        RECT  0.445 0.340 0.515 0.770 ;
        RECT  0.105 0.195 0.125 0.335 ;
        RECT  0.105 0.850 0.125 1.030 ;
        RECT  0.035 0.195 0.105 1.030 ;
    END
END MUX3ND4BWP40

MACRO MUX4D0BWP40
    CLASS CORE ;
    FOREIGN MUX4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.195 3.465 1.045 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.355 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.480 1.365 0.800 ;
        RECT  1.205 0.480 1.275 0.670 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.015400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.495 0.945 0.800 ;
        RECT  0.800 0.495 0.865 0.650 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.485 2.205 0.775 ;
        RECT  2.095 0.485 2.135 0.655 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.015600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.480 1.505 0.800 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.115 3.500 0.115 ;
        RECT  3.180 -0.115 3.260 0.280 ;
        RECT  2.300 -0.115 3.180 0.115 ;
        RECT  2.180 -0.115 2.300 0.125 ;
        RECT  1.355 -0.115 2.180 0.115 ;
        RECT  1.265 -0.115 1.355 0.260 ;
        RECT  1.050 -0.115 1.265 0.115 ;
        RECT  0.980 -0.115 1.050 0.235 ;
        RECT  0.140 -0.115 0.980 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.145 3.500 1.375 ;
        RECT  3.180 0.930 3.260 1.375 ;
        RECT  2.300 1.145 3.180 1.375 ;
        RECT  2.180 1.135 2.300 1.375 ;
        RECT  1.380 1.145 2.180 1.375 ;
        RECT  1.260 1.050 1.380 1.375 ;
        RECT  0.980 1.145 1.260 1.375 ;
        RECT  0.860 1.050 0.980 1.375 ;
        RECT  0.130 1.145 0.860 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.220 0.370 3.290 0.810 ;
        RECT  3.040 0.370 3.220 0.440 ;
        RECT  3.080 0.740 3.220 0.810 ;
        RECT  2.880 0.530 3.150 0.650 ;
        RECT  3.000 0.740 3.080 1.065 ;
        RECT  2.970 0.195 3.040 0.440 ;
        RECT  1.850 0.195 2.970 0.265 ;
        RECT  2.810 0.345 2.880 0.980 ;
        RECT  2.630 0.345 2.700 1.065 ;
        RECT  2.580 0.345 2.630 0.420 ;
        RECT  2.600 0.785 2.630 1.065 ;
        RECT  1.540 0.995 2.600 1.065 ;
        RECT  2.500 0.555 2.560 0.675 ;
        RECT  2.430 0.350 2.500 0.915 ;
        RECT  2.025 0.335 2.100 0.405 ;
        RECT  2.025 0.855 2.090 0.925 ;
        RECT  1.955 0.335 2.025 0.925 ;
        RECT  1.780 0.195 1.850 0.925 ;
        RECT  1.495 0.195 1.710 0.270 ;
        RECT  1.575 0.360 1.645 0.800 ;
        RECT  1.470 0.910 1.540 1.065 ;
        RECT  1.425 0.195 1.495 0.400 ;
        RECT  0.510 0.910 1.470 0.980 ;
        RECT  1.125 0.330 1.425 0.400 ;
        RECT  1.055 0.330 1.125 0.830 ;
        RECT  0.900 0.330 1.055 0.400 ;
        RECT  0.820 0.195 0.900 0.400 ;
        RECT  0.550 0.195 0.820 0.265 ;
        RECT  0.660 0.355 0.730 0.840 ;
        RECT  0.510 0.380 0.570 0.460 ;
        RECT  0.430 0.380 0.510 0.980 ;
        RECT  0.270 0.215 0.340 0.990 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.220 0.910 0.270 0.990 ;
    END
END MUX4D0BWP40

MACRO MUX4D1BWP40
    CLASS CORE ;
    FOREIGN MUX4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.375 0.195 3.465 1.045 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.355 2.355 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.480 1.365 0.800 ;
        RECT  1.205 0.480 1.275 0.670 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.017600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.495 0.945 0.800 ;
        RECT  0.800 0.495 0.865 0.650 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.485 2.205 0.775 ;
        RECT  2.095 0.485 2.135 0.655 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.480 1.505 0.800 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.115 3.500 0.115 ;
        RECT  3.180 -0.115 3.260 0.290 ;
        RECT  2.300 -0.115 3.180 0.115 ;
        RECT  2.180 -0.115 2.300 0.125 ;
        RECT  1.355 -0.115 2.180 0.115 ;
        RECT  1.265 -0.115 1.355 0.260 ;
        RECT  1.050 -0.115 1.265 0.115 ;
        RECT  0.980 -0.115 1.050 0.235 ;
        RECT  0.140 -0.115 0.980 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.145 3.500 1.375 ;
        RECT  3.180 0.890 3.260 1.375 ;
        RECT  2.300 1.145 3.180 1.375 ;
        RECT  2.180 1.135 2.300 1.375 ;
        RECT  1.380 1.145 2.180 1.375 ;
        RECT  1.260 1.050 1.380 1.375 ;
        RECT  0.980 1.145 1.260 1.375 ;
        RECT  0.860 1.050 0.980 1.375 ;
        RECT  0.130 1.145 0.860 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.220 0.370 3.290 0.810 ;
        RECT  3.040 0.370 3.220 0.440 ;
        RECT  3.080 0.740 3.220 0.810 ;
        RECT  2.880 0.530 3.150 0.650 ;
        RECT  3.000 0.740 3.080 1.065 ;
        RECT  2.970 0.195 3.040 0.440 ;
        RECT  1.850 0.195 2.970 0.265 ;
        RECT  2.810 0.345 2.880 0.980 ;
        RECT  2.630 0.345 2.700 1.065 ;
        RECT  2.580 0.345 2.630 0.420 ;
        RECT  2.600 0.785 2.630 1.065 ;
        RECT  1.540 0.995 2.600 1.065 ;
        RECT  2.500 0.555 2.560 0.675 ;
        RECT  2.430 0.350 2.500 0.915 ;
        RECT  2.025 0.335 2.100 0.405 ;
        RECT  2.025 0.855 2.090 0.925 ;
        RECT  1.955 0.335 2.025 0.925 ;
        RECT  1.780 0.195 1.850 0.925 ;
        RECT  1.495 0.195 1.710 0.270 ;
        RECT  1.575 0.360 1.645 0.800 ;
        RECT  1.470 0.910 1.540 1.065 ;
        RECT  1.425 0.195 1.495 0.400 ;
        RECT  0.510 0.910 1.470 0.980 ;
        RECT  1.125 0.330 1.425 0.400 ;
        RECT  1.055 0.330 1.125 0.830 ;
        RECT  0.900 0.330 1.055 0.400 ;
        RECT  0.820 0.195 0.900 0.400 ;
        RECT  0.550 0.195 0.820 0.265 ;
        RECT  0.660 0.355 0.730 0.840 ;
        RECT  0.510 0.380 0.570 0.460 ;
        RECT  0.430 0.380 0.510 0.980 ;
        RECT  0.270 0.215 0.340 0.990 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.220 0.910 0.270 0.990 ;
    END
END MUX4D1BWP40

MACRO MUX4D2BWP40
    CLASS CORE ;
    FOREIGN MUX4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.136000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 0.195 4.165 1.045 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.355 3.060 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.047600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.525 0.480 1.645 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.640 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 0.495 1.085 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 0.485 2.905 0.775 ;
        RECT  2.770 0.485 2.810 0.655 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.355 2.100 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.405 -0.115 4.480 0.115 ;
        RECT  4.335 -0.115 4.405 0.510 ;
        RECT  3.960 -0.115 4.335 0.115 ;
        RECT  3.880 -0.115 3.960 0.290 ;
        RECT  2.975 -0.115 3.880 0.115 ;
        RECT  2.855 -0.115 2.975 0.125 ;
        RECT  1.705 -0.115 2.855 0.115 ;
        RECT  1.585 -0.115 1.705 0.210 ;
        RECT  1.045 -0.115 1.585 0.115 ;
        RECT  0.935 -0.115 1.045 0.210 ;
        RECT  0.140 -0.115 0.935 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.410 1.145 4.480 1.375 ;
        RECT  4.340 0.720 4.410 1.375 ;
        RECT  3.960 1.145 4.340 1.375 ;
        RECT  3.880 0.890 3.960 1.375 ;
        RECT  2.975 1.145 3.880 1.375 ;
        RECT  2.855 1.135 2.975 1.375 ;
        RECT  1.700 1.145 2.855 1.375 ;
        RECT  1.580 1.050 1.700 1.375 ;
        RECT  0.985 1.145 1.580 1.375 ;
        RECT  0.845 1.050 0.985 1.375 ;
        RECT  0.130 1.145 0.845 1.375 ;
        RECT  0.050 0.870 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.920 0.370 3.990 0.810 ;
        RECT  3.740 0.370 3.920 0.440 ;
        RECT  3.780 0.740 3.920 0.810 ;
        RECT  3.580 0.530 3.850 0.650 ;
        RECT  3.700 0.740 3.780 1.065 ;
        RECT  3.670 0.195 3.740 0.440 ;
        RECT  2.525 0.195 3.670 0.265 ;
        RECT  3.510 0.345 3.580 0.980 ;
        RECT  3.330 0.345 3.400 1.065 ;
        RECT  3.280 0.345 3.330 0.420 ;
        RECT  3.300 0.785 3.330 1.065 ;
        RECT  2.215 0.995 3.300 1.065 ;
        RECT  3.200 0.555 3.260 0.675 ;
        RECT  3.130 0.350 3.200 0.915 ;
        RECT  2.700 0.335 2.775 0.405 ;
        RECT  2.700 0.840 2.765 0.910 ;
        RECT  2.630 0.335 2.700 0.910 ;
        RECT  2.455 0.195 2.525 0.925 ;
        RECT  1.895 0.195 2.385 0.270 ;
        RECT  2.275 0.360 2.345 0.830 ;
        RECT  2.225 0.360 2.275 0.430 ;
        RECT  1.890 0.760 2.275 0.830 ;
        RECT  2.145 0.910 2.215 1.065 ;
        RECT  0.510 0.910 2.145 0.980 ;
        RECT  1.825 0.195 1.895 0.350 ;
        RECT  1.815 0.420 1.890 0.830 ;
        RECT  1.445 0.280 1.825 0.350 ;
        RECT  1.770 0.420 1.815 0.500 ;
        RECT  1.375 0.280 1.445 0.830 ;
        RECT  0.865 0.280 1.375 0.350 ;
        RECT  1.225 0.420 1.270 0.505 ;
        RECT  1.155 0.420 1.225 0.840 ;
        RECT  0.730 0.770 1.155 0.840 ;
        RECT  0.795 0.195 0.865 0.350 ;
        RECT  0.550 0.195 0.795 0.265 ;
        RECT  0.660 0.395 0.730 0.840 ;
        RECT  0.510 0.380 0.570 0.460 ;
        RECT  0.430 0.380 0.510 0.980 ;
        RECT  0.270 0.215 0.340 0.990 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.220 0.910 0.270 0.990 ;
    END
END MUX4D2BWP40

MACRO MUX4D4BWP40
    CLASS CORE ;
    FOREIGN MUX4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.195 5.300 0.475 ;
        RECT  5.215 0.735 5.300 1.045 ;
        RECT  5.005 0.380 5.215 0.820 ;
        RECT  4.930 0.380 5.005 0.475 ;
        RECT  4.930 0.735 5.005 0.820 ;
        RECT  4.840 0.195 4.930 0.475 ;
        RECT  4.840 0.735 4.930 1.045 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.495 3.760 0.765 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.047600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.885 0.480 2.065 0.800 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.495 0.385 0.645 ;
        RECT  0.170 0.495 0.250 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.054000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.495 1.275 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.057800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.205 0.485 3.340 0.765 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.044800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.360 0.355 2.485 0.625 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.540 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.540 0.485 ;
        RECT  5.100 -0.115 5.470 0.115 ;
        RECT  5.030 -0.115 5.100 0.280 ;
        RECT  4.725 -0.115 5.030 0.115 ;
        RECT  4.645 -0.115 4.725 0.290 ;
        RECT  3.745 -0.115 4.645 0.115 ;
        RECT  3.600 -0.115 3.745 0.125 ;
        RECT  3.345 -0.115 3.600 0.115 ;
        RECT  3.190 -0.115 3.345 0.125 ;
        RECT  2.065 -0.115 3.190 0.115 ;
        RECT  1.945 -0.115 2.065 0.200 ;
        RECT  1.675 -0.115 1.945 0.115 ;
        RECT  1.550 -0.115 1.675 0.200 ;
        RECT  1.240 -0.115 1.550 0.115 ;
        RECT  1.120 -0.115 1.240 0.200 ;
        RECT  0.345 -0.115 1.120 0.115 ;
        RECT  0.215 -0.115 0.345 0.215 ;
        RECT  0.000 -0.115 0.215 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.540 1.145 5.600 1.375 ;
        RECT  5.470 0.720 5.540 1.375 ;
        RECT  5.100 1.145 5.470 1.375 ;
        RECT  5.030 0.905 5.100 1.375 ;
        RECT  4.725 1.145 5.030 1.375 ;
        RECT  4.645 0.890 4.725 1.375 ;
        RECT  3.745 1.145 4.645 1.375 ;
        RECT  3.610 1.135 3.745 1.375 ;
        RECT  3.330 1.145 3.610 1.375 ;
        RECT  3.200 1.135 3.330 1.375 ;
        RECT  2.460 1.145 3.200 1.375 ;
        RECT  2.330 1.050 2.460 1.375 ;
        RECT  2.055 1.145 2.330 1.375 ;
        RECT  1.935 1.050 2.055 1.375 ;
        RECT  1.615 1.145 1.935 1.375 ;
        RECT  1.460 1.050 1.615 1.375 ;
        RECT  1.175 1.145 1.460 1.375 ;
        RECT  1.035 1.050 1.175 1.375 ;
        RECT  0.345 1.145 1.035 1.375 ;
        RECT  0.215 1.045 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.195 5.300 0.475 ;
        RECT  5.285 0.735 5.300 1.045 ;
        RECT  4.930 0.380 4.935 0.475 ;
        RECT  4.930 0.735 4.935 0.820 ;
        RECT  4.840 0.195 4.930 0.475 ;
        RECT  4.840 0.735 4.930 1.045 ;
        RECT  4.685 0.370 4.755 0.810 ;
        RECT  4.505 0.370 4.685 0.440 ;
        RECT  4.545 0.740 4.685 0.810 ;
        RECT  4.345 0.530 4.615 0.650 ;
        RECT  4.465 0.740 4.545 1.065 ;
        RECT  4.435 0.195 4.505 0.440 ;
        RECT  2.885 0.195 4.435 0.265 ;
        RECT  4.275 0.345 4.345 0.980 ;
        RECT  4.095 0.345 4.165 1.065 ;
        RECT  4.045 0.345 4.095 0.420 ;
        RECT  4.065 0.785 4.095 1.065 ;
        RECT  2.725 0.995 4.065 1.065 ;
        RECT  3.965 0.555 4.025 0.675 ;
        RECT  3.895 0.350 3.965 0.915 ;
        RECT  3.440 0.335 3.530 0.465 ;
        RECT  3.060 0.840 3.530 0.910 ;
        RECT  3.060 0.335 3.440 0.405 ;
        RECT  2.990 0.335 3.060 0.910 ;
        RECT  2.815 0.195 2.885 0.925 ;
        RECT  2.255 0.195 2.745 0.270 ;
        RECT  2.655 0.910 2.725 1.065 ;
        RECT  2.635 0.360 2.705 0.830 ;
        RECT  0.700 0.910 2.655 0.980 ;
        RECT  2.585 0.360 2.635 0.430 ;
        RECT  2.265 0.760 2.635 0.830 ;
        RECT  2.175 0.420 2.265 0.830 ;
        RECT  2.185 0.195 2.255 0.340 ;
        RECT  1.805 0.270 2.185 0.340 ;
        RECT  2.135 0.420 2.175 0.500 ;
        RECT  1.735 0.270 1.805 0.830 ;
        RECT  1.050 0.270 1.735 0.340 ;
        RECT  1.415 0.420 1.460 0.505 ;
        RECT  1.345 0.420 1.415 0.840 ;
        RECT  0.920 0.770 1.345 0.840 ;
        RECT  0.980 0.195 1.050 0.340 ;
        RECT  0.740 0.195 0.980 0.265 ;
        RECT  0.850 0.395 0.920 0.840 ;
        RECT  0.700 0.380 0.760 0.460 ;
        RECT  0.620 0.380 0.700 0.980 ;
        RECT  0.460 0.195 0.530 0.975 ;
        RECT  0.455 0.195 0.460 0.355 ;
        RECT  0.035 0.905 0.460 0.975 ;
        RECT  0.035 0.285 0.455 0.355 ;
    END
END MUX4D4BWP40

MACRO MUX4ND0BWP40
    CLASS CORE ;
    FOREIGN MUX4ND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.064000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.790 0.195 3.885 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.655 0.665 ;
        RECT  2.555 0.495 2.625 0.770 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.830 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.945 0.765 ;
        RECT  0.730 0.545 0.870 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.355 2.095 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.445 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.625 -0.115 3.920 0.115 ;
        RECT  3.505 -0.115 3.625 0.125 ;
        RECT  2.635 -0.115 3.505 0.115 ;
        RECT  2.515 -0.115 2.635 0.125 ;
        RECT  2.225 -0.115 2.515 0.115 ;
        RECT  2.105 -0.115 2.225 0.275 ;
        RECT  1.285 -0.115 2.105 0.115 ;
        RECT  1.215 -0.115 1.285 0.260 ;
        RECT  1.015 -0.115 1.215 0.115 ;
        RECT  0.945 -0.115 1.015 0.235 ;
        RECT  0.140 -0.115 0.945 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.645 1.145 3.920 1.375 ;
        RECT  3.525 1.120 3.645 1.375 ;
        RECT  2.625 1.145 3.525 1.375 ;
        RECT  2.505 1.135 2.625 1.375 ;
        RECT  2.225 1.145 2.505 1.375 ;
        RECT  2.105 1.120 2.225 1.375 ;
        RECT  1.335 1.145 2.105 1.375 ;
        RECT  1.215 1.050 1.335 1.375 ;
        RECT  0.945 1.145 1.215 1.375 ;
        RECT  0.825 1.050 0.945 1.375 ;
        RECT  0.140 1.145 0.825 1.375 ;
        RECT  0.040 0.885 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.510 3.690 0.630 ;
        RECT  3.600 0.195 3.675 0.630 ;
        RECT  3.575 0.700 3.645 1.050 ;
        RECT  3.215 0.195 3.600 0.265 ;
        RECT  3.520 0.700 3.575 0.770 ;
        RECT  2.015 0.980 3.575 1.050 ;
        RECT  3.435 0.500 3.520 0.770 ;
        RECT  3.365 0.840 3.465 0.910 ;
        RECT  3.365 0.335 3.405 0.435 ;
        RECT  3.285 0.335 3.365 0.910 ;
        RECT  3.145 0.195 3.215 0.880 ;
        RECT  3.085 0.195 3.145 0.370 ;
        RECT  2.915 0.195 2.985 0.900 ;
        RECT  2.405 0.195 2.915 0.265 ;
        RECT  2.775 0.345 2.845 0.910 ;
        RECT  2.645 0.345 2.775 0.415 ;
        RECT  2.675 0.840 2.775 0.910 ;
        RECT  2.335 0.195 2.405 0.900 ;
        RECT  2.185 0.500 2.265 0.910 ;
        RECT  1.780 0.840 2.185 0.910 ;
        RECT  1.920 0.700 2.025 0.770 ;
        RECT  1.920 0.195 2.015 0.275 ;
        RECT  1.945 0.980 2.015 1.065 ;
        RECT  1.495 0.995 1.945 1.065 ;
        RECT  1.850 0.195 1.920 0.770 ;
        RECT  1.710 0.195 1.780 0.910 ;
        RECT  1.665 0.840 1.710 0.910 ;
        RECT  1.445 0.200 1.640 0.280 ;
        RECT  1.515 0.370 1.585 0.835 ;
        RECT  1.460 0.755 1.515 0.835 ;
        RECT  1.425 0.910 1.495 1.065 ;
        RECT  1.375 0.200 1.445 0.400 ;
        RECT  0.510 0.910 1.425 0.980 ;
        RECT  1.085 0.330 1.375 0.400 ;
        RECT  1.015 0.330 1.085 0.830 ;
        RECT  0.875 0.330 1.015 0.400 ;
        RECT  0.805 0.195 0.875 0.400 ;
        RECT  0.515 0.195 0.805 0.270 ;
        RECT  0.660 0.350 0.730 0.460 ;
        RECT  0.660 0.720 0.725 0.840 ;
        RECT  0.590 0.350 0.660 0.840 ;
        RECT  0.510 0.340 0.520 0.470 ;
        RECT  0.430 0.340 0.510 0.980 ;
        RECT  0.270 0.215 0.340 1.065 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.240 0.745 0.270 1.065 ;
    END
END MUX4ND0BWP40

MACRO MUX4ND1BWP40
    CLASS CORE ;
    FOREIGN MUX4ND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.120800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.790 0.195 3.885 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.655 0.665 ;
        RECT  2.555 0.495 2.625 0.770 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.830 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.017400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.945 0.765 ;
        RECT  0.730 0.545 0.870 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.355 2.095 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.445 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.625 -0.115 3.920 0.115 ;
        RECT  3.505 -0.115 3.625 0.125 ;
        RECT  2.635 -0.115 3.505 0.115 ;
        RECT  2.515 -0.115 2.635 0.125 ;
        RECT  2.225 -0.115 2.515 0.115 ;
        RECT  2.105 -0.115 2.225 0.275 ;
        RECT  1.285 -0.115 2.105 0.115 ;
        RECT  1.215 -0.115 1.285 0.260 ;
        RECT  1.015 -0.115 1.215 0.115 ;
        RECT  0.945 -0.115 1.015 0.235 ;
        RECT  0.140 -0.115 0.945 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.645 1.145 3.920 1.375 ;
        RECT  3.525 1.120 3.645 1.375 ;
        RECT  2.625 1.145 3.525 1.375 ;
        RECT  2.505 1.135 2.625 1.375 ;
        RECT  2.225 1.145 2.505 1.375 ;
        RECT  2.105 1.120 2.225 1.375 ;
        RECT  1.335 1.145 2.105 1.375 ;
        RECT  1.215 1.050 1.335 1.375 ;
        RECT  0.945 1.145 1.215 1.375 ;
        RECT  0.825 1.050 0.945 1.375 ;
        RECT  0.140 1.145 0.825 1.375 ;
        RECT  0.040 0.910 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.510 3.690 0.630 ;
        RECT  3.600 0.195 3.675 0.630 ;
        RECT  3.575 0.700 3.645 1.050 ;
        RECT  3.215 0.195 3.600 0.265 ;
        RECT  3.520 0.700 3.575 0.770 ;
        RECT  2.015 0.980 3.575 1.050 ;
        RECT  3.435 0.500 3.520 0.770 ;
        RECT  3.365 0.840 3.465 0.910 ;
        RECT  3.365 0.335 3.405 0.435 ;
        RECT  3.285 0.335 3.365 0.910 ;
        RECT  3.145 0.195 3.215 0.880 ;
        RECT  3.085 0.195 3.145 0.370 ;
        RECT  2.915 0.195 2.985 0.900 ;
        RECT  2.405 0.195 2.915 0.265 ;
        RECT  2.775 0.345 2.845 0.910 ;
        RECT  2.645 0.345 2.775 0.415 ;
        RECT  2.675 0.840 2.775 0.910 ;
        RECT  2.335 0.195 2.405 0.900 ;
        RECT  2.185 0.500 2.265 0.910 ;
        RECT  1.780 0.840 2.185 0.910 ;
        RECT  1.920 0.700 2.025 0.770 ;
        RECT  1.920 0.195 2.015 0.275 ;
        RECT  1.945 0.980 2.015 1.065 ;
        RECT  1.495 0.995 1.945 1.065 ;
        RECT  1.850 0.195 1.920 0.770 ;
        RECT  1.710 0.195 1.780 0.910 ;
        RECT  1.665 0.840 1.710 0.910 ;
        RECT  1.445 0.200 1.640 0.280 ;
        RECT  1.515 0.370 1.585 0.835 ;
        RECT  1.460 0.755 1.515 0.835 ;
        RECT  1.425 0.910 1.495 1.065 ;
        RECT  1.375 0.200 1.445 0.400 ;
        RECT  0.510 0.910 1.425 0.980 ;
        RECT  1.085 0.330 1.375 0.400 ;
        RECT  1.015 0.330 1.085 0.830 ;
        RECT  0.875 0.330 1.015 0.400 ;
        RECT  0.805 0.195 0.875 0.400 ;
        RECT  0.515 0.195 0.805 0.270 ;
        RECT  0.660 0.350 0.730 0.460 ;
        RECT  0.660 0.720 0.725 0.840 ;
        RECT  0.590 0.350 0.660 0.840 ;
        RECT  0.510 0.340 0.520 0.470 ;
        RECT  0.430 0.340 0.510 0.980 ;
        RECT  0.270 0.215 0.340 1.065 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.240 0.745 0.270 1.065 ;
    END
END MUX4ND1BWP40

MACRO MUX4ND2BWP40
    CLASS CORE ;
    FOREIGN MUX4ND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.113250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.830 0.495 3.885 0.765 ;
        RECT  3.815 0.195 3.830 0.765 ;
        RECT  3.760 0.195 3.815 1.045 ;
        RECT  3.745 0.195 3.760 0.465 ;
        RECT  3.745 0.710 3.760 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.655 0.665 ;
        RECT  2.555 0.495 2.625 0.770 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.480 1.225 0.830 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.017400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.870 0.495 0.945 0.765 ;
        RECT  0.730 0.545 0.870 0.640 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.355 2.095 0.630 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.018200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.445 0.640 ;
        RECT  1.295 0.495 1.365 0.770 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 -0.115 4.060 0.115 ;
        RECT  3.935 -0.115 4.005 0.435 ;
        RECT  3.625 -0.115 3.935 0.115 ;
        RECT  3.505 -0.115 3.625 0.125 ;
        RECT  2.635 -0.115 3.505 0.115 ;
        RECT  2.515 -0.115 2.635 0.125 ;
        RECT  2.225 -0.115 2.515 0.115 ;
        RECT  2.105 -0.115 2.225 0.275 ;
        RECT  1.285 -0.115 2.105 0.115 ;
        RECT  1.215 -0.115 1.285 0.260 ;
        RECT  1.015 -0.115 1.215 0.115 ;
        RECT  0.945 -0.115 1.015 0.235 ;
        RECT  0.140 -0.115 0.945 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.145 4.060 1.375 ;
        RECT  3.935 0.900 4.005 1.375 ;
        RECT  3.645 1.145 3.935 1.375 ;
        RECT  3.525 1.120 3.645 1.375 ;
        RECT  2.625 1.145 3.525 1.375 ;
        RECT  2.505 1.135 2.625 1.375 ;
        RECT  2.225 1.145 2.505 1.375 ;
        RECT  2.105 1.120 2.225 1.375 ;
        RECT  1.335 1.145 2.105 1.375 ;
        RECT  1.215 1.050 1.335 1.375 ;
        RECT  0.945 1.145 1.215 1.375 ;
        RECT  0.825 1.050 0.945 1.375 ;
        RECT  0.140 1.145 0.825 1.375 ;
        RECT  0.040 0.895 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.510 3.690 0.630 ;
        RECT  3.600 0.195 3.675 0.630 ;
        RECT  3.575 0.700 3.645 1.050 ;
        RECT  3.215 0.195 3.600 0.265 ;
        RECT  3.520 0.700 3.575 0.770 ;
        RECT  2.015 0.980 3.575 1.050 ;
        RECT  3.435 0.500 3.520 0.770 ;
        RECT  3.365 0.840 3.465 0.910 ;
        RECT  3.365 0.335 3.405 0.435 ;
        RECT  3.285 0.335 3.365 0.910 ;
        RECT  3.145 0.195 3.215 0.880 ;
        RECT  3.085 0.195 3.145 0.370 ;
        RECT  2.915 0.195 2.985 0.900 ;
        RECT  2.405 0.195 2.915 0.265 ;
        RECT  2.775 0.345 2.845 0.910 ;
        RECT  2.645 0.345 2.775 0.415 ;
        RECT  2.675 0.840 2.775 0.910 ;
        RECT  2.335 0.195 2.405 0.900 ;
        RECT  2.185 0.500 2.265 0.910 ;
        RECT  1.780 0.840 2.185 0.910 ;
        RECT  1.920 0.700 2.025 0.770 ;
        RECT  1.920 0.195 2.015 0.275 ;
        RECT  1.945 0.980 2.015 1.065 ;
        RECT  1.495 0.995 1.945 1.065 ;
        RECT  1.850 0.195 1.920 0.770 ;
        RECT  1.710 0.195 1.780 0.910 ;
        RECT  1.665 0.840 1.710 0.910 ;
        RECT  1.445 0.200 1.640 0.280 ;
        RECT  1.515 0.370 1.585 0.835 ;
        RECT  1.460 0.755 1.515 0.835 ;
        RECT  1.425 0.910 1.495 1.065 ;
        RECT  1.375 0.200 1.445 0.400 ;
        RECT  0.510 0.910 1.425 0.980 ;
        RECT  1.085 0.330 1.375 0.400 ;
        RECT  1.015 0.330 1.085 0.830 ;
        RECT  0.875 0.330 1.015 0.400 ;
        RECT  0.805 0.195 0.875 0.400 ;
        RECT  0.515 0.195 0.805 0.270 ;
        RECT  0.660 0.350 0.730 0.460 ;
        RECT  0.660 0.720 0.725 0.840 ;
        RECT  0.590 0.350 0.660 0.840 ;
        RECT  0.510 0.340 0.520 0.470 ;
        RECT  0.430 0.340 0.510 0.980 ;
        RECT  0.270 0.215 0.340 1.065 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.240 0.745 0.270 1.065 ;
    END
END MUX4ND2BWP40

MACRO MUX4ND4BWP40
    CLASS CORE ;
    FOREIGN MUX4ND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.226500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.525 0.195 5.595 0.465 ;
        RECT  5.525 0.710 5.595 1.030 ;
        RECT  5.495 0.385 5.525 0.465 ;
        RECT  5.495 0.710 5.525 0.795 ;
        RECT  5.285 0.385 5.495 0.795 ;
        RECT  5.230 0.385 5.285 0.465 ;
        RECT  5.215 0.710 5.285 0.795 ;
        RECT  5.145 0.195 5.230 0.465 ;
        RECT  5.145 0.710 5.215 1.045 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.500 0.495 3.605 0.770 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.480 1.645 0.830 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.190 0.650 ;
        RECT  0.035 0.355 0.105 0.765 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.035600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.495 1.085 0.625 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.810 0.625 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.031000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.355 2.160 0.640 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.805 -0.115 5.880 0.115 ;
        RECT  5.735 -0.115 5.805 0.470 ;
        RECT  5.405 -0.115 5.735 0.115 ;
        RECT  5.335 -0.115 5.405 0.290 ;
        RECT  5.025 -0.115 5.335 0.115 ;
        RECT  4.910 -0.115 5.025 0.125 ;
        RECT  4.575 -0.115 4.910 0.115 ;
        RECT  4.425 -0.115 4.575 0.125 ;
        RECT  3.580 -0.115 4.425 0.115 ;
        RECT  3.460 -0.115 3.580 0.125 ;
        RECT  3.345 -0.115 3.460 0.115 ;
        RECT  3.230 -0.115 3.345 0.125 ;
        RECT  2.940 -0.115 3.230 0.115 ;
        RECT  2.820 -0.115 2.940 0.275 ;
        RECT  1.675 -0.115 2.820 0.115 ;
        RECT  1.530 -0.115 1.675 0.190 ;
        RECT  1.010 -0.115 1.530 0.115 ;
        RECT  0.885 -0.115 1.010 0.190 ;
        RECT  0.140 -0.115 0.885 0.115 ;
        RECT  0.035 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.035 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.805 1.145 5.880 1.375 ;
        RECT  5.735 0.695 5.805 1.375 ;
        RECT  5.430 1.145 5.735 1.375 ;
        RECT  5.310 0.880 5.430 1.375 ;
        RECT  5.035 1.145 5.310 1.375 ;
        RECT  4.960 0.705 5.035 1.375 ;
        RECT  4.590 1.145 4.960 1.375 ;
        RECT  4.450 1.120 4.590 1.375 ;
        RECT  3.570 1.145 4.450 1.375 ;
        RECT  3.450 1.135 3.570 1.375 ;
        RECT  3.355 1.145 3.450 1.375 ;
        RECT  3.210 1.120 3.355 1.375 ;
        RECT  2.940 1.145 3.210 1.375 ;
        RECT  2.820 1.120 2.940 1.375 ;
        RECT  1.665 1.145 2.820 1.375 ;
        RECT  1.545 1.050 1.665 1.375 ;
        RECT  1.015 1.145 1.545 1.375 ;
        RECT  0.895 1.050 1.015 1.375 ;
        RECT  0.140 1.145 0.895 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.195 5.595 0.465 ;
        RECT  5.565 0.710 5.595 1.030 ;
        RECT  5.145 0.195 5.215 0.465 ;
        RECT  5.145 0.710 5.215 1.045 ;
        RECT  5.075 0.535 5.205 0.610 ;
        RECT  5.000 0.195 5.075 0.610 ;
        RECT  4.160 0.195 5.000 0.265 ;
        RECT  4.820 0.540 4.890 1.050 ;
        RECT  4.450 0.540 4.820 0.610 ;
        RECT  2.730 0.980 4.820 1.050 ;
        RECT  4.310 0.335 4.805 0.435 ;
        RECT  4.310 0.780 4.750 0.900 ;
        RECT  4.230 0.335 4.310 0.900 ;
        RECT  4.090 0.195 4.160 0.880 ;
        RECT  4.030 0.195 4.090 0.370 ;
        RECT  3.860 0.195 3.930 0.900 ;
        RECT  3.120 0.195 3.860 0.265 ;
        RECT  3.720 0.345 3.790 0.910 ;
        RECT  3.590 0.345 3.720 0.415 ;
        RECT  3.620 0.840 3.720 0.910 ;
        RECT  3.050 0.195 3.120 0.900 ;
        RECT  2.900 0.500 2.980 0.910 ;
        RECT  2.485 0.840 2.900 0.910 ;
        RECT  2.625 0.700 2.740 0.770 ;
        RECT  2.625 0.195 2.730 0.275 ;
        RECT  2.660 0.980 2.730 1.065 ;
        RECT  2.310 0.995 2.660 1.065 ;
        RECT  2.555 0.195 2.625 0.770 ;
        RECT  2.415 0.195 2.485 0.910 ;
        RECT  2.380 0.840 2.415 0.910 ;
        RECT  1.825 0.195 2.345 0.275 ;
        RECT  2.240 0.910 2.310 1.065 ;
        RECT  2.230 0.370 2.300 0.835 ;
        RECT  0.510 0.910 2.240 0.980 ;
        RECT  1.800 0.755 2.230 0.835 ;
        RECT  1.755 0.195 1.825 0.330 ;
        RECT  1.730 0.400 1.800 0.835 ;
        RECT  1.415 0.260 1.755 0.330 ;
        RECT  1.345 0.260 1.415 0.830 ;
        RECT  0.670 0.260 1.345 0.330 ;
        RECT  1.155 0.400 1.225 0.840 ;
        RECT  0.735 0.770 1.155 0.840 ;
        RECT  0.625 0.415 0.735 0.840 ;
        RECT  0.600 0.195 0.670 0.330 ;
        RECT  0.515 0.195 0.600 0.270 ;
        RECT  0.510 0.340 0.520 0.470 ;
        RECT  0.430 0.340 0.510 0.980 ;
        RECT  0.270 0.215 0.340 1.065 ;
        RECT  0.220 0.215 0.270 0.295 ;
        RECT  0.240 0.745 0.270 1.065 ;
    END
END MUX4ND4BWP40

MACRO ND2D0BWP40
    CLASS CORE ;
    FOREIGN ND2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.053875 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.195 0.525 0.915 ;
        RECT  0.435 0.195 0.455 0.320 ;
        RECT  0.315 0.845 0.455 0.915 ;
        RECT  0.245 0.845 0.315 1.050 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.560 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.145 0.560 1.375 ;
        RECT  0.410 0.985 0.520 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.955 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END ND2D0BWP40

MACRO ND2D12BWP40
    CLASS CORE ;
    FOREIGN ND2D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.110600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.445 0.755 4.515 1.045 ;
        RECT  4.420 0.755 4.445 0.915 ;
        RECT  4.340 0.345 4.420 0.915 ;
        RECT  4.230 0.345 4.340 0.415 ;
        RECT  4.140 0.845 4.340 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.740 0.845 4.060 0.915 ;
        RECT  3.660 0.845 3.740 1.075 ;
        RECT  3.480 0.845 3.660 0.915 ;
        RECT  3.480 0.345 3.570 0.415 ;
        RECT  3.410 0.345 3.480 0.915 ;
        RECT  3.355 0.755 3.410 0.915 ;
        RECT  3.285 0.755 3.355 1.045 ;
        RECT  2.975 0.755 3.285 0.915 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
        RECT  2.595 0.845 2.770 0.915 ;
        RECT  2.525 0.845 2.595 1.075 ;
        RECT  2.215 0.845 2.525 0.915 ;
        RECT  2.145 0.845 2.215 1.075 ;
        RECT  1.995 0.845 2.145 0.915 ;
        RECT  1.995 0.345 2.050 0.425 ;
        RECT  1.900 0.345 1.995 0.915 ;
        RECT  1.840 0.495 1.900 0.915 ;
        RECT  1.785 0.495 1.840 1.045 ;
        RECT  1.760 0.735 1.785 1.045 ;
        RECT  1.460 0.735 1.760 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  1.075 0.845 1.270 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.440 0.845 0.625 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.358400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 0.495 4.725 0.625 ;
        RECT  4.490 0.195 4.570 0.625 ;
        RECT  4.135 0.195 4.490 0.265 ;
        RECT  4.065 0.195 4.135 0.415 ;
        RECT  3.940 0.345 4.065 0.415 ;
        RECT  3.815 0.345 3.940 0.630 ;
        RECT  3.745 0.345 3.815 0.415 ;
        RECT  3.665 0.195 3.745 0.415 ;
        RECT  3.330 0.195 3.665 0.265 ;
        RECT  3.255 0.195 3.330 0.625 ;
        RECT  3.000 0.495 3.255 0.625 ;
        RECT  2.930 0.205 3.000 0.625 ;
        RECT  2.590 0.205 2.930 0.275 ;
        RECT  2.510 0.205 2.590 0.415 ;
        RECT  2.445 0.345 2.510 0.415 ;
        RECT  2.345 0.345 2.445 0.635 ;
        RECT  2.230 0.345 2.345 0.415 ;
        RECT  2.150 0.205 2.230 0.415 ;
        RECT  1.790 0.205 2.150 0.275 ;
        RECT  1.715 0.205 1.790 0.410 ;
        RECT  1.645 0.340 1.715 0.410 ;
        RECT  1.560 0.340 1.645 0.640 ;
        RECT  1.505 0.340 1.560 0.410 ;
        RECT  1.435 0.205 1.505 0.410 ;
        RECT  1.070 0.205 1.435 0.275 ;
        RECT  0.990 0.205 1.070 0.415 ;
        RECT  0.845 0.345 0.990 0.415 ;
        RECT  0.735 0.345 0.845 0.635 ;
        RECT  0.710 0.345 0.735 0.415 ;
        RECT  0.630 0.205 0.710 0.415 ;
        RECT  0.290 0.205 0.630 0.275 ;
        RECT  0.220 0.205 0.290 0.640 ;
        RECT  0.160 0.495 0.220 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.371200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.665 0.705 1.015 0.775 ;
        RECT  0.525 0.495 0.665 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 -0.115 4.760 0.115 ;
        RECT  4.640 -0.115 4.710 0.395 ;
        RECT  3.960 -0.115 4.640 0.115 ;
        RECT  3.840 -0.115 3.960 0.275 ;
        RECT  3.180 -0.115 3.840 0.115 ;
        RECT  3.080 -0.115 3.180 0.415 ;
        RECT  2.420 -0.115 3.080 0.115 ;
        RECT  2.320 -0.115 2.420 0.275 ;
        RECT  1.645 -0.115 2.320 0.115 ;
        RECT  1.575 -0.115 1.645 0.260 ;
        RECT  0.900 -0.115 1.575 0.115 ;
        RECT  0.800 -0.115 0.900 0.275 ;
        RECT  0.140 -0.115 0.800 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.720 1.145 4.760 1.375 ;
        RECT  4.620 0.710 4.720 1.375 ;
        RECT  4.350 1.145 4.620 1.375 ;
        RECT  4.230 0.985 4.350 1.375 ;
        RECT  3.960 1.145 4.230 1.375 ;
        RECT  3.840 0.985 3.960 1.375 ;
        RECT  3.570 1.145 3.840 1.375 ;
        RECT  3.450 1.000 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.985 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.985 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.985 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.985 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.025 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.985 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.720 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.755 4.515 1.045 ;
        RECT  4.420 0.755 4.445 0.915 ;
        RECT  4.340 0.345 4.420 0.915 ;
        RECT  4.230 0.345 4.340 0.415 ;
        RECT  4.140 0.845 4.340 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.740 0.845 4.060 0.915 ;
        RECT  3.660 0.845 3.740 1.075 ;
        RECT  1.460 0.735 1.715 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  1.075 0.845 1.270 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.440 0.845 0.625 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        RECT  4.195 0.495 4.220 0.640 ;
        RECT  4.105 0.495 4.195 0.775 ;
        RECT  3.740 0.705 4.105 0.775 ;
        RECT  3.665 0.495 3.740 0.775 ;
        RECT  3.550 0.495 3.665 0.615 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.495 2.595 0.775 ;
        RECT  2.215 0.705 2.525 0.775 ;
        RECT  2.145 0.495 2.215 0.775 ;
        RECT  2.070 0.495 2.145 0.640 ;
        RECT  2.595 0.845 2.770 0.915 ;
        RECT  2.525 0.845 2.595 1.075 ;
        RECT  2.215 0.845 2.525 0.915 ;
        RECT  2.145 0.845 2.215 1.075 ;
        RECT  2.065 0.845 2.145 0.915 ;
        RECT  3.480 0.845 3.660 0.915 ;
        RECT  3.480 0.345 3.570 0.415 ;
        RECT  3.410 0.345 3.480 0.915 ;
        RECT  3.355 0.755 3.410 0.915 ;
        RECT  3.285 0.755 3.355 1.045 ;
        RECT  2.975 0.755 3.285 0.915 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
    END
END ND2D12BWP40

MACRO ND2D16BWP40
    CLASS CORE ;
    FOREIGN ND2D16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.485600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.985 0.755 6.055 1.045 ;
        RECT  5.960 0.755 5.985 0.915 ;
        RECT  5.880 0.345 5.960 0.915 ;
        RECT  5.770 0.345 5.880 0.415 ;
        RECT  5.680 0.845 5.880 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.280 0.845 5.600 0.915 ;
        RECT  5.200 0.845 5.280 1.075 ;
        RECT  5.020 0.845 5.200 0.915 ;
        RECT  5.020 0.345 5.110 0.415 ;
        RECT  4.950 0.345 5.020 0.915 ;
        RECT  4.895 0.755 4.950 0.915 ;
        RECT  4.825 0.755 4.895 1.045 ;
        RECT  4.515 0.755 4.825 0.915 ;
        RECT  4.440 0.755 4.515 1.045 ;
        RECT  4.390 0.755 4.440 0.915 ;
        RECT  4.310 0.345 4.390 0.915 ;
        RECT  4.230 0.345 4.310 0.425 ;
        RECT  4.140 0.845 4.310 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.760 0.845 4.060 0.915 ;
        RECT  3.680 0.845 3.760 1.075 ;
        RECT  3.535 0.845 3.680 0.915 ;
        RECT  3.535 0.345 3.590 0.425 ;
        RECT  3.440 0.345 3.535 0.915 ;
        RECT  3.380 0.495 3.440 0.915 ;
        RECT  3.325 0.495 3.380 1.045 ;
        RECT  3.300 0.735 3.325 1.045 ;
        RECT  3.000 0.735 3.300 0.915 ;
        RECT  2.920 0.735 3.000 1.045 ;
        RECT  2.890 0.735 2.920 0.915 ;
        RECT  2.810 0.345 2.890 0.915 ;
        RECT  2.710 0.345 2.810 0.425 ;
        RECT  2.620 0.845 2.810 0.915 ;
        RECT  2.540 0.845 2.620 1.075 ;
        RECT  2.240 0.845 2.540 0.915 ;
        RECT  2.160 0.845 2.240 1.075 ;
        RECT  1.980 0.845 2.160 0.915 ;
        RECT  1.980 0.345 2.070 0.425 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.860 0.755 1.900 0.915 ;
        RECT  1.785 0.755 1.860 1.045 ;
        RECT  1.485 0.755 1.785 0.915 ;
        RECT  1.395 0.755 1.485 1.045 ;
        RECT  1.375 0.755 1.395 0.915 ;
        RECT  1.305 0.345 1.375 0.915 ;
        RECT  1.190 0.345 1.305 0.415 ;
        RECT  1.100 0.845 1.305 0.915 ;
        RECT  1.020 0.845 1.100 1.075 ;
        RECT  0.720 0.845 1.020 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.473600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 0.495 6.265 0.625 ;
        RECT  6.030 0.195 6.110 0.625 ;
        RECT  5.675 0.195 6.030 0.265 ;
        RECT  5.605 0.195 5.675 0.415 ;
        RECT  5.480 0.345 5.605 0.415 ;
        RECT  5.355 0.345 5.480 0.630 ;
        RECT  5.285 0.345 5.355 0.415 ;
        RECT  5.205 0.195 5.285 0.415 ;
        RECT  4.870 0.195 5.205 0.265 ;
        RECT  4.795 0.195 4.870 0.625 ;
        RECT  4.540 0.495 4.795 0.625 ;
        RECT  4.470 0.205 4.540 0.625 ;
        RECT  4.130 0.205 4.470 0.275 ;
        RECT  4.050 0.205 4.130 0.415 ;
        RECT  3.985 0.345 4.050 0.415 ;
        RECT  3.885 0.345 3.985 0.635 ;
        RECT  3.770 0.345 3.885 0.415 ;
        RECT  3.690 0.205 3.770 0.415 ;
        RECT  3.330 0.205 3.690 0.275 ;
        RECT  3.255 0.205 3.330 0.410 ;
        RECT  3.185 0.340 3.255 0.410 ;
        RECT  3.100 0.340 3.185 0.640 ;
        RECT  3.045 0.340 3.100 0.410 ;
        RECT  2.975 0.205 3.045 0.410 ;
        RECT  2.610 0.205 2.975 0.275 ;
        RECT  2.530 0.205 2.610 0.415 ;
        RECT  2.385 0.345 2.530 0.415 ;
        RECT  2.275 0.345 2.385 0.635 ;
        RECT  2.250 0.345 2.275 0.415 ;
        RECT  2.170 0.205 2.250 0.415 ;
        RECT  1.830 0.205 2.170 0.275 ;
        RECT  1.760 0.205 1.830 0.640 ;
        RECT  1.525 0.495 1.760 0.640 ;
        RECT  1.455 0.195 1.525 0.640 ;
        RECT  1.095 0.195 1.455 0.265 ;
        RECT  1.015 0.195 1.095 0.415 ;
        RECT  0.945 0.345 1.015 0.415 ;
        RECT  0.810 0.345 0.945 0.630 ;
        RECT  0.715 0.345 0.810 0.415 ;
        RECT  0.645 0.195 0.715 0.415 ;
        RECT  0.290 0.195 0.645 0.265 ;
        RECT  0.210 0.195 0.290 0.625 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.499200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.740 0.625 ;
        RECT  2.555 0.495 2.625 0.775 ;
        RECT  2.205 0.705 2.555 0.775 ;
        RECT  2.065 0.495 2.205 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 -0.115 6.300 0.115 ;
        RECT  6.180 -0.115 6.250 0.395 ;
        RECT  5.500 -0.115 6.180 0.115 ;
        RECT  5.380 -0.115 5.500 0.275 ;
        RECT  4.720 -0.115 5.380 0.115 ;
        RECT  4.620 -0.115 4.720 0.415 ;
        RECT  3.960 -0.115 4.620 0.115 ;
        RECT  3.860 -0.115 3.960 0.275 ;
        RECT  3.185 -0.115 3.860 0.115 ;
        RECT  3.115 -0.115 3.185 0.260 ;
        RECT  2.440 -0.115 3.115 0.115 ;
        RECT  2.340 -0.115 2.440 0.275 ;
        RECT  1.665 -0.115 2.340 0.115 ;
        RECT  1.595 -0.115 1.665 0.415 ;
        RECT  0.930 -0.115 1.595 0.115 ;
        RECT  0.810 -0.115 0.930 0.275 ;
        RECT  0.120 -0.115 0.810 0.115 ;
        RECT  0.050 -0.115 0.120 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.260 1.145 6.300 1.375 ;
        RECT  6.160 0.710 6.260 1.375 ;
        RECT  5.890 1.145 6.160 1.375 ;
        RECT  5.770 0.985 5.890 1.375 ;
        RECT  5.500 1.145 5.770 1.375 ;
        RECT  5.380 0.985 5.500 1.375 ;
        RECT  5.110 1.145 5.380 1.375 ;
        RECT  4.990 1.000 5.110 1.375 ;
        RECT  4.730 1.145 4.990 1.375 ;
        RECT  4.610 0.985 4.730 1.375 ;
        RECT  4.350 1.145 4.610 1.375 ;
        RECT  4.230 0.985 4.350 1.375 ;
        RECT  3.970 1.145 4.230 1.375 ;
        RECT  3.850 0.985 3.970 1.375 ;
        RECT  3.590 1.145 3.850 1.375 ;
        RECT  3.470 0.985 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.090 1.025 3.210 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 0.985 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.330 0.985 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 0.985 2.070 1.375 ;
        RECT  1.695 1.145 1.950 1.375 ;
        RECT  1.565 0.985 1.695 1.375 ;
        RECT  1.300 1.145 1.565 1.375 ;
        RECT  1.200 1.030 1.300 1.375 ;
        RECT  0.930 1.145 1.200 1.375 ;
        RECT  0.810 0.985 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.985 0.755 6.055 1.045 ;
        RECT  5.960 0.755 5.985 0.915 ;
        RECT  5.880 0.345 5.960 0.915 ;
        RECT  5.770 0.345 5.880 0.415 ;
        RECT  5.680 0.845 5.880 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.280 0.845 5.600 0.915 ;
        RECT  5.200 0.845 5.280 1.075 ;
        RECT  5.020 0.845 5.200 0.915 ;
        RECT  5.020 0.345 5.110 0.415 ;
        RECT  4.950 0.345 5.020 0.915 ;
        RECT  4.895 0.755 4.950 0.915 ;
        RECT  4.825 0.755 4.895 1.045 ;
        RECT  4.515 0.755 4.825 0.915 ;
        RECT  4.440 0.755 4.515 1.045 ;
        RECT  4.390 0.755 4.440 0.915 ;
        RECT  4.310 0.345 4.390 0.915 ;
        RECT  4.230 0.345 4.310 0.425 ;
        RECT  4.140 0.845 4.310 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.760 0.845 4.060 0.915 ;
        RECT  3.680 0.845 3.760 1.075 ;
        RECT  3.605 0.845 3.680 0.915 ;
        RECT  3.000 0.735 3.255 0.915 ;
        RECT  2.920 0.735 3.000 1.045 ;
        RECT  2.890 0.735 2.920 0.915 ;
        RECT  2.810 0.345 2.890 0.915 ;
        RECT  2.710 0.345 2.810 0.425 ;
        RECT  2.620 0.845 2.810 0.915 ;
        RECT  2.540 0.845 2.620 1.075 ;
        RECT  2.240 0.845 2.540 0.915 ;
        RECT  2.160 0.845 2.240 1.075 ;
        RECT  1.980 0.845 2.160 0.915 ;
        RECT  1.980 0.345 2.070 0.425 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.860 0.755 1.900 0.915 ;
        RECT  1.785 0.755 1.860 1.045 ;
        RECT  1.485 0.755 1.785 0.915 ;
        RECT  1.395 0.755 1.485 1.045 ;
        RECT  1.375 0.755 1.395 0.915 ;
        RECT  1.305 0.345 1.375 0.915 ;
        RECT  1.190 0.345 1.305 0.415 ;
        RECT  1.100 0.845 1.305 0.915 ;
        RECT  1.020 0.845 1.100 1.075 ;
        RECT  0.720 0.845 1.020 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  5.205 0.495 5.280 0.775 ;
        RECT  5.090 0.495 5.205 0.615 ;
        RECT  4.135 0.495 4.235 0.640 ;
        RECT  4.065 0.495 4.135 0.775 ;
        RECT  3.755 0.705 4.065 0.775 ;
        RECT  3.685 0.495 3.755 0.775 ;
        RECT  3.610 0.495 3.685 0.640 ;
        RECT  1.095 0.495 1.210 0.625 ;
        RECT  1.020 0.495 1.095 0.775 ;
        RECT  0.675 0.705 1.020 0.775 ;
        RECT  0.585 0.495 0.675 0.775 ;
        RECT  0.560 0.495 0.585 0.640 ;
        RECT  0.265 0.755 0.335 1.045 ;
        RECT  5.735 0.495 5.760 0.640 ;
        RECT  5.645 0.495 5.735 0.775 ;
        RECT  5.280 0.705 5.645 0.775 ;
    END
END ND2D16BWP40

MACRO ND2D1BWP40
    CLASS CORE ;
    FOREIGN ND2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.107750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.215 0.525 0.915 ;
        RECT  0.435 0.215 0.455 0.385 ;
        RECT  0.315 0.845 0.455 0.915 ;
        RECT  0.245 0.845 0.315 1.050 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.455 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.560 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.145 0.560 1.375 ;
        RECT  0.410 0.985 0.520 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.770 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END ND2D1BWP40

MACRO ND2D20BWP40
    CLASS CORE ;
    FOREIGN ND2D20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.860600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.520 0.735 7.600 1.045 ;
        RECT  7.495 0.735 7.520 0.945 ;
        RECT  7.425 0.345 7.495 0.945 ;
        RECT  7.310 0.345 7.425 0.415 ;
        RECT  7.220 0.845 7.425 0.945 ;
        RECT  7.140 0.845 7.220 1.075 ;
        RECT  6.820 0.845 7.140 0.915 ;
        RECT  6.740 0.845 6.820 1.075 ;
        RECT  6.540 0.845 6.740 0.915 ;
        RECT  6.540 0.345 6.650 0.415 ;
        RECT  6.460 0.345 6.540 0.915 ;
        RECT  6.435 0.755 6.460 0.915 ;
        RECT  6.365 0.755 6.435 1.045 ;
        RECT  6.055 0.755 6.365 0.915 ;
        RECT  5.985 0.755 6.055 1.045 ;
        RECT  5.960 0.755 5.985 0.915 ;
        RECT  5.880 0.345 5.960 0.915 ;
        RECT  5.770 0.345 5.880 0.415 ;
        RECT  5.680 0.845 5.880 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.280 0.845 5.600 0.915 ;
        RECT  5.200 0.845 5.280 1.075 ;
        RECT  5.020 0.845 5.200 0.915 ;
        RECT  5.020 0.345 5.110 0.415 ;
        RECT  4.950 0.345 5.020 0.915 ;
        RECT  4.895 0.755 4.950 0.915 ;
        RECT  4.825 0.755 4.895 1.045 ;
        RECT  4.515 0.755 4.825 0.915 ;
        RECT  4.440 0.755 4.515 1.045 ;
        RECT  4.390 0.755 4.440 0.915 ;
        RECT  4.310 0.345 4.390 0.915 ;
        RECT  4.230 0.345 4.310 0.425 ;
        RECT  4.140 0.845 4.310 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.760 0.845 4.060 0.915 ;
        RECT  3.680 0.845 3.760 1.075 ;
        RECT  3.535 0.845 3.680 0.915 ;
        RECT  3.535 0.345 3.590 0.425 ;
        RECT  3.440 0.345 3.535 0.915 ;
        RECT  3.380 0.495 3.440 0.915 ;
        RECT  3.325 0.495 3.380 1.045 ;
        RECT  3.300 0.735 3.325 1.045 ;
        RECT  3.000 0.735 3.300 0.915 ;
        RECT  2.920 0.735 3.000 1.045 ;
        RECT  2.890 0.735 2.920 0.915 ;
        RECT  2.810 0.345 2.890 0.915 ;
        RECT  2.710 0.345 2.810 0.425 ;
        RECT  2.620 0.845 2.810 0.915 ;
        RECT  2.540 0.845 2.620 1.075 ;
        RECT  2.240 0.845 2.540 0.915 ;
        RECT  2.160 0.845 2.240 1.075 ;
        RECT  1.980 0.845 2.160 0.915 ;
        RECT  1.980 0.345 2.070 0.425 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.860 0.755 1.900 0.915 ;
        RECT  1.785 0.755 1.860 1.045 ;
        RECT  1.485 0.755 1.785 0.915 ;
        RECT  1.395 0.755 1.485 1.045 ;
        RECT  1.375 0.755 1.395 0.915 ;
        RECT  1.305 0.345 1.375 0.915 ;
        RECT  1.190 0.345 1.305 0.415 ;
        RECT  1.100 0.845 1.305 0.915 ;
        RECT  1.020 0.845 1.100 1.075 ;
        RECT  0.720 0.845 1.020 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.588800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.645 0.495 7.705 0.640 ;
        RECT  7.575 0.195 7.645 0.640 ;
        RECT  7.215 0.195 7.575 0.265 ;
        RECT  7.145 0.195 7.215 0.415 ;
        RECT  7.050 0.345 7.145 0.415 ;
        RECT  6.895 0.345 7.050 0.630 ;
        RECT  6.825 0.345 6.895 0.415 ;
        RECT  6.745 0.195 6.825 0.415 ;
        RECT  6.390 0.195 6.745 0.265 ;
        RECT  6.320 0.195 6.390 0.625 ;
        RECT  6.110 0.495 6.320 0.625 ;
        RECT  6.030 0.195 6.110 0.625 ;
        RECT  5.675 0.195 6.030 0.265 ;
        RECT  5.605 0.195 5.675 0.415 ;
        RECT  5.480 0.345 5.605 0.415 ;
        RECT  5.355 0.345 5.480 0.630 ;
        RECT  5.285 0.345 5.355 0.415 ;
        RECT  5.205 0.195 5.285 0.415 ;
        RECT  4.870 0.195 5.205 0.265 ;
        RECT  4.795 0.195 4.870 0.625 ;
        RECT  4.540 0.495 4.795 0.625 ;
        RECT  4.470 0.205 4.540 0.625 ;
        RECT  4.130 0.205 4.470 0.275 ;
        RECT  4.050 0.205 4.130 0.415 ;
        RECT  3.985 0.345 4.050 0.415 ;
        RECT  3.885 0.345 3.985 0.635 ;
        RECT  3.770 0.345 3.885 0.415 ;
        RECT  3.690 0.205 3.770 0.415 ;
        RECT  3.330 0.205 3.690 0.275 ;
        RECT  3.255 0.205 3.330 0.410 ;
        RECT  3.185 0.340 3.255 0.410 ;
        RECT  3.100 0.340 3.185 0.640 ;
        RECT  3.045 0.340 3.100 0.410 ;
        RECT  2.975 0.205 3.045 0.410 ;
        RECT  2.610 0.205 2.975 0.275 ;
        RECT  2.530 0.205 2.610 0.415 ;
        RECT  2.385 0.345 2.530 0.415 ;
        RECT  2.275 0.345 2.385 0.635 ;
        RECT  2.250 0.345 2.275 0.415 ;
        RECT  2.170 0.205 2.250 0.415 ;
        RECT  1.830 0.205 2.170 0.275 ;
        RECT  1.760 0.205 1.830 0.640 ;
        RECT  1.525 0.495 1.760 0.640 ;
        RECT  1.455 0.195 1.525 0.640 ;
        RECT  1.095 0.195 1.455 0.265 ;
        RECT  1.015 0.195 1.095 0.415 ;
        RECT  0.945 0.345 1.015 0.415 ;
        RECT  0.810 0.345 0.945 0.630 ;
        RECT  0.715 0.345 0.810 0.415 ;
        RECT  0.645 0.195 0.715 0.415 ;
        RECT  0.290 0.195 0.645 0.265 ;
        RECT  0.210 0.195 0.290 0.625 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.627200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.235 0.640 ;
        RECT  4.065 0.495 4.165 0.775 ;
        RECT  3.755 0.705 4.065 0.775 ;
        RECT  3.675 0.495 3.755 0.775 ;
        RECT  3.610 0.495 3.675 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.785 -0.115 7.840 0.115 ;
        RECT  7.715 -0.115 7.785 0.300 ;
        RECT  7.050 -0.115 7.715 0.115 ;
        RECT  6.930 -0.115 7.050 0.275 ;
        RECT  6.250 -0.115 6.930 0.115 ;
        RECT  6.180 -0.115 6.250 0.405 ;
        RECT  5.500 -0.115 6.180 0.115 ;
        RECT  5.380 -0.115 5.500 0.275 ;
        RECT  4.720 -0.115 5.380 0.115 ;
        RECT  4.620 -0.115 4.720 0.415 ;
        RECT  3.960 -0.115 4.620 0.115 ;
        RECT  3.860 -0.115 3.960 0.275 ;
        RECT  3.185 -0.115 3.860 0.115 ;
        RECT  3.115 -0.115 3.185 0.260 ;
        RECT  2.440 -0.115 3.115 0.115 ;
        RECT  2.340 -0.115 2.440 0.275 ;
        RECT  1.665 -0.115 2.340 0.115 ;
        RECT  1.595 -0.115 1.665 0.415 ;
        RECT  0.930 -0.115 1.595 0.115 ;
        RECT  0.810 -0.115 0.930 0.275 ;
        RECT  0.120 -0.115 0.810 0.115 ;
        RECT  0.050 -0.115 0.120 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 1.145 7.840 1.375 ;
        RECT  7.700 0.730 7.800 1.375 ;
        RECT  7.420 1.145 7.700 1.375 ;
        RECT  7.320 1.030 7.420 1.375 ;
        RECT  7.030 1.145 7.320 1.375 ;
        RECT  6.910 0.985 7.030 1.375 ;
        RECT  6.650 1.145 6.910 1.375 ;
        RECT  6.530 0.985 6.650 1.375 ;
        RECT  6.260 1.145 6.530 1.375 ;
        RECT  6.160 0.985 6.260 1.375 ;
        RECT  5.890 1.145 6.160 1.375 ;
        RECT  5.770 0.985 5.890 1.375 ;
        RECT  5.500 1.145 5.770 1.375 ;
        RECT  5.380 0.985 5.500 1.375 ;
        RECT  5.110 1.145 5.380 1.375 ;
        RECT  4.990 1.000 5.110 1.375 ;
        RECT  4.730 1.145 4.990 1.375 ;
        RECT  4.610 0.985 4.730 1.375 ;
        RECT  4.350 1.145 4.610 1.375 ;
        RECT  4.230 0.985 4.350 1.375 ;
        RECT  3.970 1.145 4.230 1.375 ;
        RECT  3.850 0.985 3.970 1.375 ;
        RECT  3.590 1.145 3.850 1.375 ;
        RECT  3.470 0.985 3.590 1.375 ;
        RECT  3.210 1.145 3.470 1.375 ;
        RECT  3.090 1.025 3.210 1.375 ;
        RECT  2.830 1.145 3.090 1.375 ;
        RECT  2.710 0.985 2.830 1.375 ;
        RECT  2.450 1.145 2.710 1.375 ;
        RECT  2.330 0.985 2.450 1.375 ;
        RECT  2.070 1.145 2.330 1.375 ;
        RECT  1.950 0.985 2.070 1.375 ;
        RECT  1.695 1.145 1.950 1.375 ;
        RECT  1.565 0.985 1.695 1.375 ;
        RECT  1.300 1.145 1.565 1.375 ;
        RECT  1.200 1.030 1.300 1.375 ;
        RECT  0.930 1.145 1.200 1.375 ;
        RECT  0.810 0.985 0.930 1.375 ;
        RECT  0.550 1.145 0.810 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.520 0.735 7.600 1.045 ;
        RECT  7.495 0.735 7.520 0.945 ;
        RECT  7.425 0.345 7.495 0.945 ;
        RECT  7.310 0.345 7.425 0.415 ;
        RECT  7.220 0.845 7.425 0.945 ;
        RECT  7.140 0.845 7.220 1.075 ;
        RECT  6.820 0.845 7.140 0.915 ;
        RECT  6.740 0.845 6.820 1.075 ;
        RECT  6.540 0.845 6.740 0.915 ;
        RECT  6.540 0.345 6.650 0.415 ;
        RECT  6.460 0.345 6.540 0.915 ;
        RECT  6.435 0.755 6.460 0.915 ;
        RECT  6.365 0.755 6.435 1.045 ;
        RECT  6.055 0.755 6.365 0.915 ;
        RECT  5.985 0.755 6.055 1.045 ;
        RECT  5.960 0.755 5.985 0.915 ;
        RECT  5.880 0.345 5.960 0.915 ;
        RECT  5.770 0.345 5.880 0.415 ;
        RECT  5.680 0.845 5.880 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.280 0.845 5.600 0.915 ;
        RECT  5.200 0.845 5.280 1.075 ;
        RECT  5.020 0.845 5.200 0.915 ;
        RECT  5.020 0.345 5.110 0.415 ;
        RECT  4.950 0.345 5.020 0.915 ;
        RECT  4.895 0.755 4.950 0.915 ;
        RECT  4.825 0.755 4.895 1.045 ;
        RECT  4.515 0.755 4.825 0.915 ;
        RECT  4.440 0.755 4.515 1.045 ;
        RECT  4.390 0.755 4.440 0.915 ;
        RECT  4.310 0.345 4.390 0.915 ;
        RECT  4.230 0.345 4.310 0.425 ;
        RECT  4.140 0.845 4.310 0.915 ;
        RECT  4.060 0.845 4.140 1.075 ;
        RECT  3.760 0.845 4.060 0.915 ;
        RECT  3.680 0.845 3.760 1.075 ;
        RECT  3.605 0.845 3.680 0.915 ;
        RECT  3.000 0.735 3.255 0.915 ;
        RECT  2.920 0.735 3.000 1.045 ;
        RECT  2.890 0.735 2.920 0.915 ;
        RECT  2.810 0.345 2.890 0.915 ;
        RECT  2.710 0.345 2.810 0.425 ;
        RECT  2.620 0.845 2.810 0.915 ;
        RECT  2.540 0.845 2.620 1.075 ;
        RECT  2.240 0.845 2.540 0.915 ;
        RECT  2.160 0.845 2.240 1.075 ;
        RECT  1.980 0.845 2.160 0.915 ;
        RECT  1.980 0.345 2.070 0.425 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.860 0.755 1.900 0.915 ;
        RECT  1.785 0.755 1.860 1.045 ;
        RECT  1.485 0.755 1.785 0.915 ;
        RECT  1.395 0.755 1.485 1.045 ;
        RECT  1.375 0.755 1.395 0.915 ;
        RECT  1.305 0.345 1.375 0.915 ;
        RECT  1.190 0.345 1.305 0.415 ;
        RECT  1.100 0.845 1.305 0.915 ;
        RECT  1.020 0.845 1.100 1.075 ;
        RECT  0.720 0.845 1.020 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        RECT  7.215 0.495 7.330 0.625 ;
        RECT  7.140 0.495 7.215 0.775 ;
        RECT  6.775 0.705 7.140 0.775 ;
        RECT  6.685 0.495 6.775 0.775 ;
        RECT  6.660 0.495 6.685 0.640 ;
        RECT  5.735 0.495 5.760 0.640 ;
        RECT  5.645 0.495 5.735 0.775 ;
        RECT  5.280 0.705 5.645 0.775 ;
        RECT  5.205 0.495 5.280 0.775 ;
        RECT  5.090 0.495 5.205 0.615 ;
        RECT  2.575 0.495 2.740 0.625 ;
        RECT  2.505 0.495 2.575 0.775 ;
        RECT  2.205 0.705 2.505 0.775 ;
        RECT  2.065 0.495 2.205 0.775 ;
        RECT  1.095 0.495 1.210 0.625 ;
        RECT  1.020 0.495 1.095 0.775 ;
        RECT  0.675 0.705 1.020 0.775 ;
        RECT  0.585 0.495 0.675 0.775 ;
        RECT  0.560 0.495 0.585 0.640 ;
    END
END ND2D20BWP40

MACRO ND2D24BWP40
    CLASS CORE ;
    FOREIGN ND2D24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 2.235600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.055 0.735 9.140 1.045 ;
        RECT  9.035 0.735 9.055 0.945 ;
        RECT  8.965 0.345 9.035 0.945 ;
        RECT  8.850 0.345 8.965 0.415 ;
        RECT  8.760 0.845 8.965 0.945 ;
        RECT  8.680 0.845 8.760 1.075 ;
        RECT  8.360 0.845 8.680 0.915 ;
        RECT  8.280 0.845 8.360 1.075 ;
        RECT  8.090 0.845 8.280 0.915 ;
        RECT  8.090 0.345 8.200 0.415 ;
        RECT  8.010 0.345 8.090 0.915 ;
        RECT  7.975 0.755 8.010 0.915 ;
        RECT  7.905 0.755 7.975 1.045 ;
        RECT  7.595 0.755 7.905 0.915 ;
        RECT  7.525 0.755 7.595 1.045 ;
        RECT  7.500 0.755 7.525 0.915 ;
        RECT  7.420 0.345 7.500 0.915 ;
        RECT  7.310 0.345 7.420 0.415 ;
        RECT  7.220 0.845 7.420 0.915 ;
        RECT  7.140 0.845 7.220 1.075 ;
        RECT  6.820 0.845 7.140 0.915 ;
        RECT  6.740 0.845 6.820 1.075 ;
        RECT  6.560 0.845 6.740 0.915 ;
        RECT  6.560 0.345 6.650 0.415 ;
        RECT  6.490 0.345 6.560 0.915 ;
        RECT  6.435 0.755 6.490 0.915 ;
        RECT  6.365 0.755 6.435 1.045 ;
        RECT  6.055 0.755 6.365 0.915 ;
        RECT  5.980 0.755 6.055 1.045 ;
        RECT  5.930 0.755 5.980 0.915 ;
        RECT  5.850 0.345 5.930 0.915 ;
        RECT  5.770 0.345 5.850 0.425 ;
        RECT  5.680 0.845 5.850 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.300 0.845 5.600 0.915 ;
        RECT  5.220 0.845 5.300 1.075 ;
        RECT  5.075 0.845 5.220 0.915 ;
        RECT  5.075 0.345 5.130 0.425 ;
        RECT  4.980 0.345 5.075 0.915 ;
        RECT  4.920 0.495 4.980 0.915 ;
        RECT  4.865 0.495 4.920 1.045 ;
        RECT  4.840 0.735 4.865 1.045 ;
        RECT  4.540 0.735 4.840 0.915 ;
        RECT  4.460 0.735 4.540 1.045 ;
        RECT  4.430 0.735 4.460 0.915 ;
        RECT  4.350 0.345 4.430 0.915 ;
        RECT  4.250 0.345 4.350 0.425 ;
        RECT  4.160 0.845 4.350 0.915 ;
        RECT  4.080 0.845 4.160 1.075 ;
        RECT  3.780 0.845 4.080 0.915 ;
        RECT  3.700 0.845 3.780 1.075 ;
        RECT  3.520 0.845 3.700 0.915 ;
        RECT  3.520 0.345 3.610 0.425 ;
        RECT  3.440 0.345 3.520 0.915 ;
        RECT  3.400 0.755 3.440 0.915 ;
        RECT  3.325 0.755 3.400 1.045 ;
        RECT  3.025 0.755 3.325 0.915 ;
        RECT  2.935 0.755 3.025 1.045 ;
        RECT  2.915 0.755 2.935 0.915 ;
        RECT  2.845 0.345 2.915 0.915 ;
        RECT  2.730 0.345 2.845 0.415 ;
        RECT  2.640 0.845 2.845 0.915 ;
        RECT  2.560 0.845 2.640 1.075 ;
        RECT  2.260 0.845 2.560 0.915 ;
        RECT  2.180 0.845 2.260 1.075 ;
        RECT  1.980 0.845 2.180 0.915 ;
        RECT  1.980 0.345 2.090 0.415 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.875 0.755 1.900 0.915 ;
        RECT  1.805 0.755 1.875 1.045 ;
        RECT  1.495 0.755 1.805 0.915 ;
        RECT  1.425 0.755 1.495 1.045 ;
        RECT  1.395 0.755 1.425 0.915 ;
        RECT  1.325 0.345 1.395 0.915 ;
        RECT  1.210 0.345 1.325 0.415 ;
        RECT  1.120 0.845 1.325 0.915 ;
        RECT  1.040 0.845 1.120 1.075 ;
        RECT  0.720 0.845 1.040 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.704000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.185 0.495 9.245 0.640 ;
        RECT  9.115 0.195 9.185 0.640 ;
        RECT  8.755 0.195 9.115 0.265 ;
        RECT  8.685 0.195 8.755 0.415 ;
        RECT  8.590 0.345 8.685 0.415 ;
        RECT  8.435 0.345 8.590 0.630 ;
        RECT  8.365 0.345 8.435 0.415 ;
        RECT  8.285 0.195 8.365 0.415 ;
        RECT  7.940 0.195 8.285 0.265 ;
        RECT  7.860 0.195 7.940 0.625 ;
        RECT  7.650 0.495 7.860 0.625 ;
        RECT  7.570 0.195 7.650 0.625 ;
        RECT  7.215 0.195 7.570 0.265 ;
        RECT  7.145 0.195 7.215 0.415 ;
        RECT  7.020 0.345 7.145 0.415 ;
        RECT  6.895 0.345 7.020 0.630 ;
        RECT  6.825 0.345 6.895 0.415 ;
        RECT  6.745 0.195 6.825 0.415 ;
        RECT  6.410 0.195 6.745 0.265 ;
        RECT  6.335 0.195 6.410 0.625 ;
        RECT  6.080 0.495 6.335 0.625 ;
        RECT  6.010 0.205 6.080 0.625 ;
        RECT  5.670 0.205 6.010 0.275 ;
        RECT  5.590 0.205 5.670 0.415 ;
        RECT  5.525 0.345 5.590 0.415 ;
        RECT  5.425 0.345 5.525 0.635 ;
        RECT  5.310 0.345 5.425 0.415 ;
        RECT  5.230 0.205 5.310 0.415 ;
        RECT  4.870 0.205 5.230 0.275 ;
        RECT  4.795 0.205 4.870 0.410 ;
        RECT  4.725 0.340 4.795 0.410 ;
        RECT  4.640 0.340 4.725 0.640 ;
        RECT  4.585 0.340 4.640 0.410 ;
        RECT  4.515 0.205 4.585 0.410 ;
        RECT  4.150 0.205 4.515 0.275 ;
        RECT  4.070 0.205 4.150 0.415 ;
        RECT  3.925 0.345 4.070 0.415 ;
        RECT  3.815 0.345 3.925 0.635 ;
        RECT  3.790 0.345 3.815 0.415 ;
        RECT  3.710 0.205 3.790 0.415 ;
        RECT  3.370 0.205 3.710 0.275 ;
        RECT  3.300 0.205 3.370 0.640 ;
        RECT  3.065 0.495 3.300 0.640 ;
        RECT  2.995 0.195 3.065 0.640 ;
        RECT  2.635 0.195 2.995 0.265 ;
        RECT  2.555 0.195 2.635 0.415 ;
        RECT  2.485 0.345 2.555 0.415 ;
        RECT  2.350 0.345 2.485 0.630 ;
        RECT  2.255 0.345 2.350 0.415 ;
        RECT  2.185 0.195 2.255 0.415 ;
        RECT  1.830 0.195 2.185 0.265 ;
        RECT  1.760 0.195 1.830 0.640 ;
        RECT  1.545 0.495 1.760 0.640 ;
        RECT  1.475 0.195 1.545 0.640 ;
        RECT  1.115 0.195 1.475 0.265 ;
        RECT  1.015 0.195 1.115 0.415 ;
        RECT  0.945 0.345 1.015 0.415 ;
        RECT  0.825 0.345 0.945 0.630 ;
        RECT  0.715 0.345 0.825 0.415 ;
        RECT  0.645 0.195 0.715 0.415 ;
        RECT  0.290 0.195 0.645 0.265 ;
        RECT  0.210 0.195 0.290 0.625 ;
        RECT  0.095 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.755200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.705 0.495 5.775 0.640 ;
        RECT  5.605 0.495 5.705 0.775 ;
        RECT  5.295 0.705 5.605 0.775 ;
        RECT  5.215 0.495 5.295 0.775 ;
        RECT  5.150 0.495 5.215 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.325 -0.115 9.380 0.115 ;
        RECT  9.255 -0.115 9.325 0.300 ;
        RECT  8.590 -0.115 9.255 0.115 ;
        RECT  8.470 -0.115 8.590 0.275 ;
        RECT  7.790 -0.115 8.470 0.115 ;
        RECT  7.720 -0.115 7.790 0.400 ;
        RECT  7.040 -0.115 7.720 0.115 ;
        RECT  6.920 -0.115 7.040 0.275 ;
        RECT  6.260 -0.115 6.920 0.115 ;
        RECT  6.160 -0.115 6.260 0.415 ;
        RECT  5.500 -0.115 6.160 0.115 ;
        RECT  5.400 -0.115 5.500 0.275 ;
        RECT  4.725 -0.115 5.400 0.115 ;
        RECT  4.655 -0.115 4.725 0.260 ;
        RECT  3.980 -0.115 4.655 0.115 ;
        RECT  3.880 -0.115 3.980 0.275 ;
        RECT  3.205 -0.115 3.880 0.115 ;
        RECT  3.135 -0.115 3.205 0.415 ;
        RECT  2.470 -0.115 3.135 0.115 ;
        RECT  2.350 -0.115 2.470 0.275 ;
        RECT  1.690 -0.115 2.350 0.115 ;
        RECT  1.620 -0.115 1.690 0.415 ;
        RECT  0.940 -0.115 1.620 0.115 ;
        RECT  0.820 -0.115 0.940 0.275 ;
        RECT  0.120 -0.115 0.820 0.115 ;
        RECT  0.050 -0.115 0.120 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.340 1.145 9.380 1.375 ;
        RECT  9.240 0.730 9.340 1.375 ;
        RECT  8.960 1.145 9.240 1.375 ;
        RECT  8.860 1.030 8.960 1.375 ;
        RECT  8.570 1.145 8.860 1.375 ;
        RECT  8.450 0.985 8.570 1.375 ;
        RECT  8.190 1.145 8.450 1.375 ;
        RECT  8.070 0.985 8.190 1.375 ;
        RECT  7.800 1.145 8.070 1.375 ;
        RECT  7.700 0.985 7.800 1.375 ;
        RECT  7.430 1.145 7.700 1.375 ;
        RECT  7.310 0.985 7.430 1.375 ;
        RECT  7.040 1.145 7.310 1.375 ;
        RECT  6.920 0.985 7.040 1.375 ;
        RECT  6.650 1.145 6.920 1.375 ;
        RECT  6.530 1.000 6.650 1.375 ;
        RECT  6.270 1.145 6.530 1.375 ;
        RECT  6.150 0.985 6.270 1.375 ;
        RECT  5.890 1.145 6.150 1.375 ;
        RECT  5.770 0.985 5.890 1.375 ;
        RECT  5.510 1.145 5.770 1.375 ;
        RECT  5.390 0.985 5.510 1.375 ;
        RECT  5.130 1.145 5.390 1.375 ;
        RECT  5.010 0.985 5.130 1.375 ;
        RECT  4.750 1.145 5.010 1.375 ;
        RECT  4.630 1.025 4.750 1.375 ;
        RECT  4.370 1.145 4.630 1.375 ;
        RECT  4.250 0.985 4.370 1.375 ;
        RECT  3.990 1.145 4.250 1.375 ;
        RECT  3.870 0.985 3.990 1.375 ;
        RECT  3.610 1.145 3.870 1.375 ;
        RECT  3.490 0.985 3.610 1.375 ;
        RECT  3.230 1.145 3.490 1.375 ;
        RECT  3.105 0.985 3.230 1.375 ;
        RECT  2.840 1.145 3.105 1.375 ;
        RECT  2.740 1.030 2.840 1.375 ;
        RECT  2.470 1.145 2.740 1.375 ;
        RECT  2.350 0.985 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 0.985 2.090 1.375 ;
        RECT  1.710 1.145 1.970 1.375 ;
        RECT  1.590 0.985 1.710 1.375 ;
        RECT  1.320 1.145 1.590 1.375 ;
        RECT  1.220 1.030 1.320 1.375 ;
        RECT  0.940 1.145 1.220 1.375 ;
        RECT  0.820 0.985 0.940 1.375 ;
        RECT  0.550 1.145 0.820 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.055 0.735 9.140 1.045 ;
        RECT  9.035 0.735 9.055 0.945 ;
        RECT  8.965 0.345 9.035 0.945 ;
        RECT  8.850 0.345 8.965 0.415 ;
        RECT  8.760 0.845 8.965 0.945 ;
        RECT  8.680 0.845 8.760 1.075 ;
        RECT  8.360 0.845 8.680 0.915 ;
        RECT  8.280 0.845 8.360 1.075 ;
        RECT  8.090 0.845 8.280 0.915 ;
        RECT  8.090 0.345 8.200 0.415 ;
        RECT  8.010 0.345 8.090 0.915 ;
        RECT  7.975 0.755 8.010 0.915 ;
        RECT  7.905 0.755 7.975 1.045 ;
        RECT  7.595 0.755 7.905 0.915 ;
        RECT  7.525 0.755 7.595 1.045 ;
        RECT  7.500 0.755 7.525 0.915 ;
        RECT  7.420 0.345 7.500 0.915 ;
        RECT  7.310 0.345 7.420 0.415 ;
        RECT  7.220 0.845 7.420 0.915 ;
        RECT  2.730 0.345 2.845 0.415 ;
        RECT  2.640 0.845 2.845 0.915 ;
        RECT  2.560 0.845 2.640 1.075 ;
        RECT  2.260 0.845 2.560 0.915 ;
        RECT  2.180 0.845 2.260 1.075 ;
        RECT  1.980 0.845 2.180 0.915 ;
        RECT  1.980 0.345 2.090 0.415 ;
        RECT  1.900 0.345 1.980 0.915 ;
        RECT  1.875 0.755 1.900 0.915 ;
        RECT  1.805 0.755 1.875 1.045 ;
        RECT  1.495 0.755 1.805 0.915 ;
        RECT  1.425 0.755 1.495 1.045 ;
        RECT  1.395 0.755 1.425 0.915 ;
        RECT  1.325 0.345 1.395 0.915 ;
        RECT  1.210 0.345 1.325 0.415 ;
        RECT  1.120 0.845 1.325 0.915 ;
        RECT  1.040 0.845 1.120 1.075 ;
        RECT  0.720 0.845 1.040 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        RECT  8.755 0.495 8.870 0.625 ;
        RECT  8.680 0.495 8.755 0.775 ;
        RECT  8.315 0.705 8.680 0.775 ;
        RECT  8.225 0.495 8.315 0.775 ;
        RECT  8.200 0.495 8.225 0.640 ;
        RECT  7.275 0.495 7.300 0.640 ;
        RECT  7.185 0.495 7.275 0.775 ;
        RECT  6.820 0.705 7.185 0.775 ;
        RECT  6.745 0.495 6.820 0.775 ;
        RECT  6.630 0.495 6.745 0.615 ;
        RECT  4.115 0.495 4.280 0.625 ;
        RECT  4.045 0.495 4.115 0.775 ;
        RECT  3.745 0.705 4.045 0.775 ;
        RECT  3.605 0.495 3.745 0.775 ;
        RECT  2.635 0.495 2.750 0.625 ;
        RECT  2.560 0.495 2.635 0.775 ;
        RECT  2.215 0.705 2.560 0.775 ;
        RECT  2.125 0.495 2.215 0.775 ;
        RECT  2.100 0.495 2.125 0.640 ;
        RECT  1.115 0.495 1.230 0.625 ;
        RECT  1.040 0.495 1.115 0.775 ;
        RECT  0.675 0.705 1.040 0.775 ;
        RECT  0.585 0.495 0.675 0.775 ;
        RECT  0.560 0.495 0.585 0.640 ;
        RECT  7.140 0.845 7.220 1.075 ;
        RECT  6.820 0.845 7.140 0.915 ;
        RECT  6.740 0.845 6.820 1.075 ;
        RECT  6.560 0.845 6.740 0.915 ;
        RECT  6.560 0.345 6.650 0.415 ;
        RECT  6.490 0.345 6.560 0.915 ;
        RECT  6.435 0.755 6.490 0.915 ;
        RECT  6.365 0.755 6.435 1.045 ;
        RECT  6.055 0.755 6.365 0.915 ;
        RECT  5.980 0.755 6.055 1.045 ;
        RECT  5.930 0.755 5.980 0.915 ;
        RECT  5.850 0.345 5.930 0.915 ;
        RECT  5.770 0.345 5.850 0.425 ;
        RECT  5.680 0.845 5.850 0.915 ;
        RECT  5.600 0.845 5.680 1.075 ;
        RECT  5.300 0.845 5.600 0.915 ;
        RECT  5.220 0.845 5.300 1.075 ;
        RECT  5.145 0.845 5.220 0.915 ;
        RECT  4.540 0.735 4.795 0.915 ;
        RECT  4.460 0.735 4.540 1.045 ;
        RECT  4.430 0.735 4.460 0.915 ;
        RECT  4.350 0.345 4.430 0.915 ;
        RECT  4.250 0.345 4.350 0.425 ;
        RECT  4.160 0.845 4.350 0.915 ;
        RECT  4.080 0.845 4.160 1.075 ;
        RECT  3.780 0.845 4.080 0.915 ;
        RECT  3.700 0.845 3.780 1.075 ;
        RECT  3.520 0.845 3.700 0.915 ;
        RECT  3.520 0.345 3.610 0.425 ;
        RECT  3.440 0.345 3.520 0.915 ;
        RECT  3.400 0.755 3.440 0.915 ;
        RECT  3.325 0.755 3.400 1.045 ;
        RECT  3.025 0.755 3.325 0.915 ;
        RECT  2.935 0.755 3.025 1.045 ;
        RECT  2.915 0.755 2.935 0.915 ;
        RECT  2.845 0.345 2.915 0.915 ;
    END
END ND2D24BWP40

MACRO ND2D2BWP40
    CLASS CORE ;
    FOREIGN ND2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.187500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.835 0.720 1.035 ;
        RECT  0.390 0.835 0.640 0.915 ;
        RECT  0.355 0.345 0.390 0.915 ;
        RECT  0.315 0.345 0.355 1.045 ;
        RECT  0.240 0.345 0.315 0.415 ;
        RECT  0.260 0.705 0.315 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.675 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.355 0.105 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.980 0.115 ;
        RECT  0.630 -0.115 0.730 0.275 ;
        RECT  0.000 -0.115 0.630 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.705 0.910 1.375 ;
        RECT  0.540 1.145 0.830 1.375 ;
        RECT  0.440 0.990 0.540 1.375 ;
        RECT  0.145 1.145 0.440 1.375 ;
        RECT  0.075 0.705 0.145 1.375 ;
        RECT  0.000 1.145 0.075 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.835 0.185 0.925 0.415 ;
        RECT  0.530 0.345 0.835 0.415 ;
        RECT  0.460 0.205 0.530 0.415 ;
        RECT  0.035 0.205 0.460 0.275 ;
    END
END ND2D2BWP40

MACRO ND2D3BWP40
    CLASS CORE ;
    FOREIGN ND2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.313250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.835 1.155 1.075 ;
        RECT  0.705 0.835 1.040 0.905 ;
        RECT  0.635 0.835 0.705 1.065 ;
        RECT  0.525 0.835 0.635 0.905 ;
        RECT  0.455 0.350 0.525 0.905 ;
        RECT  0.130 0.350 0.455 0.420 ;
        RECT  0.330 0.835 0.455 0.905 ;
        RECT  0.230 0.835 0.330 1.075 ;
        RECT  0.050 0.215 0.130 0.420 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.495 1.110 0.625 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.385 0.640 ;
        RECT  0.145 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.415 ;
        RECT  0.920 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.920 0.275 ;
        RECT  0.000 -0.115 0.820 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.700 1.360 1.375 ;
        RECT  0.920 1.145 1.260 1.375 ;
        RECT  0.820 0.990 0.920 1.375 ;
        RECT  0.520 1.145 0.820 1.375 ;
        RECT  0.420 0.990 0.520 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.840 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.030 0.185 1.130 0.425 ;
        RECT  0.695 0.355 1.030 0.425 ;
        RECT  0.625 0.210 0.695 0.425 ;
        RECT  0.220 0.210 0.625 0.280 ;
    END
END ND2D3BWP40

MACRO ND2D4BWP40
    CLASS CORE ;
    FOREIGN ND2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.375000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.735 1.575 1.045 ;
        RECT  1.430 0.345 1.435 1.045 ;
        RECT  1.365 0.345 1.430 0.945 ;
        RECT  1.250 0.345 1.365 0.415 ;
        RECT  1.160 0.845 1.365 0.945 ;
        RECT  1.080 0.845 1.160 1.075 ;
        RECT  0.720 0.845 1.080 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.585 0.495 1.645 0.640 ;
        RECT  1.515 0.195 1.585 0.640 ;
        RECT  1.155 0.195 1.515 0.265 ;
        RECT  1.085 0.195 1.155 0.415 ;
        RECT  0.950 0.345 1.085 0.415 ;
        RECT  0.850 0.345 0.950 0.630 ;
        RECT  0.715 0.345 0.850 0.415 ;
        RECT  0.645 0.195 0.715 0.415 ;
        RECT  0.290 0.195 0.645 0.265 ;
        RECT  0.210 0.195 0.290 0.625 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.270 0.625 ;
        RECT  1.080 0.495 1.155 0.775 ;
        RECT  0.675 0.705 1.080 0.775 ;
        RECT  0.585 0.495 0.675 0.775 ;
        RECT  0.560 0.495 0.585 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 -0.115 1.820 0.115 ;
        RECT  1.680 -0.115 1.780 0.415 ;
        RECT  0.960 -0.115 1.680 0.115 ;
        RECT  0.840 -0.115 0.960 0.275 ;
        RECT  0.120 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.120 0.385 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.145 1.820 1.375 ;
        RECT  1.680 0.730 1.780 1.375 ;
        RECT  1.360 1.145 1.680 1.375 ;
        RECT  1.260 1.030 1.360 1.375 ;
        RECT  0.960 1.145 1.260 1.375 ;
        RECT  0.840 0.985 0.960 1.375 ;
        RECT  0.550 1.145 0.840 1.375 ;
        RECT  0.430 0.985 0.550 1.375 ;
        RECT  0.140 1.145 0.430 1.375 ;
        RECT  0.040 0.710 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.250 0.345 1.295 0.415 ;
        RECT  1.160 0.845 1.295 0.945 ;
        RECT  1.080 0.845 1.160 1.075 ;
        RECT  0.720 0.845 1.080 0.915 ;
        RECT  0.640 0.845 0.720 1.075 ;
        RECT  0.440 0.845 0.640 0.915 ;
        RECT  0.440 0.345 0.550 0.415 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.335 0.755 0.360 0.915 ;
        RECT  0.265 0.755 0.335 1.045 ;
    END
END ND2D4BWP40

MACRO ND2D6BWP40
    CLASS CORE ;
    FOREIGN ND2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.640500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.195 2.625 0.420 ;
        RECT  2.510 0.195 2.555 0.905 ;
        RECT  2.375 0.350 2.510 0.905 ;
        RECT  2.345 0.350 2.375 1.065 ;
        RECT  2.090 0.350 2.345 0.420 ;
        RECT  2.305 0.835 2.345 1.065 ;
        RECT  1.985 0.835 2.305 0.905 ;
        RECT  1.915 0.835 1.985 1.065 ;
        RECT  1.575 0.835 1.915 0.905 ;
        RECT  1.505 0.835 1.575 1.065 ;
        RECT  1.115 0.835 1.505 0.905 ;
        RECT  1.045 0.835 1.115 1.065 ;
        RECT  0.705 0.835 1.045 0.905 ;
        RECT  0.635 0.835 0.705 1.065 ;
        RECT  0.315 0.835 0.635 0.905 ;
        RECT  0.130 0.350 0.530 0.420 ;
        RECT  0.245 0.835 0.315 1.065 ;
        RECT  0.130 0.835 0.245 0.905 ;
        RECT  0.050 0.215 0.130 0.905 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.885 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.075 0.495 2.205 0.765 ;
        RECT  0.665 0.695 2.075 0.765 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.320 0.495 0.595 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 -0.115 2.660 0.115 ;
        RECT  1.700 -0.115 1.800 0.275 ;
        RECT  1.360 -0.115 1.700 0.115 ;
        RECT  1.260 -0.115 1.360 0.275 ;
        RECT  0.920 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.920 0.275 ;
        RECT  0.000 -0.115 0.820 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.145 2.660 1.375 ;
        RECT  2.520 0.990 2.620 1.375 ;
        RECT  2.200 1.145 2.520 1.375 ;
        RECT  2.100 0.990 2.200 1.375 ;
        RECT  1.800 1.145 2.100 1.375 ;
        RECT  1.700 0.990 1.800 1.375 ;
        RECT  1.360 1.145 1.700 1.375 ;
        RECT  1.260 0.990 1.360 1.375 ;
        RECT  0.920 1.145 1.260 1.375 ;
        RECT  0.820 0.990 0.920 1.375 ;
        RECT  0.520 1.145 0.820 1.375 ;
        RECT  0.420 0.990 0.520 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.990 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.090 0.350 2.275 0.420 ;
        RECT  1.985 0.835 2.275 0.905 ;
        RECT  1.915 0.835 1.985 1.065 ;
        RECT  1.575 0.835 1.915 0.905 ;
        RECT  1.505 0.835 1.575 1.065 ;
        RECT  1.115 0.835 1.505 0.905 ;
        RECT  1.045 0.835 1.115 1.065 ;
        RECT  0.705 0.835 1.045 0.905 ;
        RECT  0.635 0.835 0.705 1.065 ;
        RECT  0.315 0.835 0.635 0.905 ;
        RECT  0.130 0.350 0.530 0.420 ;
        RECT  0.245 0.835 0.315 1.065 ;
        RECT  0.130 0.835 0.245 0.905 ;
        RECT  0.050 0.215 0.130 0.905 ;
        RECT  1.995 0.210 2.400 0.280 ;
        RECT  1.925 0.210 1.995 0.425 ;
        RECT  1.575 0.355 1.925 0.425 ;
        RECT  1.505 0.195 1.575 0.425 ;
        RECT  1.115 0.355 1.505 0.425 ;
        RECT  1.045 0.195 1.115 0.425 ;
        RECT  0.695 0.355 1.045 0.425 ;
        RECT  0.625 0.210 0.695 0.425 ;
        RECT  0.220 0.210 0.625 0.280 ;
    END
END ND2D6BWP40

MACRO ND2D8BWP40
    CLASS CORE ;
    FOREIGN ND2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.735600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
        RECT  2.595 0.845 2.770 0.915 ;
        RECT  2.525 0.845 2.595 1.075 ;
        RECT  2.215 0.845 2.525 0.915 ;
        RECT  2.145 0.845 2.215 1.075 ;
        RECT  1.995 0.845 2.145 0.915 ;
        RECT  1.995 0.345 2.050 0.425 ;
        RECT  1.900 0.345 1.995 0.915 ;
        RECT  1.840 0.495 1.900 0.915 ;
        RECT  1.785 0.495 1.840 1.045 ;
        RECT  1.760 0.735 1.785 1.045 ;
        RECT  1.460 0.735 1.760 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  1.075 0.845 1.270 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.440 0.845 0.625 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.000 0.495 3.130 0.625 ;
        RECT  2.930 0.205 3.000 0.625 ;
        RECT  2.590 0.205 2.930 0.275 ;
        RECT  2.510 0.205 2.590 0.415 ;
        RECT  2.445 0.345 2.510 0.415 ;
        RECT  2.345 0.345 2.445 0.635 ;
        RECT  2.230 0.345 2.345 0.415 ;
        RECT  2.150 0.205 2.230 0.415 ;
        RECT  1.790 0.205 2.150 0.275 ;
        RECT  1.715 0.205 1.790 0.410 ;
        RECT  1.645 0.340 1.715 0.410 ;
        RECT  1.560 0.340 1.645 0.640 ;
        RECT  1.505 0.340 1.560 0.410 ;
        RECT  1.435 0.205 1.505 0.410 ;
        RECT  1.070 0.205 1.435 0.275 ;
        RECT  0.990 0.205 1.070 0.415 ;
        RECT  0.845 0.345 0.990 0.415 ;
        RECT  0.735 0.345 0.845 0.635 ;
        RECT  0.710 0.345 0.735 0.415 ;
        RECT  0.630 0.205 0.710 0.415 ;
        RECT  0.290 0.205 0.630 0.275 ;
        RECT  0.220 0.205 0.290 0.640 ;
        RECT  0.160 0.495 0.220 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.495 1.085 0.775 ;
        RECT  0.665 0.705 1.015 0.775 ;
        RECT  0.525 0.495 0.665 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 -0.115 3.220 0.115 ;
        RECT  3.080 -0.115 3.180 0.415 ;
        RECT  2.420 -0.115 3.080 0.115 ;
        RECT  2.320 -0.115 2.420 0.275 ;
        RECT  1.645 -0.115 2.320 0.115 ;
        RECT  1.575 -0.115 1.645 0.260 ;
        RECT  0.900 -0.115 1.575 0.115 ;
        RECT  0.800 -0.115 0.900 0.275 ;
        RECT  0.140 -0.115 0.800 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.145 3.220 1.375 ;
        RECT  3.090 0.720 3.170 1.375 ;
        RECT  2.810 1.145 3.090 1.375 ;
        RECT  2.690 0.985 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.985 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.985 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 1.025 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.985 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.985 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.720 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.900 0.755 2.975 1.045 ;
        RECT  2.850 0.755 2.900 0.915 ;
        RECT  2.770 0.345 2.850 0.915 ;
        RECT  2.690 0.345 2.770 0.425 ;
        RECT  2.595 0.845 2.770 0.915 ;
        RECT  2.525 0.845 2.595 1.075 ;
        RECT  2.215 0.845 2.525 0.915 ;
        RECT  2.145 0.845 2.215 1.075 ;
        RECT  2.065 0.845 2.145 0.915 ;
        RECT  1.460 0.735 1.715 0.915 ;
        RECT  1.380 0.735 1.460 1.045 ;
        RECT  1.350 0.735 1.380 0.915 ;
        RECT  1.270 0.345 1.350 0.915 ;
        RECT  1.170 0.345 1.270 0.425 ;
        RECT  1.075 0.845 1.270 0.915 ;
        RECT  1.005 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.005 0.915 ;
        RECT  0.625 0.845 0.695 1.075 ;
        RECT  0.440 0.845 0.625 0.915 ;
        RECT  0.440 0.345 0.530 0.425 ;
        RECT  0.360 0.345 0.440 0.915 ;
        RECT  0.320 0.755 0.360 0.915 ;
        RECT  0.245 0.755 0.320 1.045 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.495 2.595 0.775 ;
        RECT  2.215 0.705 2.525 0.775 ;
        RECT  2.145 0.495 2.215 0.775 ;
        RECT  2.070 0.495 2.145 0.640 ;
    END
END ND2D8BWP40

MACRO ND3D0BWP40
    CLASS CORE ;
    FOREIGN ND3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.104250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.715 0.185 0.735 0.445 ;
        RECT  0.715 0.730 0.735 1.045 ;
        RECT  0.385 0.730 0.715 0.800 ;
        RECT  0.265 0.730 0.385 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.325 0.385 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.130 0.270 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.840 1.375 ;
        RECT  0.470 0.940 0.550 1.375 ;
        RECT  0.140 1.145 0.470 1.375 ;
        RECT  0.040 0.945 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND3D0BWP40

MACRO ND3D12BWP40
    CLASS CORE ;
    FOREIGN ND3D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.539000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.055 0.355 7.060 0.425 ;
        RECT  6.950 0.705 7.050 0.970 ;
        RECT  6.670 0.705 6.950 0.815 ;
        RECT  6.570 0.705 6.670 0.970 ;
        RECT  6.290 0.705 6.570 0.815 ;
        RECT  6.190 0.705 6.290 0.970 ;
        RECT  6.055 0.705 6.190 0.815 ;
        RECT  5.900 0.355 6.055 0.815 ;
        RECT  5.845 0.355 5.900 0.990 ;
        RECT  5.040 0.355 5.845 0.425 ;
        RECT  5.820 0.705 5.845 0.990 ;
        RECT  5.520 0.705 5.820 0.815 ;
        RECT  5.440 0.705 5.520 0.990 ;
        RECT  5.140 0.705 5.440 0.815 ;
        RECT  5.060 0.705 5.140 0.990 ;
        RECT  4.580 0.705 5.060 0.815 ;
        RECT  4.500 0.705 4.580 0.990 ;
        RECT  4.200 0.705 4.500 0.815 ;
        RECT  4.120 0.705 4.200 0.990 ;
        RECT  3.820 0.705 4.120 0.815 ;
        RECT  3.740 0.705 3.820 0.990 ;
        RECT  3.440 0.705 3.740 0.815 ;
        RECT  3.360 0.705 3.440 0.990 ;
        RECT  3.060 0.705 3.360 0.815 ;
        RECT  2.980 0.705 3.060 0.990 ;
        RECT  2.680 0.705 2.980 0.815 ;
        RECT  2.600 0.705 2.680 0.990 ;
        RECT  2.300 0.705 2.600 0.815 ;
        RECT  2.220 0.705 2.300 0.990 ;
        RECT  1.920 0.705 2.220 0.815 ;
        RECT  1.840 0.705 1.920 0.990 ;
        RECT  1.540 0.705 1.840 0.815 ;
        RECT  1.460 0.705 1.540 0.990 ;
        RECT  1.160 0.705 1.460 0.815 ;
        RECT  1.080 0.705 1.160 0.990 ;
        RECT  0.790 0.705 1.080 0.815 ;
        RECT  0.690 0.705 0.790 0.970 ;
        RECT  0.410 0.705 0.690 0.815 ;
        RECT  0.310 0.705 0.410 0.970 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 0.495 2.245 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.495 4.255 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.495 5.715 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.115 7.280 0.115 ;
        RECT  2.220 -0.115 2.300 0.285 ;
        RECT  1.920 -0.115 2.220 0.115 ;
        RECT  1.840 -0.115 1.920 0.285 ;
        RECT  1.540 -0.115 1.840 0.115 ;
        RECT  1.460 -0.115 1.540 0.285 ;
        RECT  1.160 -0.115 1.460 0.115 ;
        RECT  1.080 -0.115 1.160 0.285 ;
        RECT  0.780 -0.115 1.080 0.115 ;
        RECT  0.700 -0.115 0.780 0.285 ;
        RECT  0.400 -0.115 0.700 0.115 ;
        RECT  0.320 -0.115 0.400 0.285 ;
        RECT  0.000 -0.115 0.320 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.225 1.145 7.280 1.375 ;
        RECT  7.155 0.695 7.225 1.375 ;
        RECT  6.870 1.145 7.155 1.375 ;
        RECT  6.750 0.885 6.870 1.375 ;
        RECT  6.490 1.145 6.750 1.375 ;
        RECT  6.370 0.885 6.490 1.375 ;
        RECT  6.110 1.145 6.370 1.375 ;
        RECT  5.990 0.885 6.110 1.375 ;
        RECT  5.730 1.145 5.990 1.375 ;
        RECT  5.610 0.885 5.730 1.375 ;
        RECT  5.350 1.145 5.610 1.375 ;
        RECT  5.230 0.885 5.350 1.375 ;
        RECT  4.950 1.145 5.230 1.375 ;
        RECT  4.870 0.885 4.950 1.375 ;
        RECT  4.770 1.145 4.870 1.375 ;
        RECT  4.690 0.885 4.770 1.375 ;
        RECT  4.390 1.145 4.690 1.375 ;
        RECT  4.310 0.885 4.390 1.375 ;
        RECT  4.030 1.145 4.310 1.375 ;
        RECT  3.910 0.885 4.030 1.375 ;
        RECT  3.650 1.145 3.910 1.375 ;
        RECT  3.530 0.885 3.650 1.375 ;
        RECT  3.270 1.145 3.530 1.375 ;
        RECT  3.150 0.885 3.270 1.375 ;
        RECT  2.890 1.145 3.150 1.375 ;
        RECT  2.770 0.885 2.890 1.375 ;
        RECT  2.510 1.145 2.770 1.375 ;
        RECT  2.390 0.885 2.510 1.375 ;
        RECT  2.130 1.145 2.390 1.375 ;
        RECT  2.010 0.885 2.130 1.375 ;
        RECT  1.750 1.145 2.010 1.375 ;
        RECT  1.630 0.885 1.750 1.375 ;
        RECT  1.370 1.145 1.630 1.375 ;
        RECT  1.250 0.885 1.370 1.375 ;
        RECT  0.990 1.145 1.250 1.375 ;
        RECT  0.870 0.885 0.990 1.375 ;
        RECT  0.610 1.145 0.870 1.375 ;
        RECT  0.490 0.885 0.610 1.375 ;
        RECT  0.130 1.145 0.490 1.375 ;
        RECT  0.050 0.695 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.125 0.355 7.060 0.425 ;
        RECT  6.950 0.705 7.050 0.970 ;
        RECT  6.670 0.705 6.950 0.815 ;
        RECT  6.570 0.705 6.670 0.970 ;
        RECT  6.290 0.705 6.570 0.815 ;
        RECT  6.190 0.705 6.290 0.970 ;
        RECT  6.125 0.705 6.190 0.815 ;
        RECT  5.040 0.355 5.775 0.425 ;
        RECT  5.520 0.705 5.775 0.815 ;
        RECT  5.440 0.705 5.520 0.990 ;
        RECT  5.140 0.705 5.440 0.815 ;
        RECT  5.060 0.705 5.140 0.990 ;
        RECT  4.580 0.705 5.060 0.815 ;
        RECT  4.500 0.705 4.580 0.990 ;
        RECT  4.200 0.705 4.500 0.815 ;
        RECT  4.120 0.705 4.200 0.990 ;
        RECT  3.820 0.705 4.120 0.815 ;
        RECT  3.740 0.705 3.820 0.990 ;
        RECT  3.440 0.705 3.740 0.815 ;
        RECT  3.360 0.705 3.440 0.990 ;
        RECT  3.060 0.705 3.360 0.815 ;
        RECT  2.980 0.705 3.060 0.990 ;
        RECT  2.680 0.705 2.980 0.815 ;
        RECT  2.600 0.705 2.680 0.990 ;
        RECT  2.300 0.705 2.600 0.815 ;
        RECT  2.220 0.705 2.300 0.990 ;
        RECT  1.920 0.705 2.220 0.815 ;
        RECT  1.840 0.705 1.920 0.990 ;
        RECT  1.540 0.705 1.840 0.815 ;
        RECT  1.460 0.705 1.540 0.990 ;
        RECT  1.160 0.705 1.460 0.815 ;
        RECT  1.080 0.705 1.160 0.990 ;
        RECT  0.790 0.705 1.080 0.815 ;
        RECT  0.690 0.705 0.790 0.970 ;
        RECT  0.410 0.705 0.690 0.815 ;
        RECT  0.310 0.705 0.410 0.970 ;
        RECT  7.155 0.215 7.225 0.475 ;
        RECT  2.580 0.215 7.155 0.285 ;
        RECT  6.140 0.550 6.805 0.625 ;
        RECT  2.485 0.355 4.790 0.425 ;
        RECT  2.415 0.185 2.485 0.425 ;
        RECT  2.105 0.355 2.415 0.425 ;
        RECT  2.035 0.185 2.105 0.425 ;
        RECT  1.725 0.355 2.035 0.425 ;
        RECT  1.655 0.185 1.725 0.425 ;
        RECT  1.345 0.355 1.655 0.425 ;
        RECT  1.275 0.185 1.345 0.425 ;
        RECT  0.965 0.355 1.275 0.425 ;
        RECT  0.895 0.185 0.965 0.425 ;
        RECT  0.585 0.355 0.895 0.425 ;
        RECT  0.515 0.185 0.585 0.425 ;
        RECT  0.140 0.355 0.515 0.425 ;
        RECT  0.040 0.185 0.140 0.425 ;
    END
END ND3D12BWP40

MACRO ND3D1BWP40
    CLASS CORE ;
    FOREIGN ND3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.208500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.045 ;
        RECT  0.715 0.185 0.735 0.445 ;
        RECT  0.715 0.730 0.735 1.045 ;
        RECT  0.385 0.730 0.715 0.800 ;
        RECT  0.265 0.730 0.385 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.325 0.385 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.130 -0.115 0.840 0.115 ;
        RECT  0.050 -0.115 0.130 0.410 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.145 0.840 1.375 ;
        RECT  0.470 0.870 0.550 1.375 ;
        RECT  0.140 1.145 0.470 1.375 ;
        RECT  0.040 0.775 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND3D1BWP40

MACRO ND3D2BWP40
    CLASS CORE ;
    FOREIGN ND3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.322500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.290 1.365 1.045 ;
        RECT  1.135 0.290 1.280 0.360 ;
        RECT  0.930 0.835 1.280 0.905 ;
        RECT  1.055 0.195 1.135 0.360 ;
        RECT  0.595 0.195 1.055 0.265 ;
        RECT  0.850 0.835 0.930 1.070 ;
        RECT  0.550 0.835 0.850 0.905 ;
        RECT  0.470 0.835 0.550 1.070 ;
        RECT  0.140 0.835 0.470 0.905 ;
        RECT  0.035 0.835 0.140 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 0.475 1.195 0.765 ;
        RECT  0.245 0.695 1.110 0.765 ;
        RECT  0.175 0.495 0.245 0.765 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.975 0.535 1.030 0.625 ;
        RECT  0.875 0.335 0.975 0.625 ;
        RECT  0.525 0.335 0.875 0.405 ;
        RECT  0.455 0.335 0.525 0.625 ;
        RECT  0.315 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 -0.115 1.400 0.115 ;
        RECT  1.230 -0.115 1.350 0.220 ;
        RECT  0.140 -0.115 1.230 0.115 ;
        RECT  0.070 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.145 1.400 1.375 ;
        RECT  1.040 0.975 1.120 1.375 ;
        RECT  0.740 1.145 1.040 1.375 ;
        RECT  0.660 0.975 0.740 1.375 ;
        RECT  0.350 1.145 0.660 1.375 ;
        RECT  0.270 0.975 0.350 1.375 ;
        RECT  0.000 1.145 0.270 1.375 ;
        END
    END VDD
END ND3D2BWP40

MACRO ND3D3BWP40
    CLASS CORE ;
    FOREIGN ND3D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.430500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.845 1.705 1.075 ;
        RECT  1.290 0.845 1.610 0.935 ;
        RECT  1.210 0.845 1.290 1.075 ;
        RECT  0.910 0.845 1.210 0.935 ;
        RECT  0.830 0.845 0.910 1.075 ;
        RECT  0.595 0.845 0.830 0.935 ;
        RECT  0.530 0.350 0.595 0.935 ;
        RECT  0.450 0.350 0.530 1.075 ;
        RECT  0.385 0.350 0.450 0.935 ;
        RECT  0.130 0.350 0.385 0.420 ;
        RECT  0.145 0.845 0.385 0.935 ;
        RECT  0.050 0.845 0.145 1.075 ;
        RECT  0.050 0.215 0.130 0.420 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.495 1.745 0.625 ;
        RECT  1.410 0.495 1.515 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.495 1.155 0.625 ;
        RECT  0.735 0.495 0.815 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.310 0.640 ;
        RECT  0.175 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.830 -0.115 1.910 0.425 ;
        RECT  1.510 -0.115 1.830 0.115 ;
        RECT  1.390 -0.115 1.510 0.275 ;
        RECT  0.000 -0.115 1.390 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.830 0.695 1.910 1.375 ;
        RECT  1.510 1.145 1.830 1.375 ;
        RECT  1.390 1.010 1.510 1.375 ;
        RECT  1.120 1.145 1.390 1.375 ;
        RECT  1.000 1.010 1.120 1.375 ;
        RECT  0.740 1.145 1.000 1.375 ;
        RECT  0.620 1.010 0.740 1.375 ;
        RECT  0.360 1.145 0.620 1.375 ;
        RECT  0.240 1.010 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.610 0.845 1.705 1.075 ;
        RECT  1.290 0.845 1.610 0.935 ;
        RECT  1.210 0.845 1.290 1.075 ;
        RECT  0.910 0.845 1.210 0.935 ;
        RECT  0.830 0.845 0.910 1.075 ;
        RECT  0.665 0.845 0.830 0.935 ;
        RECT  0.145 0.845 0.315 0.935 ;
        RECT  0.130 0.350 0.305 0.420 ;
        RECT  0.050 0.845 0.145 1.075 ;
        RECT  0.050 0.215 0.130 0.420 ;
        RECT  1.590 0.210 1.710 0.415 ;
        RECT  1.290 0.345 1.590 0.415 ;
        RECT  1.210 0.185 1.290 0.415 ;
        RECT  0.780 0.345 1.210 0.415 ;
        RECT  0.240 0.205 1.120 0.275 ;
    END
END ND3D3BWP40

MACRO ND3D4BWP40
    CLASS CORE ;
    FOREIGN ND3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.505450 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.320 2.625 0.905 ;
        RECT  2.410 0.320 2.555 0.390 ;
        RECT  2.345 0.735 2.555 1.055 ;
        RECT  2.340 0.195 2.410 0.390 ;
        RECT  0.130 0.985 2.345 1.055 ;
        RECT  0.615 0.195 2.340 0.265 ;
        RECT  0.035 0.745 0.130 1.055 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.460 2.485 0.640 ;
        RECT  2.215 0.460 2.380 0.530 ;
        RECT  2.135 0.335 2.215 0.530 ;
        RECT  1.365 0.335 2.135 0.405 ;
        RECT  1.265 0.335 1.365 0.630 ;
        RECT  0.270 0.335 1.265 0.405 ;
        RECT  0.175 0.335 0.270 0.625 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.113400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.230 0.600 2.270 0.710 ;
        RECT  2.135 0.600 2.230 0.915 ;
        RECT  1.725 0.845 2.135 0.915 ;
        RECT  1.590 0.615 1.725 0.915 ;
        RECT  1.045 0.845 1.590 0.915 ;
        RECT  0.915 0.615 1.045 0.915 ;
        RECT  0.525 0.845 0.915 0.915 ;
        RECT  0.450 0.520 0.525 0.915 ;
        RECT  0.370 0.520 0.450 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.113400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.795 0.475 2.065 0.625 ;
        RECT  1.520 0.475 1.795 0.545 ;
        RECT  1.435 0.475 1.520 0.775 ;
        RECT  1.185 0.705 1.435 0.775 ;
        RECT  1.115 0.475 1.185 0.775 ;
        RECT  0.845 0.475 1.115 0.545 ;
        RECT  0.595 0.475 0.845 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.600 -0.115 2.660 0.115 ;
        RECT  2.500 -0.115 2.600 0.250 ;
        RECT  1.410 -0.115 2.500 0.115 ;
        RECT  1.280 -0.115 1.410 0.125 ;
        RECT  0.120 -0.115 1.280 0.115 ;
        RECT  0.050 -0.115 0.120 0.280 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.145 2.660 1.375 ;
        RECT  2.290 1.125 2.410 1.375 ;
        RECT  2.010 1.145 2.290 1.375 ;
        RECT  1.890 1.125 2.010 1.375 ;
        RECT  1.570 1.145 1.890 1.375 ;
        RECT  1.450 1.125 1.570 1.375 ;
        RECT  1.150 1.145 1.450 1.375 ;
        RECT  1.030 1.125 1.150 1.375 ;
        RECT  0.750 1.145 1.030 1.375 ;
        RECT  0.630 1.125 0.750 1.375 ;
        RECT  0.350 1.145 0.630 1.375 ;
        RECT  0.230 1.125 0.350 1.375 ;
        RECT  0.000 1.145 0.230 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.615 0.195 2.275 0.265 ;
        RECT  0.130 0.985 2.275 1.055 ;
        RECT  0.035 0.745 0.130 1.055 ;
    END
END ND3D4BWP40

MACRO ND3D6BWP40
    CLASS CORE ;
    FOREIGN ND3D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.765000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.355 3.560 0.425 ;
        RECT  3.460 0.355 3.535 0.990 ;
        RECT  3.325 0.355 3.460 0.815 ;
        RECT  2.680 0.355 3.325 0.425 ;
        RECT  3.160 0.705 3.325 0.815 ;
        RECT  3.080 0.705 3.160 0.990 ;
        RECT  2.780 0.705 3.080 0.815 ;
        RECT  2.700 0.705 2.780 0.990 ;
        RECT  2.220 0.705 2.700 0.815 ;
        RECT  2.140 0.705 2.220 0.990 ;
        RECT  1.840 0.705 2.140 0.815 ;
        RECT  1.760 0.705 1.840 0.990 ;
        RECT  1.460 0.705 1.760 0.815 ;
        RECT  1.380 0.705 1.460 0.990 ;
        RECT  1.080 0.705 1.380 0.815 ;
        RECT  1.000 0.705 1.080 0.990 ;
        RECT  0.700 0.705 1.000 0.815 ;
        RECT  0.620 0.705 0.700 0.990 ;
        RECT  0.330 0.705 0.620 0.815 ;
        RECT  0.230 0.705 0.330 0.970 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.495 1.070 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.495 2.275 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.495 3.155 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.115 3.780 0.115 ;
        RECT  1.000 -0.115 1.080 0.285 ;
        RECT  0.700 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.700 0.285 ;
        RECT  0.320 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.320 0.285 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 1.145 3.780 1.375 ;
        RECT  3.655 0.695 3.725 1.375 ;
        RECT  3.370 1.145 3.655 1.375 ;
        RECT  3.250 0.885 3.370 1.375 ;
        RECT  2.990 1.145 3.250 1.375 ;
        RECT  2.870 0.885 2.990 1.375 ;
        RECT  2.605 1.145 2.870 1.375 ;
        RECT  2.495 0.885 2.605 1.375 ;
        RECT  2.425 1.145 2.495 1.375 ;
        RECT  2.315 0.885 2.425 1.375 ;
        RECT  2.050 1.145 2.315 1.375 ;
        RECT  1.930 0.885 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.885 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.885 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.885 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.885 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.695 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.680 0.355 3.255 0.425 ;
        RECT  3.160 0.705 3.255 0.815 ;
        RECT  3.080 0.705 3.160 0.990 ;
        RECT  2.780 0.705 3.080 0.815 ;
        RECT  2.700 0.705 2.780 0.990 ;
        RECT  2.220 0.705 2.700 0.815 ;
        RECT  2.140 0.705 2.220 0.990 ;
        RECT  1.840 0.705 2.140 0.815 ;
        RECT  1.760 0.705 1.840 0.990 ;
        RECT  1.460 0.705 1.760 0.815 ;
        RECT  1.380 0.705 1.460 0.990 ;
        RECT  1.080 0.705 1.380 0.815 ;
        RECT  1.000 0.705 1.080 0.990 ;
        RECT  0.700 0.705 1.000 0.815 ;
        RECT  0.620 0.705 0.700 0.990 ;
        RECT  0.330 0.705 0.620 0.815 ;
        RECT  0.230 0.705 0.330 0.970 ;
        RECT  0.885 0.355 1.195 0.425 ;
        RECT  0.815 0.185 0.885 0.425 ;
        RECT  0.505 0.355 0.815 0.425 ;
        RECT  0.435 0.185 0.505 0.425 ;
        RECT  0.140 0.355 0.435 0.425 ;
        RECT  0.040 0.185 0.140 0.425 ;
        RECT  3.655 0.215 3.725 0.475 ;
        RECT  1.355 0.215 3.655 0.285 ;
        RECT  1.265 0.355 2.430 0.425 ;
        RECT  1.195 0.185 1.265 0.425 ;
    END
END ND3D6BWP40

MACRO ND3D8BWP40
    CLASS CORE ;
    FOREIGN ND3D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.020000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.355 4.760 0.425 ;
        RECT  4.650 0.705 4.750 0.970 ;
        RECT  4.375 0.705 4.650 0.815 ;
        RECT  4.360 0.355 4.375 0.815 ;
        RECT  4.280 0.355 4.360 0.990 ;
        RECT  4.165 0.355 4.280 0.815 ;
        RECT  3.500 0.355 4.165 0.425 ;
        RECT  3.980 0.705 4.165 0.815 ;
        RECT  3.900 0.705 3.980 0.990 ;
        RECT  3.600 0.705 3.900 0.815 ;
        RECT  3.520 0.705 3.600 0.990 ;
        RECT  3.040 0.705 3.520 0.815 ;
        RECT  2.960 0.705 3.040 0.990 ;
        RECT  2.660 0.705 2.960 0.815 ;
        RECT  2.580 0.705 2.660 0.990 ;
        RECT  2.280 0.705 2.580 0.815 ;
        RECT  2.200 0.705 2.280 0.990 ;
        RECT  1.900 0.705 2.200 0.815 ;
        RECT  1.820 0.705 1.900 0.990 ;
        RECT  1.520 0.705 1.820 0.815 ;
        RECT  1.440 0.705 1.520 0.990 ;
        RECT  1.140 0.705 1.440 0.815 ;
        RECT  1.060 0.705 1.140 0.990 ;
        RECT  0.760 0.705 1.060 0.815 ;
        RECT  0.680 0.705 0.760 0.990 ;
        RECT  0.390 0.705 0.680 0.815 ;
        RECT  0.290 0.705 0.390 0.970 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.215 0.495 1.475 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 0.495 3.095 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.455 0.495 3.975 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.115 5.040 0.115 ;
        RECT  1.440 -0.115 1.520 0.285 ;
        RECT  1.140 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.140 0.285 ;
        RECT  0.760 -0.115 1.060 0.115 ;
        RECT  0.680 -0.115 0.760 0.285 ;
        RECT  0.380 -0.115 0.680 0.115 ;
        RECT  0.300 -0.115 0.380 0.285 ;
        RECT  0.000 -0.115 0.300 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.950 1.145 5.040 1.375 ;
        RECT  4.880 0.695 4.950 1.375 ;
        RECT  4.570 1.145 4.880 1.375 ;
        RECT  4.450 0.885 4.570 1.375 ;
        RECT  4.190 1.145 4.450 1.375 ;
        RECT  4.070 0.885 4.190 1.375 ;
        RECT  3.810 1.145 4.070 1.375 ;
        RECT  3.690 0.885 3.810 1.375 ;
        RECT  3.425 1.145 3.690 1.375 ;
        RECT  3.315 0.885 3.425 1.375 ;
        RECT  3.245 1.145 3.315 1.375 ;
        RECT  3.135 0.885 3.245 1.375 ;
        RECT  2.870 1.145 3.135 1.375 ;
        RECT  2.750 0.885 2.870 1.375 ;
        RECT  2.490 1.145 2.750 1.375 ;
        RECT  2.370 0.885 2.490 1.375 ;
        RECT  2.110 1.145 2.370 1.375 ;
        RECT  1.990 0.885 2.110 1.375 ;
        RECT  1.730 1.145 1.990 1.375 ;
        RECT  1.610 0.885 1.730 1.375 ;
        RECT  1.350 1.145 1.610 1.375 ;
        RECT  1.230 0.885 1.350 1.375 ;
        RECT  0.970 1.145 1.230 1.375 ;
        RECT  0.850 0.885 0.970 1.375 ;
        RECT  0.590 1.145 0.850 1.375 ;
        RECT  0.470 0.885 0.590 1.375 ;
        RECT  0.190 1.145 0.470 1.375 ;
        RECT  0.090 0.695 0.190 1.375 ;
        RECT  0.000 1.145 0.090 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.355 4.760 0.425 ;
        RECT  4.650 0.705 4.750 0.970 ;
        RECT  4.445 0.705 4.650 0.815 ;
        RECT  3.500 0.355 4.095 0.425 ;
        RECT  3.980 0.705 4.095 0.815 ;
        RECT  3.900 0.705 3.980 0.990 ;
        RECT  3.600 0.705 3.900 0.815 ;
        RECT  3.520 0.705 3.600 0.990 ;
        RECT  3.040 0.705 3.520 0.815 ;
        RECT  2.960 0.705 3.040 0.990 ;
        RECT  2.660 0.705 2.960 0.815 ;
        RECT  2.580 0.705 2.660 0.990 ;
        RECT  2.280 0.705 2.580 0.815 ;
        RECT  2.200 0.705 2.280 0.990 ;
        RECT  1.900 0.705 2.200 0.815 ;
        RECT  1.820 0.705 1.900 0.990 ;
        RECT  1.520 0.705 1.820 0.815 ;
        RECT  1.440 0.705 1.520 0.990 ;
        RECT  1.140 0.705 1.440 0.815 ;
        RECT  1.060 0.705 1.140 0.990 ;
        RECT  0.760 0.705 1.060 0.815 ;
        RECT  0.680 0.705 0.760 0.990 ;
        RECT  0.390 0.705 0.680 0.815 ;
        RECT  0.290 0.705 0.390 0.970 ;
        RECT  4.880 0.215 4.950 0.475 ;
        RECT  1.800 0.215 4.880 0.285 ;
        RECT  4.490 0.550 4.820 0.625 ;
        RECT  1.705 0.355 3.250 0.425 ;
        RECT  1.635 0.185 1.705 0.425 ;
        RECT  1.325 0.355 1.635 0.425 ;
        RECT  1.255 0.185 1.325 0.425 ;
        RECT  0.945 0.355 1.255 0.425 ;
        RECT  0.875 0.185 0.945 0.425 ;
        RECT  0.565 0.355 0.875 0.425 ;
        RECT  0.495 0.185 0.565 0.425 ;
        RECT  0.200 0.355 0.495 0.425 ;
        RECT  0.100 0.185 0.200 0.425 ;
    END
END ND3D8BWP40

MACRO ND4D0BWP40
    CLASS CORE ;
    FOREIGN ND4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.093875 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 0.810 ;
        RECT  0.810 0.195 0.875 0.265 ;
        RECT  0.720 0.740 0.875 0.810 ;
        RECT  0.640 0.740 0.720 1.035 ;
        RECT  0.320 0.740 0.640 0.810 ;
        RECT  0.245 0.740 0.320 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.625 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.980 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.820 1.020 0.940 1.375 ;
        RECT  0.540 1.145 0.820 1.375 ;
        RECT  0.420 1.020 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.985 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND4D0BWP40

MACRO ND4D1BWP40
    CLASS CORE ;
    FOREIGN ND4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.187750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 0.810 ;
        RECT  0.810 0.195 0.875 0.265 ;
        RECT  0.720 0.740 0.875 0.810 ;
        RECT  0.640 0.740 0.720 1.035 ;
        RECT  0.320 0.740 0.640 0.810 ;
        RECT  0.245 0.740 0.320 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.345 0.385 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.625 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 -0.115 0.980 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.820 0.880 0.940 1.375 ;
        RECT  0.540 1.145 0.820 1.375 ;
        RECT  0.420 0.880 0.540 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END ND4D1BWP40

MACRO ND4D2BWP40
    CLASS CORE ;
    FOREIGN ND4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.322500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.835 1.690 1.075 ;
        RECT  1.300 0.835 1.590 0.905 ;
        RECT  1.220 0.835 1.300 1.075 ;
        RECT  0.740 0.835 1.220 0.905 ;
        RECT  0.660 0.835 0.740 1.075 ;
        RECT  0.385 0.835 0.660 0.905 ;
        RECT  0.355 0.345 0.385 0.905 ;
        RECT  0.315 0.345 0.355 1.035 ;
        RECT  0.260 0.345 0.315 0.415 ;
        RECT  0.285 0.735 0.315 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.495 1.785 0.625 ;
        RECT  1.570 0.495 1.655 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.285 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.285 0.615 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.775 0.615 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.355 0.105 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.680 -0.115 1.960 0.115 ;
        RECT  1.600 -0.115 1.680 0.285 ;
        RECT  0.000 -0.115 1.600 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.810 0.705 1.910 1.375 ;
        RECT  1.490 1.145 1.810 1.375 ;
        RECT  1.410 0.975 1.490 1.375 ;
        RECT  1.110 1.145 1.410 1.375 ;
        RECT  1.030 0.975 1.110 1.375 ;
        RECT  0.930 1.145 1.030 1.375 ;
        RECT  0.850 0.975 0.930 1.375 ;
        RECT  0.550 1.145 0.850 1.375 ;
        RECT  0.470 0.975 0.550 1.375 ;
        RECT  0.150 1.145 0.470 1.375 ;
        RECT  0.050 0.730 0.150 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.810 0.185 1.910 0.425 ;
        RECT  1.490 0.355 1.810 0.425 ;
        RECT  1.410 0.195 1.490 0.425 ;
        RECT  1.015 0.195 1.410 0.265 ;
        RECT  0.635 0.355 1.320 0.425 ;
        RECT  0.545 0.195 0.945 0.265 ;
        RECT  0.475 0.195 0.545 0.425 ;
        RECT  0.040 0.195 0.475 0.265 ;
    END
END ND4D2BWP40

MACRO ND4D3BWP40
    CLASS CORE ;
    FOREIGN ND4D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.567750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 0.700 2.450 1.035 ;
        RECT  2.050 0.700 2.370 0.815 ;
        RECT  1.970 0.700 2.050 1.035 ;
        RECT  1.670 0.700 1.970 0.815 ;
        RECT  1.590 0.700 1.670 1.035 ;
        RECT  1.290 0.700 1.590 0.815 ;
        RECT  1.210 0.700 1.290 1.035 ;
        RECT  0.910 0.700 1.210 0.815 ;
        RECT  0.830 0.700 0.910 1.035 ;
        RECT  0.825 0.700 0.830 0.960 ;
        RECT  0.595 0.845 0.825 0.960 ;
        RECT  0.530 0.355 0.595 0.960 ;
        RECT  0.450 0.355 0.530 1.065 ;
        RECT  0.385 0.355 0.450 0.960 ;
        RECT  0.160 0.355 0.385 0.425 ;
        RECT  0.150 0.845 0.385 0.960 ;
        RECT  0.060 0.185 0.160 0.425 ;
        RECT  0.070 0.845 0.150 1.035 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.955 0.495 2.345 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.725 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.140 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.305 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 -0.115 2.520 0.115 ;
        RECT  2.370 -0.115 2.450 0.425 ;
        RECT  2.070 -0.115 2.370 0.115 ;
        RECT  1.950 -0.115 2.070 0.285 ;
        RECT  0.000 -0.115 1.950 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.145 2.520 1.375 ;
        RECT  2.140 0.885 2.260 1.375 ;
        RECT  1.880 1.145 2.140 1.375 ;
        RECT  1.760 0.885 1.880 1.375 ;
        RECT  1.500 1.145 1.760 1.375 ;
        RECT  1.380 0.885 1.500 1.375 ;
        RECT  1.120 1.145 1.380 1.375 ;
        RECT  1.000 0.885 1.120 1.375 ;
        RECT  0.740 1.145 1.000 1.375 ;
        RECT  0.620 1.030 0.740 1.375 ;
        RECT  0.360 1.145 0.620 1.375 ;
        RECT  0.240 1.030 0.360 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.370 0.700 2.450 1.035 ;
        RECT  2.050 0.700 2.370 0.815 ;
        RECT  1.970 0.700 2.050 1.035 ;
        RECT  1.670 0.700 1.970 0.815 ;
        RECT  1.590 0.700 1.670 1.035 ;
        RECT  1.290 0.700 1.590 0.815 ;
        RECT  1.210 0.700 1.290 1.035 ;
        RECT  0.910 0.700 1.210 0.815 ;
        RECT  0.830 0.700 0.910 1.035 ;
        RECT  0.825 0.700 0.830 0.960 ;
        RECT  0.665 0.845 0.825 0.960 ;
        RECT  0.160 0.355 0.315 0.425 ;
        RECT  0.150 0.845 0.315 0.960 ;
        RECT  0.060 0.185 0.160 0.425 ;
        RECT  0.070 0.845 0.150 1.035 ;
        RECT  2.150 0.185 2.250 0.425 ;
        RECT  1.860 0.355 2.150 0.425 ;
        RECT  1.780 0.215 1.860 0.425 ;
        RECT  1.380 0.215 1.780 0.285 ;
        RECT  1.290 0.355 1.690 0.425 ;
        RECT  1.210 0.190 1.290 0.425 ;
        RECT  0.780 0.355 1.210 0.425 ;
        RECT  0.240 0.205 1.120 0.275 ;
    END
END ND4D3BWP40

MACRO ND4D4BWP40
    CLASS CORE ;
    FOREIGN ND4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.615000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.185 0.700 3.255 1.020 ;
        RECT  2.875 0.700 3.185 0.815 ;
        RECT  2.805 0.700 2.875 1.020 ;
        RECT  2.495 0.700 2.805 0.815 ;
        RECT  2.425 0.700 2.495 1.020 ;
        RECT  2.115 0.700 2.425 0.815 ;
        RECT  2.045 0.700 2.115 1.020 ;
        RECT  1.455 0.700 2.045 0.815 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.075 0.700 1.385 0.815 ;
        RECT  1.005 0.700 1.075 1.020 ;
        RECT  0.695 0.700 1.005 0.815 ;
        RECT  0.595 0.345 0.720 0.430 ;
        RECT  0.625 0.700 0.695 1.020 ;
        RECT  0.595 0.700 0.625 0.815 ;
        RECT  0.385 0.345 0.595 0.815 ;
        RECT  0.220 0.345 0.385 0.430 ;
        RECT  0.315 0.700 0.385 0.815 ;
        RECT  0.245 0.700 0.315 1.020 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.495 3.325 0.630 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.555 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.495 1.460 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.545 0.255 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.115 3.500 0.115 ;
        RECT  3.160 -0.115 3.280 0.275 ;
        RECT  2.900 -0.115 3.160 0.115 ;
        RECT  2.780 -0.115 2.900 0.275 ;
        RECT  0.000 -0.115 2.780 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 1.145 3.500 1.375 ;
        RECT  3.375 0.700 3.445 1.375 ;
        RECT  3.090 1.145 3.375 1.375 ;
        RECT  2.970 0.885 3.090 1.375 ;
        RECT  2.710 1.145 2.970 1.375 ;
        RECT  2.590 0.885 2.710 1.375 ;
        RECT  2.330 1.145 2.590 1.375 ;
        RECT  2.210 0.885 2.330 1.375 ;
        RECT  1.950 1.145 2.210 1.375 ;
        RECT  1.830 0.885 1.950 1.375 ;
        RECT  1.670 1.145 1.830 1.375 ;
        RECT  1.550 0.885 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.885 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.885 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.885 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.185 0.700 3.255 1.020 ;
        RECT  2.875 0.700 3.185 0.815 ;
        RECT  2.805 0.700 2.875 1.020 ;
        RECT  2.495 0.700 2.805 0.815 ;
        RECT  2.425 0.700 2.495 1.020 ;
        RECT  2.115 0.700 2.425 0.815 ;
        RECT  2.045 0.700 2.115 1.020 ;
        RECT  1.455 0.700 2.045 0.815 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.075 0.700 1.385 0.815 ;
        RECT  1.005 0.700 1.075 1.020 ;
        RECT  0.695 0.700 1.005 0.815 ;
        RECT  0.665 0.345 0.720 0.430 ;
        RECT  0.665 0.700 0.695 1.020 ;
        RECT  0.220 0.345 0.315 0.430 ;
        RECT  0.245 0.700 0.315 1.020 ;
        RECT  3.360 0.185 3.460 0.425 ;
        RECT  3.070 0.355 3.360 0.425 ;
        RECT  2.990 0.190 3.070 0.425 ;
        RECT  2.690 0.355 2.990 0.425 ;
        RECT  2.610 0.190 2.690 0.425 ;
        RECT  1.830 0.355 2.610 0.425 ;
        RECT  0.980 0.205 2.520 0.275 ;
        RECT  0.885 0.345 1.670 0.415 ;
        RECT  0.815 0.205 0.885 0.415 ;
        RECT  0.130 0.205 0.815 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END ND4D4BWP40

MACRO ND4D6BWP40
    CLASS CORE ;
    FOREIGN ND4D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.922500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.700 4.795 1.020 ;
        RECT  4.415 0.700 4.725 0.815 ;
        RECT  4.345 0.700 4.415 1.020 ;
        RECT  4.035 0.700 4.345 0.815 ;
        RECT  3.965 0.700 4.035 1.020 ;
        RECT  3.655 0.700 3.965 0.815 ;
        RECT  3.585 0.700 3.655 1.020 ;
        RECT  3.275 0.700 3.585 0.815 ;
        RECT  3.205 0.700 3.275 1.020 ;
        RECT  2.895 0.700 3.205 0.815 ;
        RECT  2.825 0.700 2.895 1.020 ;
        RECT  2.230 0.700 2.825 0.815 ;
        RECT  2.145 0.700 2.230 1.020 ;
        RECT  1.835 0.700 2.145 0.815 ;
        RECT  1.765 0.700 1.835 1.020 ;
        RECT  1.455 0.700 1.765 0.815 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.075 0.700 1.385 0.815 ;
        RECT  0.595 0.345 1.100 0.420 ;
        RECT  1.005 0.700 1.075 1.020 ;
        RECT  0.695 0.700 1.005 0.815 ;
        RECT  0.625 0.700 0.695 1.020 ;
        RECT  0.595 0.700 0.625 0.815 ;
        RECT  0.385 0.345 0.595 0.815 ;
        RECT  0.220 0.345 0.385 0.430 ;
        RECT  0.315 0.700 0.385 0.815 ;
        RECT  0.245 0.700 0.315 1.020 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.955 0.495 4.865 0.630 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.495 3.745 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 2.265 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.495 1.145 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.820 0.275 ;
        RECT  4.440 -0.115 4.700 0.115 ;
        RECT  4.320 -0.115 4.440 0.275 ;
        RECT  4.060 -0.115 4.320 0.115 ;
        RECT  3.940 -0.115 4.060 0.275 ;
        RECT  0.000 -0.115 3.940 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 1.145 5.040 1.375 ;
        RECT  4.915 0.700 4.985 1.375 ;
        RECT  4.630 1.145 4.915 1.375 ;
        RECT  4.510 0.885 4.630 1.375 ;
        RECT  4.250 1.145 4.510 1.375 ;
        RECT  4.130 0.885 4.250 1.375 ;
        RECT  3.870 1.145 4.130 1.375 ;
        RECT  3.750 0.885 3.870 1.375 ;
        RECT  3.490 1.145 3.750 1.375 ;
        RECT  3.370 0.885 3.490 1.375 ;
        RECT  3.110 1.145 3.370 1.375 ;
        RECT  2.990 0.885 3.110 1.375 ;
        RECT  2.730 1.145 2.990 1.375 ;
        RECT  2.610 0.885 2.730 1.375 ;
        RECT  2.450 1.145 2.610 1.375 ;
        RECT  2.325 0.885 2.450 1.375 ;
        RECT  2.050 1.145 2.325 1.375 ;
        RECT  1.930 0.885 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.885 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.885 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.885 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.885 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.705 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.700 4.795 1.020 ;
        RECT  4.415 0.700 4.725 0.815 ;
        RECT  4.345 0.700 4.415 1.020 ;
        RECT  4.035 0.700 4.345 0.815 ;
        RECT  3.965 0.700 4.035 1.020 ;
        RECT  3.655 0.700 3.965 0.815 ;
        RECT  3.585 0.700 3.655 1.020 ;
        RECT  3.275 0.700 3.585 0.815 ;
        RECT  3.205 0.700 3.275 1.020 ;
        RECT  2.895 0.700 3.205 0.815 ;
        RECT  2.825 0.700 2.895 1.020 ;
        RECT  2.230 0.700 2.825 0.815 ;
        RECT  2.145 0.700 2.230 1.020 ;
        RECT  1.835 0.700 2.145 0.815 ;
        RECT  1.765 0.700 1.835 1.020 ;
        RECT  1.455 0.700 1.765 0.815 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.075 0.700 1.385 0.815 ;
        RECT  0.665 0.345 1.100 0.420 ;
        RECT  1.005 0.700 1.075 1.020 ;
        RECT  0.695 0.700 1.005 0.815 ;
        RECT  0.665 0.700 0.695 1.020 ;
        RECT  0.220 0.345 0.315 0.430 ;
        RECT  0.245 0.700 0.315 1.020 ;
        RECT  4.900 0.185 5.000 0.425 ;
        RECT  4.610 0.355 4.900 0.425 ;
        RECT  4.530 0.190 4.610 0.425 ;
        RECT  4.230 0.355 4.530 0.425 ;
        RECT  4.150 0.190 4.230 0.425 ;
        RECT  3.850 0.355 4.150 0.425 ;
        RECT  3.770 0.190 3.850 0.425 ;
        RECT  2.610 0.355 3.770 0.425 ;
        RECT  1.360 0.205 3.680 0.275 ;
        RECT  1.265 0.345 2.450 0.415 ;
        RECT  1.195 0.205 1.265 0.415 ;
        RECT  0.130 0.205 1.195 0.275 ;
        RECT  0.050 0.205 0.130 0.455 ;
    END
END ND4D6BWP40

MACRO ND4D8BWP40
    CLASS CORE ;
    FOREIGN ND4D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.230000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.245 0.700 6.315 1.020 ;
        RECT  5.935 0.700 6.245 0.815 ;
        RECT  5.865 0.700 5.935 1.020 ;
        RECT  5.555 0.700 5.865 0.815 ;
        RECT  5.485 0.700 5.555 1.020 ;
        RECT  5.175 0.700 5.485 0.815 ;
        RECT  5.105 0.700 5.175 1.020 ;
        RECT  4.795 0.700 5.105 0.815 ;
        RECT  4.725 0.700 4.795 1.020 ;
        RECT  4.415 0.700 4.725 0.815 ;
        RECT  4.345 0.700 4.415 1.020 ;
        RECT  4.035 0.700 4.345 0.815 ;
        RECT  3.965 0.700 4.035 1.020 ;
        RECT  3.655 0.700 3.965 0.815 ;
        RECT  3.585 0.700 3.655 1.020 ;
        RECT  2.975 0.700 3.585 0.815 ;
        RECT  2.905 0.700 2.975 1.020 ;
        RECT  2.595 0.700 2.905 0.815 ;
        RECT  2.525 0.700 2.595 1.020 ;
        RECT  2.215 0.700 2.525 0.815 ;
        RECT  2.145 0.700 2.215 1.020 ;
        RECT  1.835 0.700 2.145 0.815 ;
        RECT  1.765 0.700 1.835 1.020 ;
        RECT  1.455 0.700 1.765 0.815 ;
        RECT  1.015 0.345 1.480 0.425 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.075 0.700 1.385 0.815 ;
        RECT  1.015 0.700 1.075 1.045 ;
        RECT  1.005 0.345 1.015 1.045 ;
        RECT  0.805 0.345 1.005 0.815 ;
        RECT  0.220 0.345 0.805 0.425 ;
        RECT  0.695 0.700 0.805 0.815 ;
        RECT  0.625 0.700 0.695 1.020 ;
        RECT  0.315 0.700 0.625 0.815 ;
        RECT  0.245 0.700 0.315 1.020 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 0.495 6.405 0.630 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.530 0.495 4.865 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.675 0.495 2.995 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.495 0.680 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.340 -0.115 6.580 0.115 ;
        RECT  6.220 -0.115 6.340 0.275 ;
        RECT  5.960 -0.115 6.220 0.115 ;
        RECT  5.840 -0.115 5.960 0.275 ;
        RECT  5.580 -0.115 5.840 0.115 ;
        RECT  5.460 -0.115 5.580 0.275 ;
        RECT  5.200 -0.115 5.460 0.115 ;
        RECT  5.080 -0.115 5.200 0.275 ;
        RECT  0.000 -0.115 5.080 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 1.145 6.580 1.375 ;
        RECT  6.455 0.700 6.525 1.375 ;
        RECT  6.150 1.145 6.455 1.375 ;
        RECT  6.030 0.885 6.150 1.375 ;
        RECT  5.770 1.145 6.030 1.375 ;
        RECT  5.650 0.885 5.770 1.375 ;
        RECT  5.390 1.145 5.650 1.375 ;
        RECT  5.270 0.885 5.390 1.375 ;
        RECT  5.010 1.145 5.270 1.375 ;
        RECT  4.890 0.885 5.010 1.375 ;
        RECT  4.630 1.145 4.890 1.375 ;
        RECT  4.510 0.885 4.630 1.375 ;
        RECT  4.250 1.145 4.510 1.375 ;
        RECT  4.130 0.885 4.250 1.375 ;
        RECT  3.870 1.145 4.130 1.375 ;
        RECT  3.750 0.885 3.870 1.375 ;
        RECT  3.490 1.145 3.750 1.375 ;
        RECT  3.370 0.885 3.490 1.375 ;
        RECT  3.190 1.145 3.370 1.375 ;
        RECT  3.070 0.885 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.885 2.810 1.375 ;
        RECT  2.430 1.145 2.690 1.375 ;
        RECT  2.310 0.885 2.430 1.375 ;
        RECT  2.050 1.145 2.310 1.375 ;
        RECT  1.930 0.885 2.050 1.375 ;
        RECT  1.670 1.145 1.930 1.375 ;
        RECT  1.550 0.885 1.670 1.375 ;
        RECT  1.290 1.145 1.550 1.375 ;
        RECT  1.170 0.885 1.290 1.375 ;
        RECT  0.910 1.145 1.170 1.375 ;
        RECT  0.790 0.885 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 0.885 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.705 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.245 0.700 6.315 1.020 ;
        RECT  5.935 0.700 6.245 0.815 ;
        RECT  5.865 0.700 5.935 1.020 ;
        RECT  5.555 0.700 5.865 0.815 ;
        RECT  5.485 0.700 5.555 1.020 ;
        RECT  5.175 0.700 5.485 0.815 ;
        RECT  5.105 0.700 5.175 1.020 ;
        RECT  4.795 0.700 5.105 0.815 ;
        RECT  4.725 0.700 4.795 1.020 ;
        RECT  4.415 0.700 4.725 0.815 ;
        RECT  4.345 0.700 4.415 1.020 ;
        RECT  4.035 0.700 4.345 0.815 ;
        RECT  3.965 0.700 4.035 1.020 ;
        RECT  3.655 0.700 3.965 0.815 ;
        RECT  3.585 0.700 3.655 1.020 ;
        RECT  2.975 0.700 3.585 0.815 ;
        RECT  2.905 0.700 2.975 1.020 ;
        RECT  2.595 0.700 2.905 0.815 ;
        RECT  2.525 0.700 2.595 1.020 ;
        RECT  2.215 0.700 2.525 0.815 ;
        RECT  2.145 0.700 2.215 1.020 ;
        RECT  1.835 0.700 2.145 0.815 ;
        RECT  1.765 0.700 1.835 1.020 ;
        RECT  1.455 0.700 1.765 0.815 ;
        RECT  1.085 0.345 1.480 0.425 ;
        RECT  1.385 0.700 1.455 1.020 ;
        RECT  1.085 0.700 1.385 0.815 ;
        RECT  0.220 0.345 0.735 0.425 ;
        RECT  0.695 0.700 0.735 0.815 ;
        RECT  0.625 0.700 0.695 1.020 ;
        RECT  0.315 0.700 0.625 0.815 ;
        RECT  0.245 0.700 0.315 1.020 ;
        RECT  6.440 0.185 6.540 0.425 ;
        RECT  6.130 0.355 6.440 0.425 ;
        RECT  6.050 0.190 6.130 0.425 ;
        RECT  5.750 0.355 6.050 0.425 ;
        RECT  5.670 0.190 5.750 0.425 ;
        RECT  5.370 0.355 5.670 0.425 ;
        RECT  5.290 0.190 5.370 0.425 ;
        RECT  4.990 0.355 5.290 0.425 ;
        RECT  4.910 0.190 4.990 0.425 ;
        RECT  3.370 0.355 4.910 0.425 ;
        RECT  1.740 0.205 4.820 0.275 ;
        RECT  1.645 0.345 3.190 0.415 ;
        RECT  1.575 0.205 1.645 0.415 ;
        RECT  0.130 0.205 1.575 0.275 ;
        RECT  1.090 0.495 1.560 0.615 ;
        RECT  0.050 0.205 0.130 0.455 ;
    END
END ND4D8BWP40

MACRO NR2D0BWP40
    CLASS CORE ;
    FOREIGN NR2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.052125 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.325 0.525 1.045 ;
        RECT  0.325 0.325 0.455 0.395 ;
        RECT  0.435 0.915 0.455 1.045 ;
        RECT  0.235 0.210 0.325 0.395 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.255 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.145 0.560 1.375 ;
        RECT  0.050 0.950 0.125 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END NR2D0BWP40

MACRO NR2D12BWP40
    CLASS CORE ;
    FOREIGN NR2D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.999000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 0.210 4.515 0.370 ;
        RECT  4.340 0.210 4.420 0.915 ;
        RECT  3.480 0.210 4.340 0.280 ;
        RECT  4.230 0.845 4.340 0.915 ;
        RECT  3.480 0.845 3.570 0.915 ;
        RECT  3.410 0.210 3.480 0.915 ;
        RECT  2.850 0.210 3.410 0.370 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  1.995 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.995 0.835 2.065 0.915 ;
        RECT  1.910 0.210 1.995 0.915 ;
        RECT  1.785 0.210 1.910 0.625 ;
        RECT  1.350 0.210 1.785 0.350 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.348800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 0.495 4.680 0.625 ;
        RECT  4.490 0.495 4.570 1.065 ;
        RECT  4.135 0.995 4.490 1.065 ;
        RECT  4.065 0.845 4.135 1.065 ;
        RECT  3.940 0.845 4.065 0.915 ;
        RECT  3.815 0.495 3.940 0.915 ;
        RECT  3.745 0.845 3.815 0.915 ;
        RECT  3.665 0.845 3.745 1.065 ;
        RECT  3.330 0.995 3.665 1.065 ;
        RECT  3.255 0.495 3.330 1.065 ;
        RECT  3.000 0.495 3.255 0.625 ;
        RECT  2.930 0.495 3.000 1.055 ;
        RECT  2.590 0.985 2.930 1.055 ;
        RECT  2.510 0.845 2.590 1.055 ;
        RECT  2.445 0.845 2.510 0.915 ;
        RECT  2.345 0.525 2.445 0.915 ;
        RECT  2.230 0.845 2.345 0.915 ;
        RECT  2.135 0.845 2.230 1.065 ;
        RECT  1.790 0.995 2.135 1.065 ;
        RECT  1.715 0.710 1.790 1.065 ;
        RECT  1.655 0.710 1.715 0.780 ;
        RECT  1.575 0.495 1.655 0.780 ;
        RECT  1.505 0.710 1.575 0.780 ;
        RECT  1.435 0.710 1.505 1.055 ;
        RECT  1.085 0.985 1.435 1.055 ;
        RECT  0.990 0.845 1.085 1.055 ;
        RECT  0.845 0.845 0.990 0.915 ;
        RECT  0.735 0.495 0.845 0.915 ;
        RECT  0.710 0.845 0.735 0.915 ;
        RECT  0.630 0.845 0.710 1.055 ;
        RECT  0.290 0.985 0.630 1.055 ;
        RECT  0.220 0.495 0.290 1.055 ;
        RECT  0.160 0.495 0.220 0.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.374400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.350 1.085 0.625 ;
        RECT  0.665 0.350 1.015 0.420 ;
        RECT  0.525 0.350 0.665 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.720 -0.115 4.760 0.115 ;
        RECT  4.620 -0.115 4.720 0.410 ;
        RECT  4.350 -0.115 4.620 0.115 ;
        RECT  4.230 -0.115 4.350 0.140 ;
        RECT  3.960 -0.115 4.230 0.115 ;
        RECT  3.840 -0.115 3.960 0.140 ;
        RECT  3.570 -0.115 3.840 0.115 ;
        RECT  3.450 -0.115 3.570 0.140 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.140 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.140 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.140 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.140 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.140 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.140 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.145 4.760 1.375 ;
        RECT  4.640 0.720 4.710 1.375 ;
        RECT  3.960 1.145 4.640 1.375 ;
        RECT  3.840 0.985 3.960 1.375 ;
        RECT  3.180 1.145 3.840 1.375 ;
        RECT  3.080 0.845 3.180 1.375 ;
        RECT  2.420 1.145 3.080 1.375 ;
        RECT  2.320 0.985 2.420 1.375 ;
        RECT  1.645 1.145 2.320 1.375 ;
        RECT  1.575 0.860 1.645 1.375 ;
        RECT  0.900 1.145 1.575 1.375 ;
        RECT  0.800 0.985 0.900 1.375 ;
        RECT  0.140 1.145 0.800 1.375 ;
        RECT  0.040 0.730 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.420 0.210 4.515 0.370 ;
        RECT  4.340 0.210 4.420 0.915 ;
        RECT  3.480 0.210 4.340 0.280 ;
        RECT  4.230 0.845 4.340 0.915 ;
        RECT  3.480 0.845 3.570 0.915 ;
        RECT  3.410 0.210 3.480 0.915 ;
        RECT  2.850 0.210 3.410 0.370 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  2.065 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.350 0.210 1.715 0.350 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        RECT  4.195 0.520 4.220 0.665 ;
        RECT  4.105 0.350 4.195 0.665 ;
        RECT  3.725 0.350 4.105 0.420 ;
        RECT  3.650 0.350 3.725 0.630 ;
        RECT  3.550 0.510 3.650 0.630 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.350 2.595 0.640 ;
        RECT  2.215 0.350 2.525 0.420 ;
        RECT  2.145 0.350 2.215 0.665 ;
        RECT  2.070 0.495 2.145 0.665 ;
    END
END NR2D12BWP40

MACRO NR2D16BWP40
    CLASS CORE ;
    FOREIGN NR2D16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.335300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.960 0.210 6.055 0.370 ;
        RECT  5.880 0.210 5.960 0.915 ;
        RECT  5.020 0.210 5.880 0.280 ;
        RECT  5.770 0.845 5.880 0.915 ;
        RECT  5.020 0.845 5.110 0.915 ;
        RECT  4.950 0.210 5.020 0.915 ;
        RECT  4.390 0.210 4.950 0.370 ;
        RECT  4.310 0.210 4.390 0.915 ;
        RECT  3.535 0.210 4.310 0.280 ;
        RECT  4.230 0.835 4.310 0.915 ;
        RECT  3.535 0.835 3.605 0.915 ;
        RECT  3.450 0.210 3.535 0.915 ;
        RECT  3.325 0.210 3.450 0.625 ;
        RECT  2.890 0.210 3.325 0.350 ;
        RECT  2.810 0.210 2.890 0.915 ;
        RECT  1.980 0.210 2.810 0.280 ;
        RECT  2.710 0.835 2.810 0.915 ;
        RECT  1.980 0.835 2.070 0.915 ;
        RECT  1.900 0.210 1.980 0.915 ;
        RECT  1.355 0.210 1.900 0.370 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.190 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.460800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.110 0.495 6.205 0.625 ;
        RECT  6.030 0.495 6.110 1.065 ;
        RECT  5.675 0.995 6.030 1.065 ;
        RECT  5.605 0.845 5.675 1.065 ;
        RECT  5.480 0.845 5.605 0.915 ;
        RECT  5.355 0.495 5.480 0.915 ;
        RECT  5.285 0.845 5.355 0.915 ;
        RECT  5.205 0.845 5.285 1.065 ;
        RECT  4.870 0.995 5.205 1.065 ;
        RECT  4.795 0.495 4.870 1.065 ;
        RECT  4.540 0.495 4.795 0.625 ;
        RECT  4.470 0.495 4.540 1.055 ;
        RECT  4.130 0.985 4.470 1.055 ;
        RECT  4.050 0.845 4.130 1.055 ;
        RECT  3.985 0.845 4.050 0.915 ;
        RECT  3.885 0.525 3.985 0.915 ;
        RECT  3.770 0.845 3.885 0.915 ;
        RECT  3.675 0.845 3.770 1.065 ;
        RECT  3.330 0.995 3.675 1.065 ;
        RECT  3.255 0.710 3.330 1.065 ;
        RECT  3.195 0.710 3.255 0.780 ;
        RECT  3.115 0.495 3.195 0.780 ;
        RECT  3.045 0.710 3.115 0.780 ;
        RECT  2.975 0.710 3.045 1.055 ;
        RECT  2.625 0.985 2.975 1.055 ;
        RECT  2.530 0.845 2.625 1.055 ;
        RECT  2.385 0.845 2.530 0.915 ;
        RECT  2.275 0.495 2.385 0.915 ;
        RECT  2.250 0.845 2.275 0.915 ;
        RECT  2.170 0.845 2.250 1.055 ;
        RECT  1.830 0.985 2.170 1.055 ;
        RECT  1.760 0.495 1.830 1.055 ;
        RECT  1.515 0.495 1.760 0.665 ;
        RECT  1.435 0.495 1.515 1.065 ;
        RECT  1.095 0.995 1.435 1.065 ;
        RECT  1.015 0.845 1.095 1.065 ;
        RECT  0.945 0.845 1.015 0.915 ;
        RECT  0.735 0.495 0.945 0.915 ;
        RECT  0.695 0.845 0.735 0.915 ;
        RECT  0.625 0.845 0.695 1.065 ;
        RECT  0.270 0.995 0.625 1.065 ;
        RECT  0.190 0.495 0.270 1.065 ;
        RECT  0.080 0.495 0.190 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.499200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.740 0.625 ;
        RECT  2.555 0.350 2.625 0.625 ;
        RECT  2.205 0.350 2.555 0.420 ;
        RECT  2.065 0.350 2.205 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.260 -0.115 6.300 0.115 ;
        RECT  6.160 -0.115 6.260 0.410 ;
        RECT  5.890 -0.115 6.160 0.115 ;
        RECT  5.770 -0.115 5.890 0.140 ;
        RECT  5.500 -0.115 5.770 0.115 ;
        RECT  5.380 -0.115 5.500 0.140 ;
        RECT  5.110 -0.115 5.380 0.115 ;
        RECT  4.990 -0.115 5.110 0.140 ;
        RECT  4.730 -0.115 4.990 0.115 ;
        RECT  4.610 -0.115 4.730 0.140 ;
        RECT  4.350 -0.115 4.610 0.115 ;
        RECT  4.230 -0.115 4.350 0.140 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.140 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.140 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.140 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.140 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.140 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.140 ;
        RECT  1.695 -0.115 1.950 0.115 ;
        RECT  1.565 -0.115 1.695 0.140 ;
        RECT  1.310 -0.115 1.565 0.115 ;
        RECT  1.190 -0.115 1.310 0.140 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.920 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.145 6.300 1.375 ;
        RECT  6.180 0.720 6.250 1.375 ;
        RECT  5.500 1.145 6.180 1.375 ;
        RECT  5.380 0.985 5.500 1.375 ;
        RECT  4.720 1.145 5.380 1.375 ;
        RECT  4.620 0.845 4.720 1.375 ;
        RECT  3.960 1.145 4.620 1.375 ;
        RECT  3.860 0.985 3.960 1.375 ;
        RECT  3.185 1.145 3.860 1.375 ;
        RECT  3.115 0.860 3.185 1.375 ;
        RECT  2.440 1.145 3.115 1.375 ;
        RECT  2.340 0.985 2.440 1.375 ;
        RECT  1.670 1.145 2.340 1.375 ;
        RECT  1.600 0.815 1.670 1.375 ;
        RECT  0.920 1.145 1.600 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.120 1.145 0.800 1.375 ;
        RECT  0.050 0.720 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.960 0.210 6.055 0.370 ;
        RECT  5.880 0.210 5.960 0.915 ;
        RECT  5.020 0.210 5.880 0.280 ;
        RECT  5.770 0.845 5.880 0.915 ;
        RECT  5.020 0.845 5.110 0.915 ;
        RECT  4.950 0.210 5.020 0.915 ;
        RECT  4.390 0.210 4.950 0.370 ;
        RECT  4.310 0.210 4.390 0.915 ;
        RECT  1.980 0.210 2.810 0.280 ;
        RECT  2.710 0.835 2.810 0.915 ;
        RECT  1.980 0.835 2.070 0.915 ;
        RECT  1.900 0.210 1.980 0.915 ;
        RECT  1.355 0.210 1.900 0.370 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.190 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        RECT  5.735 0.520 5.760 0.665 ;
        RECT  5.645 0.350 5.735 0.665 ;
        RECT  5.265 0.350 5.645 0.420 ;
        RECT  5.190 0.350 5.265 0.630 ;
        RECT  5.090 0.510 5.190 0.630 ;
        RECT  4.135 0.495 4.235 0.640 ;
        RECT  4.065 0.350 4.135 0.640 ;
        RECT  3.755 0.350 4.065 0.420 ;
        RECT  3.685 0.350 3.755 0.665 ;
        RECT  3.610 0.495 3.685 0.665 ;
        RECT  1.100 0.495 1.165 0.640 ;
        RECT  1.025 0.355 1.100 0.640 ;
        RECT  0.650 0.355 1.025 0.425 ;
        RECT  0.565 0.355 0.650 0.640 ;
        RECT  0.540 0.495 0.565 0.640 ;
        RECT  3.605 0.210 4.310 0.280 ;
        RECT  4.230 0.835 4.310 0.915 ;
        RECT  2.890 0.210 3.255 0.350 ;
        RECT  2.810 0.210 2.890 0.915 ;
    END
END NR2D16BWP40

MACRO NR2D1BWP40
    CLASS CORE ;
    FOREIGN NR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.104250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.325 0.525 1.045 ;
        RECT  0.325 0.325 0.455 0.395 ;
        RECT  0.435 0.915 0.455 1.045 ;
        RECT  0.235 0.210 0.325 0.395 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.510 -0.115 0.560 0.115 ;
        RECT  0.430 -0.115 0.510 0.255 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.145 0.560 1.375 ;
        RECT  0.050 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
END NR2D1BWP40

MACRO NR2D20BWP40
    CLASS CORE ;
    FOREIGN NR2D20BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.671600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.480 0.210 7.610 0.395 ;
        RECT  7.410 0.210 7.480 0.915 ;
        RECT  6.540 0.210 7.410 0.285 ;
        RECT  7.310 0.845 7.410 0.915 ;
        RECT  6.540 0.845 6.650 0.915 ;
        RECT  6.460 0.210 6.540 0.915 ;
        RECT  5.930 0.210 6.460 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.020 0.210 5.850 0.280 ;
        RECT  5.770 0.845 5.850 0.915 ;
        RECT  5.020 0.845 5.110 0.915 ;
        RECT  4.950 0.210 5.020 0.915 ;
        RECT  4.390 0.210 4.950 0.370 ;
        RECT  4.310 0.210 4.390 0.915 ;
        RECT  3.535 0.210 4.310 0.280 ;
        RECT  4.230 0.835 4.310 0.915 ;
        RECT  3.535 0.835 3.605 0.915 ;
        RECT  3.450 0.210 3.535 0.915 ;
        RECT  3.325 0.210 3.450 0.625 ;
        RECT  2.890 0.210 3.325 0.350 ;
        RECT  2.810 0.210 2.890 0.915 ;
        RECT  1.980 0.210 2.810 0.280 ;
        RECT  2.710 0.835 2.810 0.915 ;
        RECT  1.980 0.835 2.070 0.915 ;
        RECT  1.900 0.210 1.980 0.915 ;
        RECT  1.355 0.210 1.900 0.370 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.190 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.572800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 0.495 7.755 0.625 ;
        RECT  7.570 0.495 7.640 1.065 ;
        RECT  7.215 0.995 7.570 1.065 ;
        RECT  7.145 0.845 7.215 1.065 ;
        RECT  7.010 0.845 7.145 0.915 ;
        RECT  6.895 0.495 7.010 0.915 ;
        RECT  6.825 0.845 6.895 0.915 ;
        RECT  6.745 0.845 6.825 1.065 ;
        RECT  6.390 0.995 6.745 1.065 ;
        RECT  6.310 0.495 6.390 1.065 ;
        RECT  6.090 0.495 6.310 0.625 ;
        RECT  6.010 0.495 6.090 1.065 ;
        RECT  5.675 0.995 6.010 1.065 ;
        RECT  5.605 0.845 5.675 1.065 ;
        RECT  5.480 0.845 5.605 0.915 ;
        RECT  5.355 0.495 5.480 0.915 ;
        RECT  5.285 0.845 5.355 0.915 ;
        RECT  5.205 0.845 5.285 1.065 ;
        RECT  4.870 0.995 5.205 1.065 ;
        RECT  4.795 0.495 4.870 1.065 ;
        RECT  4.540 0.495 4.795 0.625 ;
        RECT  4.470 0.495 4.540 1.055 ;
        RECT  4.130 0.985 4.470 1.055 ;
        RECT  4.050 0.845 4.130 1.055 ;
        RECT  3.985 0.845 4.050 0.915 ;
        RECT  3.885 0.525 3.985 0.915 ;
        RECT  3.770 0.845 3.885 0.915 ;
        RECT  3.675 0.845 3.770 1.065 ;
        RECT  3.330 0.995 3.675 1.065 ;
        RECT  3.255 0.710 3.330 1.065 ;
        RECT  3.195 0.710 3.255 0.780 ;
        RECT  3.115 0.495 3.195 0.780 ;
        RECT  3.045 0.710 3.115 0.780 ;
        RECT  2.975 0.710 3.045 1.055 ;
        RECT  2.625 0.985 2.975 1.055 ;
        RECT  2.530 0.845 2.625 1.055 ;
        RECT  2.385 0.845 2.530 0.915 ;
        RECT  2.275 0.495 2.385 0.915 ;
        RECT  2.250 0.845 2.275 0.915 ;
        RECT  2.170 0.845 2.250 1.055 ;
        RECT  1.830 0.985 2.170 1.055 ;
        RECT  1.760 0.495 1.830 1.055 ;
        RECT  1.515 0.495 1.760 0.665 ;
        RECT  1.435 0.495 1.515 1.065 ;
        RECT  1.095 0.995 1.435 1.065 ;
        RECT  1.015 0.845 1.095 1.065 ;
        RECT  0.945 0.845 1.015 0.915 ;
        RECT  0.735 0.495 0.945 0.915 ;
        RECT  0.695 0.845 0.735 0.915 ;
        RECT  0.625 0.845 0.695 1.065 ;
        RECT  0.270 0.995 0.625 1.065 ;
        RECT  0.190 0.495 0.270 1.065 ;
        RECT  0.085 0.495 0.190 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.624000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.495 2.740 0.625 ;
        RECT  2.555 0.350 2.625 0.625 ;
        RECT  2.205 0.350 2.555 0.420 ;
        RECT  2.065 0.350 2.205 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 -0.115 7.840 0.115 ;
        RECT  7.700 -0.115 7.800 0.410 ;
        RECT  7.430 -0.115 7.700 0.115 ;
        RECT  7.310 -0.115 7.430 0.140 ;
        RECT  7.045 -0.115 7.310 0.115 ;
        RECT  6.905 -0.115 7.045 0.140 ;
        RECT  6.650 -0.115 6.905 0.115 ;
        RECT  6.530 -0.115 6.650 0.140 ;
        RECT  6.275 -0.115 6.530 0.115 ;
        RECT  6.145 -0.115 6.275 0.140 ;
        RECT  5.890 -0.115 6.145 0.115 ;
        RECT  5.770 -0.115 5.890 0.140 ;
        RECT  5.500 -0.115 5.770 0.115 ;
        RECT  5.380 -0.115 5.500 0.140 ;
        RECT  5.110 -0.115 5.380 0.115 ;
        RECT  4.990 -0.115 5.110 0.140 ;
        RECT  4.730 -0.115 4.990 0.115 ;
        RECT  4.610 -0.115 4.730 0.140 ;
        RECT  4.350 -0.115 4.610 0.115 ;
        RECT  4.230 -0.115 4.350 0.140 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.140 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.140 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.140 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.140 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.140 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.140 ;
        RECT  1.695 -0.115 1.950 0.115 ;
        RECT  1.565 -0.115 1.695 0.140 ;
        RECT  1.310 -0.115 1.565 0.115 ;
        RECT  1.190 -0.115 1.310 0.140 ;
        RECT  0.920 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.920 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.785 1.145 7.840 1.375 ;
        RECT  7.715 0.720 7.785 1.375 ;
        RECT  7.040 1.145 7.715 1.375 ;
        RECT  6.920 0.985 7.040 1.375 ;
        RECT  6.240 1.145 6.920 1.375 ;
        RECT  6.170 0.805 6.240 1.375 ;
        RECT  5.500 1.145 6.170 1.375 ;
        RECT  5.380 0.985 5.500 1.375 ;
        RECT  4.720 1.145 5.380 1.375 ;
        RECT  4.620 0.845 4.720 1.375 ;
        RECT  3.960 1.145 4.620 1.375 ;
        RECT  3.860 0.985 3.960 1.375 ;
        RECT  3.185 1.145 3.860 1.375 ;
        RECT  3.115 0.860 3.185 1.375 ;
        RECT  2.440 1.145 3.115 1.375 ;
        RECT  2.340 0.985 2.440 1.375 ;
        RECT  1.670 1.145 2.340 1.375 ;
        RECT  1.600 0.815 1.670 1.375 ;
        RECT  0.920 1.145 1.600 1.375 ;
        RECT  0.800 0.985 0.920 1.375 ;
        RECT  0.120 1.145 0.800 1.375 ;
        RECT  0.050 0.720 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.480 0.210 7.610 0.395 ;
        RECT  7.410 0.210 7.480 0.915 ;
        RECT  6.540 0.210 7.410 0.285 ;
        RECT  7.310 0.845 7.410 0.915 ;
        RECT  6.540 0.845 6.650 0.915 ;
        RECT  6.460 0.210 6.540 0.915 ;
        RECT  5.930 0.210 6.460 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.020 0.210 5.850 0.280 ;
        RECT  5.770 0.845 5.850 0.915 ;
        RECT  5.020 0.845 5.110 0.915 ;
        RECT  4.950 0.210 5.020 0.915 ;
        RECT  4.390 0.210 4.950 0.370 ;
        RECT  4.310 0.210 4.390 0.915 ;
        RECT  3.605 0.210 4.310 0.280 ;
        RECT  4.230 0.835 4.310 0.915 ;
        RECT  2.890 0.210 3.255 0.350 ;
        RECT  2.810 0.210 2.890 0.915 ;
        RECT  1.980 0.210 2.810 0.280 ;
        RECT  2.710 0.835 2.810 0.915 ;
        RECT  1.980 0.835 2.070 0.915 ;
        RECT  1.900 0.210 1.980 0.915 ;
        RECT  1.355 0.210 1.900 0.370 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.190 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        RECT  7.215 0.495 7.285 0.640 ;
        RECT  7.140 0.355 7.215 0.640 ;
        RECT  6.775 0.355 7.140 0.425 ;
        RECT  6.685 0.355 6.775 0.640 ;
        RECT  6.660 0.495 6.685 0.640 ;
        RECT  5.735 0.520 5.760 0.665 ;
        RECT  5.645 0.350 5.735 0.665 ;
        RECT  5.265 0.350 5.645 0.420 ;
        RECT  5.190 0.350 5.265 0.630 ;
        RECT  5.090 0.510 5.190 0.630 ;
        RECT  1.025 0.355 1.100 0.640 ;
        RECT  0.650 0.355 1.025 0.425 ;
        RECT  0.565 0.355 0.650 0.640 ;
        RECT  0.540 0.495 0.565 0.640 ;
        RECT  4.135 0.495 4.235 0.640 ;
        RECT  4.065 0.350 4.135 0.640 ;
        RECT  3.755 0.350 4.065 0.420 ;
        RECT  3.685 0.350 3.755 0.665 ;
        RECT  3.610 0.495 3.685 0.665 ;
        RECT  1.100 0.495 1.165 0.640 ;
    END
END NR2D20BWP40

MACRO NR2D24BWP40
    CLASS CORE ;
    FOREIGN NR2D24BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 2.007900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.010 0.210 9.145 0.395 ;
        RECT  8.940 0.210 9.010 0.915 ;
        RECT  8.080 0.210 8.940 0.285 ;
        RECT  8.850 0.845 8.940 0.915 ;
        RECT  8.080 0.845 8.190 0.915 ;
        RECT  8.000 0.210 8.080 0.915 ;
        RECT  7.470 0.210 8.000 0.370 ;
        RECT  7.390 0.210 7.470 0.915 ;
        RECT  6.560 0.210 7.390 0.280 ;
        RECT  7.310 0.845 7.390 0.915 ;
        RECT  6.560 0.845 6.650 0.915 ;
        RECT  6.490 0.210 6.560 0.915 ;
        RECT  5.930 0.210 6.490 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.075 0.210 5.850 0.280 ;
        RECT  5.770 0.835 5.850 0.915 ;
        RECT  5.075 0.835 5.145 0.915 ;
        RECT  4.990 0.210 5.075 0.915 ;
        RECT  4.865 0.210 4.990 0.625 ;
        RECT  4.430 0.210 4.865 0.350 ;
        RECT  4.350 0.210 4.430 0.915 ;
        RECT  3.520 0.210 4.350 0.280 ;
        RECT  4.250 0.835 4.350 0.915 ;
        RECT  3.520 0.835 3.610 0.915 ;
        RECT  3.440 0.210 3.520 0.915 ;
        RECT  2.895 0.210 3.440 0.370 ;
        RECT  2.825 0.210 2.895 0.915 ;
        RECT  1.960 0.210 2.825 0.285 ;
        RECT  2.730 0.845 2.825 0.915 ;
        RECT  1.960 0.845 2.070 0.915 ;
        RECT  1.880 0.210 1.960 0.915 ;
        RECT  1.355 0.210 1.880 0.375 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.170 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.682800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.170 0.495 9.285 0.625 ;
        RECT  9.100 0.495 9.170 1.065 ;
        RECT  8.755 0.995 9.100 1.065 ;
        RECT  8.685 0.845 8.755 1.065 ;
        RECT  8.550 0.845 8.685 0.915 ;
        RECT  8.435 0.495 8.550 0.915 ;
        RECT  8.365 0.845 8.435 0.915 ;
        RECT  8.285 0.845 8.365 1.065 ;
        RECT  7.930 0.995 8.285 1.065 ;
        RECT  7.850 0.495 7.930 1.065 ;
        RECT  7.630 0.495 7.850 0.625 ;
        RECT  7.550 0.495 7.630 1.065 ;
        RECT  7.215 0.995 7.550 1.065 ;
        RECT  7.145 0.845 7.215 1.065 ;
        RECT  7.020 0.845 7.145 0.915 ;
        RECT  6.895 0.495 7.020 0.915 ;
        RECT  6.825 0.845 6.895 0.915 ;
        RECT  6.745 0.845 6.825 1.065 ;
        RECT  6.410 0.995 6.745 1.065 ;
        RECT  6.335 0.495 6.410 1.065 ;
        RECT  6.080 0.495 6.335 0.625 ;
        RECT  6.010 0.495 6.080 1.055 ;
        RECT  5.670 0.985 6.010 1.055 ;
        RECT  5.590 0.845 5.670 1.055 ;
        RECT  5.525 0.845 5.590 0.915 ;
        RECT  5.425 0.525 5.525 0.915 ;
        RECT  5.310 0.845 5.425 0.915 ;
        RECT  5.215 0.845 5.310 1.065 ;
        RECT  4.870 0.995 5.215 1.065 ;
        RECT  4.795 0.710 4.870 1.065 ;
        RECT  4.735 0.710 4.795 0.780 ;
        RECT  4.655 0.495 4.735 0.780 ;
        RECT  4.585 0.710 4.655 0.780 ;
        RECT  4.515 0.710 4.585 1.055 ;
        RECT  4.165 0.985 4.515 1.055 ;
        RECT  4.070 0.845 4.165 1.055 ;
        RECT  3.925 0.845 4.070 0.915 ;
        RECT  3.815 0.495 3.925 0.915 ;
        RECT  3.790 0.845 3.815 0.915 ;
        RECT  3.710 0.845 3.790 1.055 ;
        RECT  3.370 0.985 3.710 1.055 ;
        RECT  3.300 0.495 3.370 1.055 ;
        RECT  3.055 0.495 3.300 0.665 ;
        RECT  2.975 0.495 3.055 1.065 ;
        RECT  2.635 0.995 2.975 1.065 ;
        RECT  2.555 0.845 2.635 1.065 ;
        RECT  2.485 0.845 2.555 0.915 ;
        RECT  2.275 0.495 2.485 0.915 ;
        RECT  2.235 0.845 2.275 0.915 ;
        RECT  2.165 0.845 2.235 1.065 ;
        RECT  1.810 0.995 2.165 1.065 ;
        RECT  1.730 0.495 1.810 1.065 ;
        RECT  1.515 0.495 1.730 0.625 ;
        RECT  1.430 0.495 1.515 1.065 ;
        RECT  1.085 0.995 1.430 1.065 ;
        RECT  1.015 0.845 1.085 1.065 ;
        RECT  0.905 0.845 1.015 0.915 ;
        RECT  0.805 0.495 0.905 0.915 ;
        RECT  0.695 0.845 0.805 0.915 ;
        RECT  0.625 0.845 0.695 1.065 ;
        RECT  0.270 0.995 0.625 1.065 ;
        RECT  0.190 0.495 0.270 1.065 ;
        RECT  0.075 0.495 0.190 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.748800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.280 0.625 ;
        RECT  4.095 0.350 4.165 0.625 ;
        RECT  3.745 0.350 4.095 0.420 ;
        RECT  3.605 0.350 3.745 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.340 -0.115 9.380 0.115 ;
        RECT  9.240 -0.115 9.340 0.410 ;
        RECT  8.970 -0.115 9.240 0.115 ;
        RECT  8.850 -0.115 8.970 0.140 ;
        RECT  8.585 -0.115 8.850 0.115 ;
        RECT  8.445 -0.115 8.585 0.140 ;
        RECT  8.190 -0.115 8.445 0.115 ;
        RECT  8.070 -0.115 8.190 0.140 ;
        RECT  7.815 -0.115 8.070 0.115 ;
        RECT  7.685 -0.115 7.815 0.140 ;
        RECT  7.430 -0.115 7.685 0.115 ;
        RECT  7.310 -0.115 7.430 0.140 ;
        RECT  7.040 -0.115 7.310 0.115 ;
        RECT  6.920 -0.115 7.040 0.140 ;
        RECT  6.650 -0.115 6.920 0.115 ;
        RECT  6.530 -0.115 6.650 0.140 ;
        RECT  6.270 -0.115 6.530 0.115 ;
        RECT  6.150 -0.115 6.270 0.140 ;
        RECT  5.890 -0.115 6.150 0.115 ;
        RECT  5.770 -0.115 5.890 0.140 ;
        RECT  5.510 -0.115 5.770 0.115 ;
        RECT  5.390 -0.115 5.510 0.140 ;
        RECT  5.130 -0.115 5.390 0.115 ;
        RECT  5.010 -0.115 5.130 0.140 ;
        RECT  4.750 -0.115 5.010 0.115 ;
        RECT  4.630 -0.115 4.750 0.140 ;
        RECT  4.370 -0.115 4.630 0.115 ;
        RECT  4.250 -0.115 4.370 0.140 ;
        RECT  3.990 -0.115 4.250 0.115 ;
        RECT  3.870 -0.115 3.990 0.140 ;
        RECT  3.610 -0.115 3.870 0.115 ;
        RECT  3.490 -0.115 3.610 0.140 ;
        RECT  3.235 -0.115 3.490 0.115 ;
        RECT  3.105 -0.115 3.235 0.140 ;
        RECT  2.850 -0.115 3.105 0.115 ;
        RECT  2.730 -0.115 2.850 0.140 ;
        RECT  2.460 -0.115 2.730 0.115 ;
        RECT  2.330 -0.115 2.460 0.140 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.140 ;
        RECT  1.695 -0.115 1.950 0.115 ;
        RECT  1.560 -0.115 1.695 0.140 ;
        RECT  1.300 -0.115 1.560 0.115 ;
        RECT  1.180 -0.115 1.300 0.140 ;
        RECT  0.910 -0.115 1.180 0.115 ;
        RECT  0.785 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.785 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.325 1.145 9.380 1.375 ;
        RECT  9.255 0.720 9.325 1.375 ;
        RECT  8.580 1.145 9.255 1.375 ;
        RECT  8.460 0.985 8.580 1.375 ;
        RECT  7.780 1.145 8.460 1.375 ;
        RECT  7.710 0.805 7.780 1.375 ;
        RECT  7.040 1.145 7.710 1.375 ;
        RECT  6.920 0.985 7.040 1.375 ;
        RECT  6.260 1.145 6.920 1.375 ;
        RECT  6.160 0.845 6.260 1.375 ;
        RECT  5.500 1.145 6.160 1.375 ;
        RECT  5.400 0.985 5.500 1.375 ;
        RECT  4.725 1.145 5.400 1.375 ;
        RECT  4.655 0.860 4.725 1.375 ;
        RECT  3.980 1.145 4.655 1.375 ;
        RECT  3.880 0.985 3.980 1.375 ;
        RECT  3.210 1.145 3.880 1.375 ;
        RECT  3.140 0.815 3.210 1.375 ;
        RECT  2.460 1.145 3.140 1.375 ;
        RECT  2.340 0.985 2.460 1.375 ;
        RECT  1.660 1.145 2.340 1.375 ;
        RECT  1.590 0.800 1.660 1.375 ;
        RECT  0.910 1.145 1.590 1.375 ;
        RECT  0.790 0.985 0.910 1.375 ;
        RECT  0.120 1.145 0.790 1.375 ;
        RECT  0.050 0.720 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.010 0.210 9.145 0.395 ;
        RECT  8.940 0.210 9.010 0.915 ;
        RECT  8.080 0.210 8.940 0.285 ;
        RECT  8.850 0.845 8.940 0.915 ;
        RECT  8.080 0.845 8.190 0.915 ;
        RECT  8.000 0.210 8.080 0.915 ;
        RECT  7.470 0.210 8.000 0.370 ;
        RECT  7.390 0.210 7.470 0.915 ;
        RECT  6.560 0.210 7.390 0.280 ;
        RECT  7.310 0.845 7.390 0.915 ;
        RECT  6.560 0.845 6.650 0.915 ;
        RECT  6.490 0.210 6.560 0.915 ;
        RECT  5.930 0.210 6.490 0.370 ;
        RECT  5.850 0.210 5.930 0.915 ;
        RECT  5.145 0.210 5.850 0.280 ;
        RECT  5.770 0.835 5.850 0.915 ;
        RECT  4.430 0.210 4.795 0.350 ;
        RECT  4.350 0.210 4.430 0.915 ;
        RECT  3.520 0.210 4.350 0.280 ;
        RECT  4.250 0.835 4.350 0.915 ;
        RECT  3.520 0.835 3.610 0.915 ;
        RECT  3.440 0.210 3.520 0.915 ;
        RECT  2.895 0.210 3.440 0.370 ;
        RECT  2.825 0.210 2.895 0.915 ;
        RECT  1.960 0.210 2.825 0.285 ;
        RECT  2.730 0.845 2.825 0.915 ;
        RECT  1.960 0.845 2.070 0.915 ;
        RECT  1.880 0.210 1.960 0.915 ;
        RECT  1.355 0.210 1.880 0.375 ;
        RECT  1.285 0.210 1.355 0.915 ;
        RECT  0.420 0.210 1.285 0.285 ;
        RECT  1.170 0.845 1.285 0.915 ;
        RECT  0.420 0.845 0.530 0.915 ;
        RECT  0.340 0.210 0.420 0.915 ;
        RECT  0.245 0.210 0.340 0.375 ;
        RECT  8.755 0.495 8.825 0.640 ;
        RECT  8.680 0.355 8.755 0.640 ;
        RECT  8.315 0.355 8.680 0.425 ;
        RECT  8.225 0.355 8.315 0.640 ;
        RECT  8.200 0.495 8.225 0.640 ;
        RECT  7.275 0.520 7.300 0.665 ;
        RECT  7.185 0.350 7.275 0.665 ;
        RECT  6.805 0.350 7.185 0.420 ;
        RECT  6.730 0.350 6.805 0.630 ;
        RECT  6.630 0.510 6.730 0.630 ;
        RECT  5.675 0.495 5.775 0.640 ;
        RECT  5.605 0.350 5.675 0.640 ;
        RECT  5.295 0.350 5.605 0.420 ;
        RECT  5.225 0.350 5.295 0.665 ;
        RECT  5.150 0.495 5.225 0.665 ;
        RECT  2.640 0.495 2.705 0.640 ;
        RECT  2.565 0.355 2.640 0.640 ;
        RECT  2.190 0.355 2.565 0.425 ;
        RECT  2.105 0.355 2.190 0.640 ;
        RECT  2.080 0.495 2.105 0.640 ;
        RECT  1.085 0.495 1.155 0.640 ;
        RECT  1.010 0.355 1.085 0.640 ;
        RECT  0.655 0.355 1.010 0.425 ;
        RECT  0.565 0.355 0.655 0.640 ;
        RECT  0.540 0.495 0.565 0.640 ;
    END
END NR2D24BWP40

MACRO NR2D2BWP40
    CLASS CORE ;
    FOREIGN NR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.172500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.225 0.720 0.425 ;
        RECT  0.390 0.345 0.640 0.425 ;
        RECT  0.355 0.345 0.390 0.915 ;
        RECT  0.315 0.215 0.355 0.915 ;
        RECT  0.260 0.215 0.315 0.425 ;
        RECT  0.175 0.845 0.315 0.915 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 0.495 0.815 0.625 ;
        RECT  0.595 0.495 0.680 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.425 ;
        RECT  0.540 -0.115 0.830 0.115 ;
        RECT  0.440 -0.115 0.540 0.270 ;
        RECT  0.145 -0.115 0.440 0.115 ;
        RECT  0.075 -0.115 0.145 0.420 ;
        RECT  0.000 -0.115 0.075 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.145 0.980 1.375 ;
        RECT  0.630 0.985 0.730 1.375 ;
        RECT  0.000 1.145 0.630 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 0.755 0.910 1.005 ;
        RECT  0.530 0.845 0.830 0.915 ;
        RECT  0.460 0.845 0.530 1.055 ;
        RECT  0.035 0.985 0.460 1.055 ;
    END
END NR2D2BWP40

MACRO NR2D3BWP40
    CLASS CORE ;
    FOREIGN NR2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.290750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.185 1.130 0.425 ;
        RECT  0.720 0.355 1.030 0.425 ;
        RECT  0.620 0.185 0.720 0.425 ;
        RECT  0.525 0.355 0.620 0.425 ;
        RECT  0.455 0.355 0.525 0.905 ;
        RECT  0.330 0.355 0.455 0.425 ;
        RECT  0.140 0.835 0.455 0.905 ;
        RECT  0.230 0.185 0.330 0.425 ;
        RECT  0.035 0.835 0.140 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.495 1.110 0.625 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.385 0.640 ;
        RECT  0.145 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.420 ;
        RECT  0.920 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.920 0.270 ;
        RECT  0.520 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.520 0.270 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.420 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.725 1.360 1.375 ;
        RECT  0.920 1.145 1.260 1.375 ;
        RECT  0.820 0.985 0.920 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.030 0.835 1.130 1.075 ;
        RECT  0.695 0.835 1.030 0.905 ;
        RECT  0.625 0.835 0.695 1.050 ;
        RECT  0.220 0.980 0.625 1.050 ;
    END
END NR2D3BWP40

MACRO NR2D4BWP40
    CLASS CORE ;
    FOREIGN NR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.336300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.215 1.575 0.525 ;
        RECT  1.365 0.215 1.435 0.915 ;
        RECT  0.440 0.215 1.365 0.285 ;
        RECT  1.250 0.845 1.365 0.915 ;
        RECT  0.440 0.845 0.550 0.915 ;
        RECT  0.360 0.215 0.440 0.915 ;
        RECT  0.265 0.215 0.360 0.375 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.122800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.595 1.675 0.665 ;
        RECT  1.525 0.595 1.595 1.065 ;
        RECT  1.155 0.995 1.525 1.065 ;
        RECT  1.085 0.720 1.155 1.065 ;
        RECT  0.950 0.720 1.085 0.790 ;
        RECT  0.850 0.495 0.950 0.790 ;
        RECT  0.715 0.720 0.850 0.790 ;
        RECT  0.645 0.720 0.715 1.065 ;
        RECT  0.290 0.995 0.645 1.065 ;
        RECT  0.210 0.495 0.290 1.065 ;
        RECT  0.035 0.495 0.210 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.640 ;
        RECT  1.080 0.355 1.155 0.640 ;
        RECT  0.675 0.355 1.080 0.425 ;
        RECT  0.585 0.355 0.675 0.640 ;
        RECT  0.560 0.495 0.585 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 -0.115 1.820 0.115 ;
        RECT  1.680 -0.115 1.780 0.410 ;
        RECT  1.370 -0.115 1.680 0.115 ;
        RECT  1.250 -0.115 1.370 0.145 ;
        RECT  0.960 -0.115 1.250 0.115 ;
        RECT  0.840 -0.115 0.960 0.145 ;
        RECT  0.550 -0.115 0.840 0.115 ;
        RECT  0.430 -0.115 0.550 0.140 ;
        RECT  0.140 -0.115 0.430 0.115 ;
        RECT  0.040 -0.115 0.140 0.410 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.145 1.820 1.375 ;
        RECT  1.680 0.845 1.780 1.375 ;
        RECT  0.960 1.145 1.680 1.375 ;
        RECT  0.840 0.890 0.960 1.375 ;
        RECT  0.120 1.145 0.840 1.375 ;
        RECT  0.050 0.720 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.440 0.215 1.295 0.285 ;
        RECT  1.250 0.845 1.295 0.915 ;
        RECT  0.440 0.845 0.550 0.915 ;
        RECT  0.360 0.215 0.440 0.915 ;
        RECT  0.265 0.215 0.360 0.375 ;
    END
END NR2D4BWP40

MACRO NR2D6BWP40
    CLASS CORE ;
    FOREIGN NR2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.599500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.840 2.625 1.045 ;
        RECT  2.510 0.355 2.555 1.045 ;
        RECT  2.380 0.355 2.510 0.910 ;
        RECT  2.345 0.195 2.380 0.910 ;
        RECT  2.300 0.195 2.345 0.425 ;
        RECT  2.090 0.840 2.345 0.910 ;
        RECT  1.990 0.355 2.300 0.425 ;
        RECT  1.910 0.195 1.990 0.425 ;
        RECT  1.580 0.355 1.910 0.425 ;
        RECT  1.500 0.195 1.580 0.425 ;
        RECT  1.120 0.355 1.500 0.425 ;
        RECT  1.040 0.195 1.120 0.425 ;
        RECT  0.710 0.355 1.040 0.425 ;
        RECT  0.630 0.195 0.710 0.425 ;
        RECT  0.320 0.355 0.630 0.425 ;
        RECT  0.130 0.840 0.530 0.910 ;
        RECT  0.240 0.195 0.320 0.425 ;
        RECT  0.130 0.355 0.240 0.425 ;
        RECT  0.050 0.355 0.130 1.065 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 1.885 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.075 0.495 2.205 0.765 ;
        RECT  0.665 0.695 2.075 0.765 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.320 0.495 0.595 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.620 -0.115 2.660 0.115 ;
        RECT  2.520 -0.115 2.620 0.270 ;
        RECT  2.200 -0.115 2.520 0.115 ;
        RECT  2.100 -0.115 2.200 0.270 ;
        RECT  1.800 -0.115 2.100 0.115 ;
        RECT  1.700 -0.115 1.800 0.270 ;
        RECT  1.360 -0.115 1.700 0.115 ;
        RECT  1.260 -0.115 1.360 0.270 ;
        RECT  0.920 -0.115 1.260 0.115 ;
        RECT  0.820 -0.115 0.920 0.270 ;
        RECT  0.520 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.520 0.270 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.270 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.145 2.660 1.375 ;
        RECT  1.700 0.985 1.800 1.375 ;
        RECT  1.360 1.145 1.700 1.375 ;
        RECT  1.260 0.985 1.360 1.375 ;
        RECT  0.920 1.145 1.260 1.375 ;
        RECT  0.820 0.985 0.920 1.375 ;
        RECT  0.000 1.145 0.820 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.990 0.355 2.275 0.425 ;
        RECT  2.090 0.840 2.275 0.910 ;
        RECT  1.910 0.195 1.990 0.425 ;
        RECT  1.580 0.355 1.910 0.425 ;
        RECT  1.500 0.195 1.580 0.425 ;
        RECT  1.120 0.355 1.500 0.425 ;
        RECT  1.040 0.195 1.120 0.425 ;
        RECT  0.710 0.355 1.040 0.425 ;
        RECT  0.630 0.195 0.710 0.425 ;
        RECT  0.320 0.355 0.630 0.425 ;
        RECT  0.130 0.840 0.530 0.910 ;
        RECT  0.240 0.195 0.320 0.425 ;
        RECT  0.130 0.355 0.240 0.425 ;
        RECT  0.050 0.355 0.130 1.065 ;
        RECT  1.995 0.980 2.400 1.050 ;
        RECT  1.925 0.835 1.995 1.050 ;
        RECT  1.580 0.835 1.925 0.905 ;
        RECT  1.500 0.835 1.580 1.065 ;
        RECT  1.120 0.835 1.500 0.905 ;
        RECT  1.040 0.835 1.120 1.065 ;
        RECT  0.695 0.835 1.040 0.905 ;
        RECT  0.625 0.835 0.695 1.050 ;
        RECT  0.220 0.980 0.625 1.050 ;
    END
END NR2D6BWP40

MACRO NR2D8BWP40
    CLASS CORE ;
    FOREIGN NR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.220 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.666000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.210 2.975 0.370 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  1.995 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.995 0.825 2.065 0.905 ;
        RECT  1.910 0.210 1.995 0.905 ;
        RECT  1.785 0.210 1.910 0.625 ;
        RECT  1.350 0.210 1.785 0.350 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.236800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.000 0.495 3.110 0.635 ;
        RECT  2.930 0.495 3.000 1.055 ;
        RECT  2.590 0.985 2.930 1.055 ;
        RECT  2.510 0.845 2.590 1.055 ;
        RECT  2.445 0.845 2.510 0.915 ;
        RECT  2.345 0.495 2.445 0.915 ;
        RECT  2.230 0.845 2.345 0.915 ;
        RECT  2.135 0.845 2.230 1.055 ;
        RECT  1.790 0.985 2.135 1.055 ;
        RECT  1.715 0.710 1.790 1.055 ;
        RECT  1.655 0.710 1.715 0.780 ;
        RECT  1.575 0.495 1.655 0.780 ;
        RECT  1.505 0.710 1.575 0.780 ;
        RECT  1.435 0.710 1.505 1.055 ;
        RECT  1.085 0.985 1.435 1.055 ;
        RECT  0.990 0.845 1.085 1.055 ;
        RECT  0.845 0.845 0.990 0.915 ;
        RECT  0.735 0.495 0.845 0.915 ;
        RECT  0.710 0.845 0.735 0.915 ;
        RECT  0.630 0.845 0.710 1.055 ;
        RECT  0.290 0.985 0.630 1.055 ;
        RECT  0.220 0.495 0.290 1.055 ;
        RECT  0.150 0.495 0.220 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.249600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.200 0.625 ;
        RECT  1.015 0.350 1.085 0.625 ;
        RECT  0.665 0.350 1.015 0.420 ;
        RECT  0.525 0.350 0.665 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.170 -0.115 3.220 0.115 ;
        RECT  3.090 -0.115 3.170 0.420 ;
        RECT  2.810 -0.115 3.090 0.115 ;
        RECT  2.690 -0.115 2.810 0.140 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.140 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.140 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.140 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.140 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.420 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.145 3.220 1.375 ;
        RECT  3.080 0.730 3.180 1.375 ;
        RECT  2.420 1.145 3.080 1.375 ;
        RECT  2.320 0.985 2.420 1.375 ;
        RECT  1.645 1.145 2.320 1.375 ;
        RECT  1.575 0.860 1.645 1.375 ;
        RECT  0.900 1.145 1.575 1.375 ;
        RECT  0.800 0.985 0.900 1.375 ;
        RECT  0.140 1.145 0.800 1.375 ;
        RECT  0.040 0.725 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 0.210 2.975 0.370 ;
        RECT  2.770 0.210 2.850 0.915 ;
        RECT  2.065 0.210 2.770 0.280 ;
        RECT  2.690 0.835 2.770 0.915 ;
        RECT  1.350 0.210 1.715 0.350 ;
        RECT  1.270 0.210 1.350 0.915 ;
        RECT  0.440 0.210 1.270 0.280 ;
        RECT  1.170 0.835 1.270 0.915 ;
        RECT  0.440 0.835 0.530 0.915 ;
        RECT  0.360 0.210 0.440 0.915 ;
        RECT  0.245 0.210 0.360 0.370 ;
        RECT  2.595 0.495 2.695 0.640 ;
        RECT  2.525 0.350 2.595 0.640 ;
        RECT  2.215 0.350 2.525 0.420 ;
        RECT  2.145 0.350 2.215 0.665 ;
        RECT  2.070 0.495 2.145 0.665 ;
    END
END NR2D8BWP40

MACRO NR3D0BWP40
    CLASS CORE ;
    FOREIGN NR3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.072250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.915 ;
        RECT  0.525 0.345 0.735 0.415 ;
        RECT  0.545 0.845 0.735 0.915 ;
        RECT  0.455 0.845 0.545 1.045 ;
        RECT  0.455 0.215 0.525 0.415 ;
        RECT  0.140 0.345 0.455 0.415 ;
        RECT  0.130 0.970 0.455 1.045 ;
        RECT  0.035 0.205 0.140 0.415 ;
        RECT  0.035 0.915 0.130 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.825 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.840 0.115 ;
        RECT  0.640 -0.115 0.760 0.235 ;
        RECT  0.350 -0.115 0.640 0.115 ;
        RECT  0.230 -0.115 0.350 0.215 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.840 1.375 ;
        RECT  0.640 0.985 0.760 1.375 ;
        RECT  0.000 1.145 0.640 1.375 ;
        END
    END VDD
END NR3D0BWP40

MACRO NR3D12BWP40
    CLASS CORE ;
    FOREIGN NR3D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.350000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.835 7.020 0.905 ;
        RECT  5.915 0.305 7.010 0.415 ;
        RECT  5.705 0.305 5.915 0.905 ;
        RECT  0.250 0.305 5.705 0.415 ;
        RECT  5.000 0.835 5.705 0.905 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 0.495 2.185 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.495 4.195 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.384000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.905 0.495 5.625 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.225 -0.115 7.280 0.115 ;
        RECT  7.155 -0.115 7.225 0.425 ;
        RECT  6.830 -0.115 7.155 0.115 ;
        RECT  6.710 -0.115 6.830 0.235 ;
        RECT  6.450 -0.115 6.710 0.115 ;
        RECT  6.330 -0.115 6.450 0.235 ;
        RECT  6.070 -0.115 6.330 0.115 ;
        RECT  5.950 -0.115 6.070 0.235 ;
        RECT  5.690 -0.115 5.950 0.115 ;
        RECT  5.570 -0.115 5.690 0.235 ;
        RECT  5.310 -0.115 5.570 0.115 ;
        RECT  5.190 -0.115 5.310 0.235 ;
        RECT  4.930 -0.115 5.190 0.115 ;
        RECT  4.810 -0.115 4.930 0.235 ;
        RECT  4.730 -0.115 4.810 0.115 ;
        RECT  4.610 -0.115 4.730 0.235 ;
        RECT  4.350 -0.115 4.610 0.115 ;
        RECT  4.230 -0.115 4.350 0.235 ;
        RECT  3.970 -0.115 4.230 0.115 ;
        RECT  3.850 -0.115 3.970 0.235 ;
        RECT  3.590 -0.115 3.850 0.115 ;
        RECT  3.470 -0.115 3.590 0.235 ;
        RECT  3.210 -0.115 3.470 0.115 ;
        RECT  3.090 -0.115 3.210 0.235 ;
        RECT  2.830 -0.115 3.090 0.115 ;
        RECT  2.710 -0.115 2.830 0.235 ;
        RECT  2.450 -0.115 2.710 0.115 ;
        RECT  2.330 -0.115 2.450 0.235 ;
        RECT  2.070 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.070 0.235 ;
        RECT  1.690 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.690 0.235 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.235 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.235 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.550 0.235 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.145 7.280 1.375 ;
        RECT  2.160 0.975 2.240 1.375 ;
        RECT  1.860 1.145 2.160 1.375 ;
        RECT  1.780 0.975 1.860 1.375 ;
        RECT  1.480 1.145 1.780 1.375 ;
        RECT  1.400 0.975 1.480 1.375 ;
        RECT  1.100 1.145 1.400 1.375 ;
        RECT  1.020 0.975 1.100 1.375 ;
        RECT  0.720 1.145 1.020 1.375 ;
        RECT  0.640 0.975 0.720 1.375 ;
        RECT  0.340 1.145 0.640 1.375 ;
        RECT  0.260 0.975 0.340 1.375 ;
        RECT  0.000 1.145 0.260 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.985 0.835 7.020 0.905 ;
        RECT  5.985 0.305 7.010 0.415 ;
        RECT  0.250 0.305 5.635 0.415 ;
        RECT  5.000 0.835 5.635 0.905 ;
        RECT  7.155 0.785 7.225 1.045 ;
        RECT  2.520 0.975 7.155 1.045 ;
        RECT  6.050 0.545 6.715 0.615 ;
        RECT  2.425 0.835 4.730 0.905 ;
        RECT  2.355 0.835 2.425 1.075 ;
        RECT  2.045 0.835 2.355 0.905 ;
        RECT  1.975 0.835 2.045 1.075 ;
        RECT  1.665 0.835 1.975 0.905 ;
        RECT  1.595 0.835 1.665 1.075 ;
        RECT  1.285 0.835 1.595 0.905 ;
        RECT  1.215 0.835 1.285 1.075 ;
        RECT  0.905 0.835 1.215 0.905 ;
        RECT  0.835 0.835 0.905 1.075 ;
        RECT  0.525 0.835 0.835 0.905 ;
        RECT  0.455 0.835 0.525 1.075 ;
        RECT  0.140 0.835 0.455 0.905 ;
        RECT  0.040 0.835 0.140 1.075 ;
    END
END NR3D12BWP40

MACRO NR3D1BWP40
    CLASS CORE ;
    FOREIGN NR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.144500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.915 ;
        RECT  0.565 0.355 0.735 0.425 ;
        RECT  0.545 0.845 0.735 0.915 ;
        RECT  0.495 0.285 0.565 0.425 ;
        RECT  0.455 0.845 0.545 1.045 ;
        RECT  0.140 0.285 0.495 0.355 ;
        RECT  0.130 0.970 0.455 1.045 ;
        RECT  0.035 0.215 0.140 0.355 ;
        RECT  0.035 0.910 0.130 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.425 0.385 0.825 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.840 0.115 ;
        RECT  0.640 -0.115 0.760 0.285 ;
        RECT  0.350 -0.115 0.640 0.115 ;
        RECT  0.230 -0.115 0.350 0.215 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.145 0.840 1.375 ;
        RECT  0.640 0.985 0.760 1.375 ;
        RECT  0.000 1.145 0.640 1.375 ;
        END
    END VDD
END NR3D1BWP40

MACRO NR3D2BWP40
    CLASS CORE ;
    FOREIGN NR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.262200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 0.210 1.365 0.970 ;
        RECT  0.165 0.210 1.280 0.280 ;
        RECT  0.595 0.900 1.280 0.970 ;
        RECT  0.035 0.210 0.165 0.420 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.475 1.195 0.810 ;
        RECT  0.245 0.740 1.125 0.810 ;
        RECT  0.175 0.495 0.245 0.810 ;
        RECT  0.035 0.495 0.175 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.545 1.040 0.615 ;
        RECT  0.875 0.350 0.945 0.615 ;
        RECT  0.525 0.350 0.875 0.420 ;
        RECT  0.455 0.350 0.525 0.625 ;
        RECT  0.315 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.155 -0.115 1.400 0.115 ;
        RECT  1.025 -0.115 1.155 0.140 ;
        RECT  0.760 -0.115 1.025 0.115 ;
        RECT  0.640 -0.115 0.760 0.140 ;
        RECT  0.370 -0.115 0.640 0.115 ;
        RECT  0.250 -0.115 0.370 0.140 ;
        RECT  0.000 -0.115 0.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.145 1.400 1.375 ;
        RECT  1.230 1.040 1.350 1.375 ;
        RECT  0.140 1.145 1.230 1.375 ;
        RECT  0.070 0.880 0.140 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
END NR3D2BWP40

MACRO NR3D3BWP40
    CLASS CORE ;
    FOREIGN NR3D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.385500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.185 1.705 0.415 ;
        RECT  1.290 0.325 1.610 0.415 ;
        RECT  1.210 0.185 1.290 0.415 ;
        RECT  0.910 0.325 1.210 0.415 ;
        RECT  0.830 0.185 0.910 0.415 ;
        RECT  0.595 0.325 0.830 0.415 ;
        RECT  0.530 0.325 0.595 0.915 ;
        RECT  0.450 0.185 0.530 0.915 ;
        RECT  0.385 0.325 0.450 0.915 ;
        RECT  0.130 0.325 0.385 0.415 ;
        RECT  0.130 0.845 0.385 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.495 1.745 0.625 ;
        RECT  1.410 0.495 1.515 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.495 1.155 0.625 ;
        RECT  0.735 0.495 0.815 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.310 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.830 -0.115 1.910 0.425 ;
        RECT  1.510 -0.115 1.830 0.115 ;
        RECT  1.390 -0.115 1.510 0.250 ;
        RECT  1.120 -0.115 1.390 0.115 ;
        RECT  1.000 -0.115 1.120 0.250 ;
        RECT  0.740 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.740 0.250 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.250 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 1.960 1.375 ;
        RECT  1.830 0.685 1.910 1.375 ;
        RECT  1.510 1.145 1.830 1.375 ;
        RECT  1.390 0.985 1.510 1.375 ;
        RECT  0.000 1.145 1.390 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.610 0.185 1.705 0.415 ;
        RECT  1.290 0.325 1.610 0.415 ;
        RECT  1.210 0.185 1.290 0.415 ;
        RECT  0.910 0.325 1.210 0.415 ;
        RECT  0.830 0.185 0.910 0.415 ;
        RECT  0.665 0.325 0.830 0.415 ;
        RECT  0.130 0.325 0.315 0.415 ;
        RECT  0.130 0.845 0.305 0.915 ;
        RECT  0.050 0.185 0.130 0.415 ;
        RECT  0.050 0.845 0.130 1.045 ;
        RECT  1.590 0.845 1.710 1.050 ;
        RECT  1.290 0.845 1.590 0.915 ;
        RECT  1.210 0.845 1.290 1.075 ;
        RECT  0.780 0.845 1.210 0.915 ;
        RECT  0.240 0.985 1.120 1.055 ;
    END
END NR3D3BWP40

MACRO NR3D4BWP40
    CLASS CORE ;
    FOREIGN NR3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.514975 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.215 2.625 0.790 ;
        RECT  2.535 0.215 2.555 0.970 ;
        RECT  2.530 0.215 2.535 0.495 ;
        RECT  2.415 0.720 2.535 0.970 ;
        RECT  0.130 0.215 2.530 0.285 ;
        RECT  2.345 0.720 2.415 1.055 ;
        RECT  0.605 0.985 2.345 1.055 ;
        RECT  0.035 0.215 0.130 0.345 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.123200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.355 2.455 0.640 ;
        RECT  1.365 0.355 2.380 0.425 ;
        RECT  1.265 0.355 1.365 0.630 ;
        RECT  0.270 0.355 1.265 0.425 ;
        RECT  0.200 0.355 0.270 0.625 ;
        RECT  0.035 0.495 0.200 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.116200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.230 0.495 2.290 0.620 ;
        RECT  2.120 0.495 2.230 0.915 ;
        RECT  1.725 0.845 2.120 0.915 ;
        RECT  1.590 0.635 1.725 0.915 ;
        RECT  1.045 0.845 1.590 0.915 ;
        RECT  0.915 0.635 1.045 0.915 ;
        RECT  0.525 0.775 0.915 0.915 ;
        RECT  0.435 0.495 0.525 0.915 ;
        RECT  0.370 0.495 0.435 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.117800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.795 0.495 2.020 0.625 ;
        RECT  1.520 0.495 1.795 0.565 ;
        RECT  1.435 0.495 1.520 0.775 ;
        RECT  1.185 0.705 1.435 0.775 ;
        RECT  1.115 0.495 1.185 0.775 ;
        RECT  0.845 0.495 1.115 0.565 ;
        RECT  0.595 0.495 0.845 0.685 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 -0.115 2.660 0.115 ;
        RECT  2.290 -0.115 2.410 0.145 ;
        RECT  2.000 -0.115 2.290 0.115 ;
        RECT  1.880 -0.115 2.000 0.145 ;
        RECT  1.620 -0.115 1.880 0.115 ;
        RECT  1.500 -0.115 1.620 0.145 ;
        RECT  1.180 -0.115 1.500 0.115 ;
        RECT  1.040 -0.115 1.180 0.145 ;
        RECT  0.760 -0.115 1.040 0.115 ;
        RECT  0.640 -0.115 0.760 0.145 ;
        RECT  0.355 -0.115 0.640 0.115 ;
        RECT  0.225 -0.115 0.355 0.145 ;
        RECT  0.000 -0.115 0.225 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.490 1.045 2.610 1.375 ;
        RECT  1.395 1.145 2.490 1.375 ;
        RECT  1.275 1.125 1.395 1.375 ;
        RECT  0.125 1.145 1.275 1.375 ;
        RECT  0.055 0.710 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.215 2.275 0.285 ;
        RECT  0.605 0.985 2.275 1.055 ;
        RECT  0.035 0.215 0.130 0.345 ;
    END
END NR3D4BWP40

MACRO NR3D6BWP40
    CLASS CORE ;
    FOREIGN NR3D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.675000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.785 3.560 0.905 ;
        RECT  3.325 0.315 3.535 0.905 ;
        RECT  2.660 0.315 3.325 0.425 ;
        RECT  2.680 0.775 3.325 0.905 ;
        RECT  2.265 0.335 2.660 0.425 ;
        RECT  0.230 0.315 2.265 0.425 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 0.495 1.070 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 0.495 2.275 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.495 3.155 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 -0.115 3.780 0.115 ;
        RECT  3.655 -0.115 3.725 0.425 ;
        RECT  3.370 -0.115 3.655 0.115 ;
        RECT  3.250 -0.115 3.370 0.235 ;
        RECT  2.990 -0.115 3.250 0.115 ;
        RECT  2.870 -0.115 2.990 0.235 ;
        RECT  2.585 -0.115 2.870 0.115 ;
        RECT  2.515 -0.115 2.585 0.255 ;
        RECT  2.405 -0.115 2.515 0.115 ;
        RECT  2.335 -0.115 2.405 0.255 ;
        RECT  2.050 -0.115 2.335 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.235 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.235 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.145 3.780 1.375 ;
        RECT  1.000 0.880 1.080 1.375 ;
        RECT  0.700 1.145 1.000 1.375 ;
        RECT  0.620 0.880 0.700 1.375 ;
        RECT  0.320 1.145 0.620 1.375 ;
        RECT  0.240 0.880 0.320 1.375 ;
        RECT  0.000 1.145 0.240 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.660 0.315 3.255 0.425 ;
        RECT  2.680 0.775 3.255 0.905 ;
        RECT  2.265 0.335 2.660 0.425 ;
        RECT  0.230 0.315 2.265 0.425 ;
        RECT  3.655 0.785 3.725 1.045 ;
        RECT  1.355 0.975 3.655 1.045 ;
        RECT  1.265 0.740 2.430 0.810 ;
        RECT  1.195 0.740 1.265 0.980 ;
        RECT  0.885 0.740 1.195 0.810 ;
        RECT  0.815 0.740 0.885 0.980 ;
        RECT  0.505 0.740 0.815 0.810 ;
        RECT  0.435 0.740 0.505 0.980 ;
        RECT  0.140 0.740 0.435 0.810 ;
        RECT  0.040 0.740 0.140 0.980 ;
    END
END NR3D6BWP40

MACRO NR3D8BWP40
    CLASS CORE ;
    FOREIGN NR3D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.900000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.375 0.745 4.760 0.905 ;
        RECT  4.375 0.315 4.750 0.425 ;
        RECT  4.165 0.315 4.375 0.905 ;
        RECT  3.475 0.315 4.165 0.425 ;
        RECT  3.500 0.745 4.165 0.905 ;
        RECT  3.090 0.335 3.475 0.425 ;
        RECT  0.290 0.315 3.090 0.425 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.215 0.495 1.475 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 0.495 3.095 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.455 0.495 3.975 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.950 -0.115 5.040 0.115 ;
        RECT  4.880 -0.115 4.950 0.425 ;
        RECT  4.570 -0.115 4.880 0.115 ;
        RECT  4.450 -0.115 4.570 0.230 ;
        RECT  4.190 -0.115 4.450 0.115 ;
        RECT  4.070 -0.115 4.190 0.230 ;
        RECT  3.810 -0.115 4.070 0.115 ;
        RECT  3.690 -0.115 3.810 0.230 ;
        RECT  3.405 -0.115 3.690 0.115 ;
        RECT  3.335 -0.115 3.405 0.255 ;
        RECT  3.225 -0.115 3.335 0.115 ;
        RECT  3.155 -0.115 3.225 0.255 ;
        RECT  2.870 -0.115 3.155 0.115 ;
        RECT  2.750 -0.115 2.870 0.230 ;
        RECT  2.490 -0.115 2.750 0.115 ;
        RECT  2.370 -0.115 2.490 0.230 ;
        RECT  2.110 -0.115 2.370 0.115 ;
        RECT  1.990 -0.115 2.110 0.230 ;
        RECT  1.730 -0.115 1.990 0.115 ;
        RECT  1.610 -0.115 1.730 0.230 ;
        RECT  1.350 -0.115 1.610 0.115 ;
        RECT  1.230 -0.115 1.350 0.230 ;
        RECT  0.970 -0.115 1.230 0.115 ;
        RECT  0.850 -0.115 0.970 0.230 ;
        RECT  0.590 -0.115 0.850 0.115 ;
        RECT  0.470 -0.115 0.590 0.230 ;
        RECT  0.155 -0.115 0.470 0.115 ;
        RECT  0.075 -0.115 0.155 0.425 ;
        RECT  0.000 -0.115 0.075 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.145 5.040 1.375 ;
        RECT  1.440 0.880 1.520 1.375 ;
        RECT  1.140 1.145 1.440 1.375 ;
        RECT  1.060 0.880 1.140 1.375 ;
        RECT  0.760 1.145 1.060 1.375 ;
        RECT  0.680 0.880 0.760 1.375 ;
        RECT  0.380 1.145 0.680 1.375 ;
        RECT  0.300 0.880 0.380 1.375 ;
        RECT  0.000 1.145 0.300 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.745 4.760 0.905 ;
        RECT  4.445 0.315 4.750 0.425 ;
        RECT  3.475 0.315 4.095 0.425 ;
        RECT  3.500 0.745 4.095 0.905 ;
        RECT  3.090 0.335 3.475 0.425 ;
        RECT  0.290 0.315 3.090 0.425 ;
        RECT  4.880 0.785 4.950 1.045 ;
        RECT  1.800 0.975 4.880 1.045 ;
        RECT  4.490 0.545 4.820 0.615 ;
        RECT  1.705 0.735 3.250 0.805 ;
        RECT  1.635 0.735 1.705 0.970 ;
        RECT  1.325 0.735 1.635 0.805 ;
        RECT  0.875 0.735 0.945 0.970 ;
        RECT  0.565 0.735 0.875 0.805 ;
        RECT  0.495 0.735 0.565 0.970 ;
        RECT  0.200 0.735 0.495 0.805 ;
        RECT  0.100 0.735 0.200 0.975 ;
        RECT  1.255 0.735 1.325 0.970 ;
        RECT  0.945 0.735 1.255 0.805 ;
    END
END NR3D8BWP40

MACRO NR4D0BWP40
    CLASS CORE ;
    FOREIGN NR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.084125 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.320 0.945 1.065 ;
        RECT  0.720 0.320 0.875 0.390 ;
        RECT  0.810 0.995 0.875 1.065 ;
        RECT  0.640 0.195 0.720 0.390 ;
        RECT  0.320 0.320 0.640 0.390 ;
        RECT  0.245 0.200 0.320 0.390 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.820 -0.115 0.940 0.240 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.240 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.145 0.980 1.375 ;
        RECT  0.040 0.985 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END NR4D0BWP40

MACRO NR4D1BWP40
    CLASS CORE ;
    FOREIGN NR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.168250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.320 0.945 1.065 ;
        RECT  0.320 0.320 0.875 0.390 ;
        RECT  0.810 0.995 0.875 1.065 ;
        RECT  0.245 0.255 0.320 0.390 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.820 -0.115 0.940 0.240 ;
        RECT  0.540 -0.115 0.820 0.115 ;
        RECT  0.420 -0.115 0.540 0.240 ;
        RECT  0.140 -0.115 0.420 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.145 0.980 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
END NR4D1BWP40

MACRO NR4D2BWP40
    CLASS CORE ;
    FOREIGN NR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.277500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.185 1.690 0.425 ;
        RECT  1.300 0.355 1.590 0.425 ;
        RECT  1.220 0.185 1.300 0.425 ;
        RECT  0.740 0.355 1.220 0.425 ;
        RECT  0.660 0.185 0.740 0.425 ;
        RECT  0.385 0.355 0.660 0.425 ;
        RECT  0.355 0.355 0.385 0.915 ;
        RECT  0.315 0.225 0.355 0.915 ;
        RECT  0.285 0.225 0.315 0.425 ;
        RECT  0.260 0.845 0.315 0.915 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.495 1.785 0.625 ;
        RECT  1.570 0.495 1.655 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.285 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.285 0.615 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.775 0.615 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.780 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.910 -0.115 1.960 0.115 ;
        RECT  1.810 -0.115 1.910 0.415 ;
        RECT  1.490 -0.115 1.810 0.115 ;
        RECT  1.410 -0.115 1.490 0.285 ;
        RECT  1.110 -0.115 1.410 0.115 ;
        RECT  1.030 -0.115 1.110 0.285 ;
        RECT  0.930 -0.115 1.030 0.115 ;
        RECT  0.850 -0.115 0.930 0.285 ;
        RECT  0.550 -0.115 0.850 0.115 ;
        RECT  0.470 -0.115 0.550 0.285 ;
        RECT  0.150 -0.115 0.470 0.115 ;
        RECT  0.050 -0.115 0.150 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.145 1.960 1.375 ;
        RECT  1.600 0.975 1.680 1.375 ;
        RECT  0.000 1.145 1.600 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.810 0.835 1.910 1.075 ;
        RECT  1.490 0.835 1.810 0.905 ;
        RECT  1.410 0.835 1.490 1.065 ;
        RECT  1.015 0.995 1.410 1.065 ;
        RECT  0.635 0.835 1.320 0.905 ;
        RECT  0.040 0.995 0.945 1.065 ;
    END
END NR4D2BWP40

MACRO NR4D3BWP40
    CLASS CORE ;
    FOREIGN NR4D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.492250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.300 2.450 0.415 ;
        RECT  0.385 0.300 0.595 0.905 ;
        RECT  0.150 0.300 0.385 0.415 ;
        RECT  0.160 0.835 0.385 0.905 ;
        RECT  0.060 0.835 0.160 1.075 ;
        RECT  0.070 0.225 0.150 0.415 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.495 2.345 0.625 ;
        RECT  1.985 0.495 2.065 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.725 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 1.140 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.495 0.305 0.625 ;
        RECT  0.035 0.495 0.125 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.260 -0.115 2.520 0.115 ;
        RECT  2.140 -0.115 2.260 0.230 ;
        RECT  1.880 -0.115 2.140 0.115 ;
        RECT  1.760 -0.115 1.880 0.230 ;
        RECT  1.500 -0.115 1.760 0.115 ;
        RECT  1.380 -0.115 1.500 0.230 ;
        RECT  1.120 -0.115 1.380 0.115 ;
        RECT  1.000 -0.115 1.120 0.230 ;
        RECT  0.740 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.740 0.230 ;
        RECT  0.360 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.360 0.230 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.145 2.520 1.375 ;
        RECT  2.370 0.725 2.450 1.375 ;
        RECT  2.070 1.145 2.370 1.375 ;
        RECT  1.950 1.015 2.070 1.375 ;
        RECT  0.000 1.145 1.950 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.300 2.450 0.415 ;
        RECT  0.150 0.300 0.315 0.415 ;
        RECT  0.160 0.835 0.315 0.905 ;
        RECT  0.060 0.835 0.160 1.075 ;
        RECT  0.070 0.225 0.150 0.415 ;
        RECT  2.165 0.845 2.255 1.075 ;
        RECT  1.860 0.845 2.165 0.915 ;
        RECT  1.780 0.845 1.860 1.055 ;
        RECT  1.380 0.985 1.780 1.055 ;
        RECT  1.290 0.845 1.690 0.915 ;
        RECT  1.210 0.845 1.290 1.075 ;
        RECT  0.780 0.845 1.210 0.915 ;
        RECT  0.240 0.985 1.120 1.055 ;
    END
END NR4D3BWP40

MACRO NR4D4BWP40
    CLASS CORE ;
    FOREIGN NR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.525000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.305 3.255 0.420 ;
        RECT  0.595 0.830 0.720 0.915 ;
        RECT  0.385 0.305 0.595 0.915 ;
        RECT  0.245 0.305 0.385 0.420 ;
        RECT  0.220 0.830 0.385 0.915 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.495 3.325 0.630 ;
        RECT  2.830 0.495 2.910 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.075 0.495 2.555 0.630 ;
        RECT  1.995 0.495 2.075 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.495 1.460 0.625 ;
        RECT  1.010 0.495 1.090 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.255 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.115 3.500 0.115 ;
        RECT  3.375 -0.115 3.445 0.420 ;
        RECT  3.090 -0.115 3.375 0.115 ;
        RECT  2.970 -0.115 3.090 0.235 ;
        RECT  2.710 -0.115 2.970 0.115 ;
        RECT  2.590 -0.115 2.710 0.235 ;
        RECT  2.330 -0.115 2.590 0.115 ;
        RECT  2.210 -0.115 2.330 0.235 ;
        RECT  1.950 -0.115 2.210 0.115 ;
        RECT  1.830 -0.115 1.950 0.235 ;
        RECT  1.670 -0.115 1.830 0.115 ;
        RECT  1.545 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.545 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.235 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.235 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.145 3.500 1.375 ;
        RECT  3.160 0.985 3.280 1.375 ;
        RECT  2.900 1.145 3.160 1.375 ;
        RECT  2.780 0.985 2.900 1.375 ;
        RECT  0.000 1.145 2.780 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.305 3.255 0.420 ;
        RECT  0.665 0.830 0.720 0.915 ;
        RECT  0.245 0.305 0.315 0.420 ;
        RECT  0.220 0.830 0.315 0.915 ;
        RECT  3.375 0.845 3.465 1.075 ;
        RECT  3.070 0.845 3.375 0.915 ;
        RECT  2.990 0.845 3.070 1.075 ;
        RECT  2.690 0.845 2.990 0.915 ;
        RECT  2.610 0.845 2.690 1.075 ;
        RECT  1.830 0.845 2.610 0.915 ;
        RECT  0.980 0.985 2.520 1.055 ;
        RECT  0.885 0.845 1.670 0.915 ;
        RECT  0.815 0.845 0.885 1.055 ;
        RECT  0.130 0.985 0.815 1.055 ;
        RECT  0.050 0.865 0.130 1.055 ;
    END
END NR4D4BWP40

MACRO NR4D6BWP40
    CLASS CORE ;
    FOREIGN NR4D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.787500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.305 4.795 0.420 ;
        RECT  0.595 0.840 1.100 0.915 ;
        RECT  0.385 0.305 0.595 0.915 ;
        RECT  0.245 0.305 0.385 0.420 ;
        RECT  0.220 0.830 0.385 0.915 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 0.495 4.865 0.625 ;
        RECT  4.440 0.495 4.520 0.765 ;
        RECT  3.955 0.495 4.440 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.330 0.495 3.745 0.625 ;
        RECT  3.250 0.495 3.330 0.765 ;
        RECT  2.770 0.495 3.250 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 0.495 2.265 0.625 ;
        RECT  1.710 0.495 1.790 0.765 ;
        RECT  1.295 0.495 1.710 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.182400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.495 1.145 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.985 0.435 ;
        RECT  4.630 -0.115 4.915 0.115 ;
        RECT  4.510 -0.115 4.630 0.235 ;
        RECT  4.250 -0.115 4.510 0.115 ;
        RECT  4.130 -0.115 4.250 0.235 ;
        RECT  3.870 -0.115 4.130 0.115 ;
        RECT  3.750 -0.115 3.870 0.235 ;
        RECT  3.490 -0.115 3.750 0.115 ;
        RECT  3.370 -0.115 3.490 0.235 ;
        RECT  3.110 -0.115 3.370 0.115 ;
        RECT  2.990 -0.115 3.110 0.235 ;
        RECT  2.710 -0.115 2.990 0.115 ;
        RECT  2.590 -0.115 2.710 0.235 ;
        RECT  2.455 -0.115 2.590 0.115 ;
        RECT  2.335 -0.115 2.455 0.235 ;
        RECT  2.050 -0.115 2.335 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.235 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.235 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 1.145 5.040 1.375 ;
        RECT  4.700 0.985 4.820 1.375 ;
        RECT  4.440 1.145 4.700 1.375 ;
        RECT  4.320 0.985 4.440 1.375 ;
        RECT  4.060 1.145 4.320 1.375 ;
        RECT  3.940 0.985 4.060 1.375 ;
        RECT  0.000 1.145 3.940 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.665 0.305 4.795 0.420 ;
        RECT  0.665 0.840 1.100 0.915 ;
        RECT  0.245 0.305 0.315 0.420 ;
        RECT  0.220 0.830 0.315 0.915 ;
        RECT  4.915 0.845 5.005 1.075 ;
        RECT  4.610 0.845 4.915 0.915 ;
        RECT  4.530 0.845 4.610 1.075 ;
        RECT  4.230 0.845 4.530 0.915 ;
        RECT  4.150 0.845 4.230 1.075 ;
        RECT  3.850 0.845 4.150 0.915 ;
        RECT  3.770 0.845 3.850 1.075 ;
        RECT  2.610 0.845 3.770 0.915 ;
        RECT  1.360 0.985 3.680 1.055 ;
        RECT  1.265 0.845 2.440 0.915 ;
        RECT  1.195 0.845 1.265 1.055 ;
        RECT  0.130 0.985 1.195 1.055 ;
        RECT  0.050 0.865 0.130 1.055 ;
    END
END NR4D6BWP40

MACRO NR4D8BWP40
    CLASS CORE ;
    FOREIGN NR4D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.050000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.305 6.315 0.420 ;
        RECT  1.015 0.835 1.480 0.915 ;
        RECT  0.805 0.305 1.015 0.915 ;
        RECT  0.245 0.305 0.805 0.420 ;
        RECT  0.220 0.835 0.805 0.915 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.780 0.495 6.405 0.630 ;
        RECT  5.700 0.495 5.780 0.765 ;
        RECT  5.040 0.495 5.700 0.630 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.495 4.865 0.630 ;
        RECT  4.370 0.495 4.450 0.765 ;
        RECT  3.530 0.495 4.370 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.495 2.995 0.625 ;
        RECT  2.130 0.495 2.210 0.765 ;
        RECT  1.675 0.495 2.130 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.243200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.680 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 -0.115 6.580 0.115 ;
        RECT  6.455 -0.115 6.525 0.420 ;
        RECT  6.150 -0.115 6.455 0.115 ;
        RECT  6.030 -0.115 6.150 0.235 ;
        RECT  5.770 -0.115 6.030 0.115 ;
        RECT  5.650 -0.115 5.770 0.235 ;
        RECT  5.390 -0.115 5.650 0.115 ;
        RECT  5.270 -0.115 5.390 0.235 ;
        RECT  5.010 -0.115 5.270 0.115 ;
        RECT  4.890 -0.115 5.010 0.235 ;
        RECT  4.630 -0.115 4.890 0.115 ;
        RECT  4.510 -0.115 4.630 0.235 ;
        RECT  4.250 -0.115 4.510 0.115 ;
        RECT  4.130 -0.115 4.250 0.235 ;
        RECT  3.870 -0.115 4.130 0.115 ;
        RECT  3.750 -0.115 3.870 0.235 ;
        RECT  3.490 -0.115 3.750 0.115 ;
        RECT  3.370 -0.115 3.490 0.235 ;
        RECT  3.190 -0.115 3.370 0.115 ;
        RECT  3.070 -0.115 3.190 0.235 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.235 ;
        RECT  2.430 -0.115 2.690 0.115 ;
        RECT  2.310 -0.115 2.430 0.235 ;
        RECT  2.050 -0.115 2.310 0.115 ;
        RECT  1.930 -0.115 2.050 0.235 ;
        RECT  1.670 -0.115 1.930 0.115 ;
        RECT  1.550 -0.115 1.670 0.235 ;
        RECT  1.290 -0.115 1.550 0.115 ;
        RECT  1.170 -0.115 1.290 0.235 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.235 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.235 ;
        RECT  0.140 -0.115 0.410 0.115 ;
        RECT  0.040 -0.115 0.140 0.415 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.340 1.145 6.580 1.375 ;
        RECT  6.220 0.985 6.340 1.375 ;
        RECT  5.960 1.145 6.220 1.375 ;
        RECT  5.840 0.985 5.960 1.375 ;
        RECT  5.580 1.145 5.840 1.375 ;
        RECT  5.460 0.985 5.580 1.375 ;
        RECT  5.200 1.145 5.460 1.375 ;
        RECT  5.080 0.985 5.200 1.375 ;
        RECT  0.000 1.145 5.080 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 0.305 6.315 0.420 ;
        RECT  1.085 0.835 1.480 0.915 ;
        RECT  0.245 0.305 0.735 0.420 ;
        RECT  0.220 0.835 0.735 0.915 ;
        RECT  6.455 0.845 6.545 1.075 ;
        RECT  6.130 0.845 6.455 0.915 ;
        RECT  6.050 0.845 6.130 1.075 ;
        RECT  5.750 0.845 6.050 0.915 ;
        RECT  5.670 0.845 5.750 1.075 ;
        RECT  5.370 0.845 5.670 0.915 ;
        RECT  5.290 0.845 5.370 1.075 ;
        RECT  4.990 0.845 5.290 0.915 ;
        RECT  4.910 0.845 4.990 1.075 ;
        RECT  3.370 0.845 4.910 0.915 ;
        RECT  1.740 0.985 4.820 1.055 ;
        RECT  1.645 0.845 3.190 0.915 ;
        RECT  1.575 0.845 1.645 1.055 ;
        RECT  0.130 0.985 1.575 1.055 ;
        RECT  1.090 0.495 1.560 0.630 ;
        RECT  0.050 0.865 0.130 1.055 ;
    END
END NR4D8BWP40

MACRO OA211D0BWP40
    CLASS CORE ;
    FOREIGN OA211D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.077700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.195 1.225 1.065 ;
        RECT  1.030 0.195 1.155 0.265 ;
        RECT  1.115 0.995 1.155 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.805 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 -0.115 1.260 0.115 ;
        RECT  0.870 -0.115 0.950 0.265 ;
        RECT  0.000 -0.115 0.870 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.145 1.260 1.375 ;
        RECT  0.830 1.050 0.950 1.375 ;
        RECT  0.550 1.145 0.830 1.375 ;
        RECT  0.430 1.050 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.045 0.345 1.085 0.835 ;
        RECT  1.015 0.345 1.045 0.975 ;
        RECT  0.220 0.345 1.015 0.415 ;
        RECT  0.975 0.770 1.015 0.975 ;
        RECT  0.130 0.905 0.975 0.975 ;
        RECT  0.035 0.200 0.540 0.270 ;
        RECT  0.050 0.905 0.130 1.060 ;
    END
END OA211D0BWP40

MACRO OA211D1BWP40
    CLASS CORE ;
    FOREIGN OA211D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.148000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.195 1.225 1.065 ;
        RECT  1.030 0.195 1.155 0.265 ;
        RECT  1.115 0.995 1.155 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.805 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 -0.115 1.260 0.115 ;
        RECT  0.865 -0.115 0.945 0.265 ;
        RECT  0.000 -0.115 0.865 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.145 1.260 1.375 ;
        RECT  0.830 1.050 0.950 1.375 ;
        RECT  0.550 1.145 0.830 1.375 ;
        RECT  0.430 1.050 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.045 0.345 1.085 0.865 ;
        RECT  1.015 0.345 1.045 0.975 ;
        RECT  0.220 0.345 1.015 0.415 ;
        RECT  0.975 0.785 1.015 0.975 ;
        RECT  0.130 0.905 0.975 0.975 ;
        RECT  0.130 0.200 0.540 0.270 ;
        RECT  0.055 0.200 0.130 0.400 ;
        RECT  0.055 0.905 0.130 1.060 ;
    END
END OA211D1BWP40

MACRO OA211D2BWP40
    CLASS CORE ;
    FOREIGN OA211D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.205 0.495 1.365 0.625 ;
        RECT  1.135 0.195 1.205 1.065 ;
        RECT  1.030 0.195 1.135 0.265 ;
        RECT  1.030 0.985 1.135 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.840 0.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.695 0.425 0.765 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.275 -0.115 1.345 0.400 ;
        RECT  0.920 -0.115 1.275 0.115 ;
        RECT  0.840 -0.115 0.920 0.265 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.275 0.720 1.345 1.375 ;
        RECT  0.930 1.145 1.275 1.375 ;
        RECT  0.850 0.985 0.930 1.375 ;
        RECT  0.550 1.145 0.850 1.375 ;
        RECT  0.430 1.010 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.345 1.055 0.915 ;
        RECT  0.220 0.345 0.985 0.415 ;
        RECT  0.035 0.845 0.985 0.915 ;
        RECT  0.130 0.200 0.540 0.270 ;
        RECT  0.055 0.200 0.130 0.370 ;
    END
END OA211D2BWP40

MACRO OA211D4BWP40
    CLASS CORE ;
    FOREIGN OA211D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.415 1.035 ;
        RECT  2.205 0.355 2.325 0.790 ;
        RECT  2.015 0.355 2.205 0.465 ;
        RECT  2.015 0.695 2.205 0.790 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.695 2.015 1.035 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.375 0.495 0.665 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.255 0.695 0.735 0.765 ;
        RECT  0.165 0.495 0.255 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.390 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.575 0.765 ;
        RECT  0.995 0.695 1.505 0.765 ;
        RECT  0.875 0.495 0.995 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.475 ;
        RECT  2.230 -0.115 2.530 0.115 ;
        RECT  2.110 -0.115 2.230 0.280 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.740 -0.115 1.840 0.275 ;
        RECT  0.530 -0.115 1.740 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.675 2.610 1.375 ;
        RECT  2.230 1.145 2.530 1.375 ;
        RECT  2.110 0.885 2.230 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.740 0.975 1.840 1.375 ;
        RECT  1.660 1.145 1.740 1.375 ;
        RECT  1.560 0.975 1.660 1.375 ;
        RECT  0.900 1.145 1.560 1.375 ;
        RECT  0.800 0.975 0.900 1.375 ;
        RECT  0.520 1.145 0.800 1.375 ;
        RECT  0.420 0.975 0.520 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.835 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.015 0.355 2.135 0.465 ;
        RECT  2.015 0.695 2.135 0.790 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.695 2.015 1.035 ;
        RECT  1.715 0.545 2.060 0.615 ;
        RECT  1.645 0.345 1.715 0.905 ;
        RECT  0.885 0.195 1.670 0.265 ;
        RECT  0.980 0.345 1.645 0.415 ;
        RECT  1.280 0.835 1.645 0.905 ;
        RECT  1.180 0.835 1.280 1.075 ;
        RECT  0.710 0.835 1.180 0.905 ;
        RECT  0.815 0.195 0.885 0.415 ;
        RECT  0.130 0.345 0.815 0.415 ;
        RECT  0.610 0.835 0.710 1.075 ;
        RECT  0.330 0.835 0.610 0.905 ;
        RECT  0.230 0.835 0.330 1.075 ;
        RECT  0.050 0.265 0.130 0.415 ;
    END
END OA211D4BWP40

MACRO OA21D0BWP40
    CLASS CORE ;
    FOREIGN OA21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.050500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.185 0.945 1.075 ;
        RECT  0.855 0.185 0.875 0.295 ;
        RECT  0.855 0.965 0.875 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.980 0.115 ;
        RECT  0.610 -0.115 0.730 0.275 ;
        RECT  0.000 -0.115 0.610 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.145 0.980 1.375 ;
        RECT  0.610 0.985 0.730 1.375 ;
        RECT  0.140 1.145 0.610 1.375 ;
        RECT  0.040 0.960 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.915 ;
        RECT  0.215 0.345 0.735 0.415 ;
        RECT  0.530 0.845 0.735 0.915 ;
        RECT  0.035 0.195 0.530 0.265 ;
        RECT  0.455 0.845 0.530 1.055 ;
        RECT  0.390 0.985 0.455 1.055 ;
    END
END OA21D0BWP40

MACRO OA21D1BWP40
    CLASS CORE ;
    FOREIGN OA21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.101000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.195 0.945 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.580 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 -0.115 0.980 0.115 ;
        RECT  0.610 -0.115 0.730 0.275 ;
        RECT  0.000 -0.115 0.610 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.145 0.980 1.375 ;
        RECT  0.610 0.985 0.730 1.375 ;
        RECT  0.140 1.145 0.610 1.375 ;
        RECT  0.040 0.960 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.705 0.345 0.775 0.915 ;
        RECT  0.215 0.345 0.705 0.415 ;
        RECT  0.530 0.845 0.705 0.915 ;
        RECT  0.035 0.195 0.530 0.265 ;
        RECT  0.455 0.845 0.530 1.055 ;
        RECT  0.390 0.985 0.455 1.055 ;
    END
END OA21D1BWP40

MACRO OA21D2BWP40
    CLASS CORE ;
    FOREIGN OA21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.195 0.945 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.805 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.200 -0.115 1.260 0.115 ;
        RECT  1.120 -0.115 1.200 0.425 ;
        RECT  0.730 -0.115 1.120 0.115 ;
        RECT  0.610 -0.115 0.730 0.275 ;
        RECT  0.000 -0.115 0.610 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.205 1.145 1.260 1.375 ;
        RECT  1.135 0.695 1.205 1.375 ;
        RECT  0.730 1.145 1.135 1.375 ;
        RECT  0.610 1.000 0.730 1.375 ;
        RECT  0.125 1.145 0.610 1.375 ;
        RECT  0.055 0.865 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.345 0.805 0.915 ;
        RECT  0.215 0.345 0.735 0.415 ;
        RECT  0.530 0.845 0.735 0.915 ;
        RECT  0.135 0.195 0.530 0.265 ;
        RECT  0.455 0.845 0.530 0.985 ;
        RECT  0.415 0.915 0.455 0.985 ;
        RECT  0.050 0.195 0.135 0.375 ;
    END
END OA21D2BWP40

MACRO OA21D4BWP40
    CLASS CORE ;
    FOREIGN OA21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.185 1.995 1.045 ;
        RECT  1.855 0.355 1.865 1.045 ;
        RECT  1.785 0.355 1.855 0.810 ;
        RECT  1.535 0.355 1.785 0.465 ;
        RECT  1.535 0.695 1.785 0.810 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.695 1.535 1.010 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.065 0.495 1.225 0.915 ;
        RECT  0.245 0.845 1.065 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.125 0.495 0.175 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.515 0.495 0.805 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.980 0.775 ;
        RECT  0.405 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.405 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 -0.115 2.240 0.115 ;
        RECT  2.090 -0.115 2.170 0.475 ;
        RECT  1.760 -0.115 2.090 0.115 ;
        RECT  1.640 -0.115 1.760 0.275 ;
        RECT  1.340 -0.115 1.640 0.115 ;
        RECT  1.220 -0.115 1.340 0.275 ;
        RECT  0.130 -0.115 1.220 0.115 ;
        RECT  0.050 -0.115 0.130 0.425 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.145 2.240 1.375 ;
        RECT  2.090 0.675 2.170 1.375 ;
        RECT  1.760 1.145 2.090 1.375 ;
        RECT  1.640 0.880 1.760 1.375 ;
        RECT  1.340 1.145 1.640 1.375 ;
        RECT  1.220 1.125 1.340 1.375 ;
        RECT  0.730 1.145 1.220 1.375 ;
        RECT  0.610 1.125 0.730 1.375 ;
        RECT  0.120 1.145 0.610 1.375 ;
        RECT  0.050 0.960 0.120 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.535 0.355 1.715 0.465 ;
        RECT  1.535 0.695 1.715 0.810 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.695 1.535 1.010 ;
        RECT  1.375 0.545 1.635 0.615 ;
        RECT  1.305 0.345 1.375 1.055 ;
        RECT  0.410 0.345 1.305 0.415 ;
        RECT  0.220 0.985 1.305 1.055 ;
        RECT  0.315 0.205 1.120 0.275 ;
        RECT  0.240 0.205 0.315 0.365 ;
    END
END OA21D4BWP40

MACRO OA221D0BWP40
    CLASS CORE ;
    FOREIGN OA221D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.075 ;
        RECT  1.415 0.185 1.435 0.305 ;
        RECT  1.415 0.945 1.435 1.075 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.355 1.365 0.495 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.085 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.805 0.625 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 0.355 0.525 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.280 0.250 ;
        RECT  0.000 -0.115 1.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.145 1.540 1.375 ;
        RECT  1.200 0.990 1.280 1.375 ;
        RECT  0.710 1.145 1.200 1.375 ;
        RECT  0.590 1.115 0.710 1.375 ;
        RECT  0.140 1.145 0.590 1.375 ;
        RECT  0.040 0.965 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.275 0.620 1.345 0.905 ;
        RECT  1.110 0.835 1.275 0.905 ;
        RECT  1.040 0.835 1.110 0.990 ;
        RECT  1.000 0.185 1.080 0.415 ;
        RECT  0.340 0.920 1.040 0.990 ;
        RECT  0.615 0.345 1.000 0.415 ;
        RECT  0.035 0.195 0.920 0.265 ;
        RECT  0.270 0.350 0.340 0.990 ;
    END
END OA221D0BWP40

MACRO OA221D1BWP40
    CLASS CORE ;
    FOREIGN OA221D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.108000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.185 1.505 1.065 ;
        RECT  1.415 0.185 1.435 0.300 ;
        RECT  1.395 0.995 1.435 1.065 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.495 1.225 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.975 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.805 0.625 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 0.355 0.525 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.280 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.280 0.395 ;
        RECT  0.000 -0.115 1.200 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.180 1.045 1.300 1.375 ;
        RECT  0.730 1.145 1.180 1.375 ;
        RECT  0.610 1.045 0.730 1.375 ;
        RECT  0.140 1.145 0.610 1.375 ;
        RECT  0.040 0.940 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.520 1.365 0.915 ;
        RECT  1.215 0.845 1.295 0.915 ;
        RECT  1.145 0.845 1.215 0.945 ;
        RECT  1.085 0.875 1.145 0.945 ;
        RECT  0.995 0.185 1.115 0.415 ;
        RECT  1.015 0.875 1.085 1.045 ;
        RECT  0.525 0.875 1.015 0.945 ;
        RECT  0.615 0.345 0.995 0.415 ;
        RECT  0.130 0.195 0.920 0.265 ;
        RECT  0.415 0.875 0.525 1.045 ;
        RECT  0.340 0.875 0.415 0.945 ;
        RECT  0.270 0.350 0.340 0.945 ;
        RECT  0.050 0.195 0.130 0.395 ;
    END
END OA221D1BWP40

MACRO OA221D2BWP40
    CLASS CORE ;
    FOREIGN OA221D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.128000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.585 0.495 1.785 0.625 ;
        RECT  1.505 0.185 1.585 1.075 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.495 1.225 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.975 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 0.355 0.525 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.115 1.820 0.115 ;
        RECT  1.695 -0.115 1.765 0.410 ;
        RECT  1.350 -0.115 1.695 0.115 ;
        RECT  1.270 -0.115 1.350 0.435 ;
        RECT  0.000 -0.115 1.270 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 1.145 1.820 1.375 ;
        RECT  1.695 0.720 1.765 1.375 ;
        RECT  1.370 1.145 1.695 1.375 ;
        RECT  1.250 0.975 1.370 1.375 ;
        RECT  0.710 1.145 1.250 1.375 ;
        RECT  0.590 0.985 0.710 1.375 ;
        RECT  0.125 1.145 0.590 1.375 ;
        RECT  0.055 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.355 0.520 1.425 0.905 ;
        RECT  1.125 0.835 1.355 0.905 ;
        RECT  1.035 0.185 1.145 0.415 ;
        RECT  1.055 0.835 1.125 1.065 ;
        RECT  0.505 0.835 1.055 0.905 ;
        RECT  0.615 0.345 1.035 0.415 ;
        RECT  0.130 0.195 0.920 0.265 ;
        RECT  0.435 0.835 0.505 1.065 ;
        RECT  0.340 0.835 0.435 0.905 ;
        RECT  0.270 0.350 0.340 0.905 ;
        RECT  0.050 0.195 0.130 0.395 ;
    END
END OA221D2BWP40

MACRO OA221D4BWP40
    CLASS CORE ;
    FOREIGN OA221D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.185 2.835 0.465 ;
        RECT  2.825 0.695 2.835 1.035 ;
        RECT  2.765 0.185 2.825 1.035 ;
        RECT  2.625 0.355 2.765 0.815 ;
        RECT  2.455 0.355 2.625 0.465 ;
        RECT  2.455 0.695 2.625 0.815 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.695 2.455 1.035 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.065 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.435 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.545 0.495 1.645 0.775 ;
        RECT  1.085 0.705 1.545 0.775 ;
        RECT  0.990 0.495 1.085 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.495 0.760 0.640 ;
        RECT  0.625 0.495 0.695 0.775 ;
        RECT  0.245 0.705 0.625 0.775 ;
        RECT  0.155 0.495 0.245 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.635 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.475 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.550 -0.115 2.670 0.280 ;
        RECT  2.270 -0.115 2.550 0.115 ;
        RECT  2.190 -0.115 2.270 0.435 ;
        RECT  1.900 -0.115 2.190 0.115 ;
        RECT  1.800 -0.115 1.900 0.275 ;
        RECT  0.000 -0.115 1.800 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.675 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.550 0.885 2.670 1.375 ;
        RECT  2.290 1.145 2.550 1.375 ;
        RECT  2.170 0.985 2.290 1.375 ;
        RECT  1.900 1.145 2.170 1.375 ;
        RECT  1.800 0.985 1.900 1.375 ;
        RECT  1.720 1.145 1.800 1.375 ;
        RECT  1.620 0.985 1.720 1.375 ;
        RECT  0.940 1.145 1.620 1.375 ;
        RECT  0.820 1.025 0.940 1.375 ;
        RECT  0.140 1.145 0.820 1.375 ;
        RECT  0.040 0.855 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.455 0.355 2.555 0.465 ;
        RECT  2.455 0.695 2.555 0.815 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.695 2.455 1.035 ;
        RECT  2.300 0.545 2.430 0.615 ;
        RECT  2.230 0.545 2.300 0.915 ;
        RECT  2.080 0.845 2.230 0.915 ;
        RECT  1.990 0.185 2.090 0.425 ;
        RECT  2.000 0.845 2.080 1.075 ;
        RECT  0.910 0.845 2.000 0.915 ;
        RECT  1.040 0.355 1.990 0.425 ;
        RECT  0.130 0.205 1.730 0.275 ;
        RECT  1.040 0.995 1.545 1.065 ;
        RECT  0.840 0.345 0.910 0.915 ;
        RECT  0.220 0.345 0.840 0.415 ;
        RECT  0.410 0.845 0.840 0.915 ;
        RECT  0.220 0.985 0.725 1.055 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA221D4BWP40

MACRO OA222D0BWP40
    CLASS CORE ;
    FOREIGN OA222D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.062000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.195 1.785 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.435 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 -0.115 1.820 0.115 ;
        RECT  1.445 -0.115 1.525 0.290 ;
        RECT  1.145 -0.115 1.445 0.115 ;
        RECT  1.025 -0.115 1.145 0.230 ;
        RECT  0.000 -0.115 1.025 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.145 1.820 1.375 ;
        RECT  1.425 0.985 1.545 1.375 ;
        RECT  0.965 1.145 1.425 1.375 ;
        RECT  0.845 1.115 0.965 1.375 ;
        RECT  0.170 1.145 0.845 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.520 0.520 1.590 0.915 ;
        RECT  1.320 0.845 1.520 0.915 ;
        RECT  1.245 0.195 1.345 0.415 ;
        RECT  1.250 0.845 1.320 1.045 ;
        RECT  0.395 0.975 1.250 1.045 ;
        RECT  0.620 0.345 1.245 0.415 ;
        RECT  0.050 0.195 0.945 0.265 ;
        RECT  0.325 0.890 0.395 1.045 ;
        RECT  0.105 0.345 0.360 0.415 ;
        RECT  0.105 0.890 0.325 0.960 ;
        RECT  0.035 0.345 0.105 0.960 ;
    END
END OA222D0BWP40

MACRO OA222D1BWP40
    CLASS CORE ;
    FOREIGN OA222D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.124000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.195 1.785 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.630 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.435 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.905 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.023000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 -0.115 1.820 0.115 ;
        RECT  1.445 -0.115 1.525 0.400 ;
        RECT  1.145 -0.115 1.445 0.115 ;
        RECT  1.025 -0.115 1.145 0.265 ;
        RECT  0.000 -0.115 1.025 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.145 1.820 1.375 ;
        RECT  1.425 0.985 1.545 1.375 ;
        RECT  0.965 1.145 1.425 1.375 ;
        RECT  0.845 1.115 0.965 1.375 ;
        RECT  0.170 1.145 0.845 1.375 ;
        RECT  0.050 1.030 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.520 0.520 1.590 0.915 ;
        RECT  1.320 0.845 1.520 0.915 ;
        RECT  0.620 0.345 1.355 0.415 ;
        RECT  1.250 0.845 1.320 1.045 ;
        RECT  0.395 0.975 1.250 1.045 ;
        RECT  0.050 0.195 0.945 0.265 ;
        RECT  0.325 0.890 0.395 1.045 ;
        RECT  0.105 0.345 0.360 0.415 ;
        RECT  0.105 0.890 0.325 0.960 ;
        RECT  0.035 0.345 0.105 0.960 ;
    END
END OA222D1BWP40

MACRO OA222D2BWP40
    CLASS CORE ;
    FOREIGN OA222D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.495 1.925 0.625 ;
        RECT  1.645 0.195 1.730 1.045 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.090 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.435 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.700 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.495 0.945 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.290 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.905 -0.115 1.960 0.115 ;
        RECT  1.835 -0.115 1.905 0.415 ;
        RECT  1.520 -0.115 1.835 0.115 ;
        RECT  1.450 -0.115 1.520 0.405 ;
        RECT  1.145 -0.115 1.450 0.115 ;
        RECT  1.025 -0.115 1.145 0.265 ;
        RECT  0.000 -0.115 1.025 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.145 1.960 1.375 ;
        RECT  1.830 0.720 1.900 1.375 ;
        RECT  1.550 1.145 1.830 1.375 ;
        RECT  1.420 0.985 1.550 1.375 ;
        RECT  0.965 1.145 1.420 1.375 ;
        RECT  0.845 0.995 0.965 1.375 ;
        RECT  0.170 1.145 0.845 1.375 ;
        RECT  0.050 0.995 0.170 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.520 1.575 0.915 ;
        RECT  1.120 0.845 1.505 0.915 ;
        RECT  0.620 0.345 1.335 0.415 ;
        RECT  1.050 0.845 1.120 1.075 ;
        RECT  0.525 0.845 1.050 0.915 ;
        RECT  0.525 0.195 0.945 0.265 ;
        RECT  0.455 0.195 0.525 0.425 ;
        RECT  0.455 0.845 0.525 1.075 ;
        RECT  0.050 0.195 0.455 0.265 ;
        RECT  0.105 0.845 0.455 0.915 ;
        RECT  0.105 0.345 0.360 0.415 ;
        RECT  0.035 0.345 0.105 0.915 ;
    END
END OA222D2BWP40

MACRO OA222D4BWP40
    CLASS CORE ;
    FOREIGN OA222D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.185 3.255 0.465 ;
        RECT  3.245 0.695 3.255 1.035 ;
        RECT  3.185 0.185 3.245 1.035 ;
        RECT  3.045 0.355 3.185 0.815 ;
        RECT  2.875 0.355 3.045 0.465 ;
        RECT  2.875 0.695 3.045 0.815 ;
        RECT  2.805 0.185 2.875 0.465 ;
        RECT  2.805 0.695 2.875 1.035 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.365 0.640 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.475 0.495 2.555 0.785 ;
        RECT  2.065 0.715 2.475 0.785 ;
        RECT  1.945 0.495 2.065 0.785 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.380 0.635 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.495 1.645 0.785 ;
        RECT  1.055 0.715 1.560 0.785 ;
        RECT  0.985 0.495 1.055 0.785 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.495 0.760 0.640 ;
        RECT  0.625 0.495 0.695 0.785 ;
        RECT  0.245 0.715 0.625 0.785 ;
        RECT  0.155 0.495 0.245 0.785 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.645 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.475 ;
        RECT  3.090 -0.115 3.370 0.115 ;
        RECT  2.970 -0.115 3.090 0.280 ;
        RECT  2.680 -0.115 2.970 0.115 ;
        RECT  2.600 -0.115 2.680 0.425 ;
        RECT  2.290 -0.115 2.600 0.115 ;
        RECT  2.210 -0.115 2.290 0.285 ;
        RECT  1.910 -0.115 2.210 0.115 ;
        RECT  1.830 -0.115 1.910 0.285 ;
        RECT  0.000 -0.115 1.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.675 3.450 1.375 ;
        RECT  3.090 1.145 3.370 1.375 ;
        RECT  2.970 0.885 3.090 1.375 ;
        RECT  2.700 1.145 2.970 1.375 ;
        RECT  2.580 1.045 2.700 1.375 ;
        RECT  1.920 1.145 2.580 1.375 ;
        RECT  1.805 1.025 1.920 1.375 ;
        RECT  1.725 1.145 1.805 1.375 ;
        RECT  1.620 1.010 1.725 1.375 ;
        RECT  0.940 1.145 1.620 1.375 ;
        RECT  0.820 1.040 0.940 1.375 ;
        RECT  0.140 1.145 0.820 1.375 ;
        RECT  0.040 0.865 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.875 0.355 2.975 0.465 ;
        RECT  2.875 0.695 2.975 0.815 ;
        RECT  2.805 0.185 2.875 0.465 ;
        RECT  2.805 0.695 2.875 1.035 ;
        RECT  2.725 0.545 2.850 0.615 ;
        RECT  2.655 0.545 2.725 0.925 ;
        RECT  0.905 0.855 2.655 0.925 ;
        RECT  2.380 0.215 2.500 0.425 ;
        RECT  2.000 0.995 2.500 1.065 ;
        RECT  2.095 0.355 2.380 0.425 ;
        RECT  2.025 0.190 2.095 0.425 ;
        RECT  1.040 0.355 2.025 0.425 ;
        RECT  0.130 0.205 1.735 0.275 ;
        RECT  1.040 0.995 1.540 1.065 ;
        RECT  0.835 0.345 0.905 0.925 ;
        RECT  0.220 0.345 0.835 0.415 ;
        RECT  0.410 0.855 0.835 0.925 ;
        RECT  0.220 0.995 0.725 1.065 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA222D4BWP40

MACRO OA22D0BWP40
    CLASS CORE ;
    FOREIGN OA22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.070000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.185 1.365 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.110 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.530 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.115 1.400 0.115 ;
        RECT  0.980 -0.115 1.080 0.275 ;
        RECT  0.340 -0.115 0.980 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.400 1.375 ;
        RECT  0.990 0.980 1.070 1.375 ;
        RECT  0.890 1.145 0.990 1.375 ;
        RECT  0.810 0.980 0.890 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.040 0.940 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.345 1.160 0.905 ;
        RECT  0.600 0.345 1.070 0.415 ;
        RECT  0.705 0.835 1.070 0.905 ;
        RECT  0.510 0.195 0.910 0.265 ;
        RECT  0.635 0.835 0.705 1.045 ;
        RECT  0.410 0.975 0.635 1.045 ;
        RECT  0.430 0.195 0.510 0.415 ;
        RECT  0.035 0.345 0.430 0.415 ;
    END
END OA22D0BWP40

MACRO OA22D1BWP40
    CLASS CORE ;
    FOREIGN OA22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.140000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.185 1.365 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.850 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.115 1.400 0.115 ;
        RECT  0.980 -0.115 1.080 0.275 ;
        RECT  0.340 -0.115 0.980 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.145 1.400 1.375 ;
        RECT  0.990 0.980 1.070 1.375 ;
        RECT  0.890 1.145 0.990 1.375 ;
        RECT  0.810 0.980 0.890 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.040 0.965 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.345 1.160 0.905 ;
        RECT  0.600 0.345 1.070 0.415 ;
        RECT  0.705 0.835 1.070 0.905 ;
        RECT  0.510 0.195 0.910 0.265 ;
        RECT  0.635 0.835 0.705 1.045 ;
        RECT  0.410 0.975 0.635 1.045 ;
        RECT  0.430 0.195 0.510 0.415 ;
        RECT  0.035 0.345 0.430 0.415 ;
    END
END OA22D1BWP40

MACRO OA22D2BWP40
    CLASS CORE ;
    FOREIGN OA22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.132000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 0.495 1.505 0.630 ;
        RECT  1.200 0.185 1.305 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.840 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 -0.115 1.540 0.115 ;
        RECT  1.390 -0.115 1.470 0.410 ;
        RECT  1.080 -0.115 1.390 0.115 ;
        RECT  0.980 -0.115 1.080 0.275 ;
        RECT  0.340 -0.115 0.980 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.145 1.540 1.375 ;
        RECT  1.395 0.720 1.470 1.375 ;
        RECT  1.070 1.145 1.395 1.375 ;
        RECT  0.990 0.980 1.070 1.375 ;
        RECT  0.890 1.145 0.990 1.375 ;
        RECT  0.810 0.980 0.890 1.375 ;
        RECT  0.140 1.145 0.810 1.375 ;
        RECT  0.040 0.855 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.345 1.120 0.905 ;
        RECT  0.600 0.345 1.050 0.415 ;
        RECT  0.705 0.835 1.050 0.905 ;
        RECT  0.510 0.195 0.910 0.265 ;
        RECT  0.635 0.835 0.705 0.990 ;
        RECT  0.410 0.920 0.635 0.990 ;
        RECT  0.430 0.195 0.510 0.415 ;
        RECT  0.125 0.345 0.430 0.415 ;
        RECT  0.055 0.240 0.125 0.415 ;
    END
END OA22D2BWP40

MACRO OA22D4BWP40
    CLASS CORE ;
    FOREIGN OA22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.395 0.465 2.415 0.770 ;
        RECT  2.325 0.185 2.395 1.050 ;
        RECT  2.205 0.355 2.325 0.905 ;
        RECT  2.015 0.355 2.205 0.465 ;
        RECT  2.015 0.770 2.205 0.905 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.770 2.015 1.050 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 0.495 0.805 0.775 ;
        RECT  0.245 0.705 0.705 0.775 ;
        RECT  0.135 0.495 0.245 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.540 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.575 0.775 ;
        RECT  0.960 0.705 1.505 0.775 ;
        RECT  0.875 0.495 0.960 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.495 1.375 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.465 ;
        RECT  2.230 -0.115 2.510 0.115 ;
        RECT  2.110 -0.115 2.230 0.280 ;
        RECT  1.840 -0.115 2.110 0.115 ;
        RECT  1.740 -0.115 1.840 0.275 ;
        RECT  0.700 -0.115 1.740 0.115 ;
        RECT  0.620 -0.115 0.700 0.275 ;
        RECT  0.320 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.320 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.675 2.590 1.375 ;
        RECT  2.230 1.145 2.510 1.375 ;
        RECT  2.110 0.980 2.230 1.375 ;
        RECT  1.840 1.145 2.110 1.375 ;
        RECT  1.740 0.985 1.840 1.375 ;
        RECT  1.660 1.145 1.740 1.375 ;
        RECT  1.565 0.985 1.660 1.375 ;
        RECT  0.905 1.145 1.565 1.375 ;
        RECT  0.805 1.000 0.905 1.375 ;
        RECT  0.140 1.145 0.805 1.375 ;
        RECT  0.040 0.895 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.015 0.355 2.135 0.465 ;
        RECT  2.015 0.770 2.135 0.905 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.945 0.770 2.015 1.050 ;
        RECT  1.715 0.545 2.060 0.615 ;
        RECT  1.645 0.345 1.715 0.915 ;
        RECT  0.885 0.195 1.670 0.265 ;
        RECT  0.980 0.345 1.645 0.415 ;
        RECT  0.410 0.845 1.645 0.915 ;
        RECT  0.980 0.995 1.485 1.065 ;
        RECT  0.815 0.195 0.885 0.415 ;
        RECT  0.520 0.345 0.815 0.415 ;
        RECT  0.220 0.995 0.725 1.065 ;
        RECT  0.420 0.190 0.520 0.415 ;
        RECT  0.130 0.345 0.420 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OA22D4BWP40

MACRO OA31D0BWP40
    CLASS CORE ;
    FOREIGN OA31D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.070000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.195 1.225 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.870 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 -0.115 1.260 0.115 ;
        RECT  0.830 -0.115 0.950 0.135 ;
        RECT  0.000 -0.115 0.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.145 1.260 1.375 ;
        RECT  0.830 1.050 0.950 1.375 ;
        RECT  0.140 1.145 0.830 1.375 ;
        RECT  0.040 0.965 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.205 1.055 0.980 ;
        RECT  0.035 0.205 0.985 0.275 ;
        RECT  0.710 0.910 0.985 0.980 ;
        RECT  0.220 0.345 0.725 0.415 ;
        RECT  0.610 0.910 0.710 1.050 ;
    END
END OA31D0BWP40

MACRO OA31D1BWP40
    CLASS CORE ;
    FOREIGN OA31D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.138250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.195 1.225 1.045 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.870 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.640 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 -0.115 1.260 0.115 ;
        RECT  0.830 -0.115 0.950 0.135 ;
        RECT  0.000 -0.115 0.830 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.145 1.260 1.375 ;
        RECT  0.830 0.995 0.950 1.375 ;
        RECT  0.140 1.145 0.830 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.205 1.055 0.915 ;
        RECT  0.035 0.205 0.985 0.275 ;
        RECT  0.700 0.845 0.985 0.915 ;
        RECT  0.220 0.345 0.725 0.415 ;
        RECT  0.605 0.845 0.700 1.075 ;
    END
END OA31D1BWP40

MACRO OA31D2BWP40
    CLASS CORE ;
    FOREIGN OA31D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.132600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.495 1.365 0.625 ;
        RECT  1.080 0.245 1.150 1.065 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.870 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.275 -0.115 1.345 0.425 ;
        RECT  0.930 -0.115 1.275 0.115 ;
        RECT  0.795 -0.115 0.930 0.130 ;
        RECT  0.000 -0.115 0.795 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.275 0.720 1.345 1.375 ;
        RECT  0.920 1.145 1.275 1.375 ;
        RECT  0.800 1.015 0.920 1.375 ;
        RECT  0.140 1.145 0.800 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 0.200 1.010 0.935 ;
        RECT  0.035 0.200 0.940 0.270 ;
        RECT  0.695 0.845 0.940 0.935 ;
        RECT  0.220 0.340 0.725 0.410 ;
        RECT  0.600 0.845 0.695 1.075 ;
    END
END OA31D2BWP40

MACRO OA31D4BWP40
    CLASS CORE ;
    FOREIGN OA31D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.225 2.395 0.535 ;
        RECT  2.325 0.760 2.395 1.075 ;
        RECT  2.275 0.440 2.325 0.535 ;
        RECT  2.275 0.760 2.325 0.905 ;
        RECT  2.065 0.440 2.275 0.905 ;
        RECT  2.015 0.440 2.065 0.535 ;
        RECT  2.015 0.760 2.065 0.905 ;
        RECT  1.945 0.225 2.015 0.535 ;
        RECT  1.945 0.760 2.015 1.075 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.660 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 0.495 0.805 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.000 0.770 ;
        RECT  0.400 0.700 0.875 0.770 ;
        RECT  0.310 0.490 0.400 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.495 1.225 0.910 ;
        RECT  0.130 0.840 1.115 0.910 ;
        RECT  0.130 0.495 0.235 0.625 ;
        RECT  0.035 0.495 0.130 0.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.485 ;
        RECT  2.230 -0.115 2.510 0.115 ;
        RECT  2.110 -0.115 2.230 0.370 ;
        RECT  1.850 -0.115 2.110 0.115 ;
        RECT  1.750 -0.115 1.850 0.265 ;
        RECT  1.485 -0.115 1.750 0.115 ;
        RECT  1.355 -0.115 1.485 0.140 ;
        RECT  0.000 -0.115 1.355 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.700 2.590 1.375 ;
        RECT  2.230 1.145 2.510 1.375 ;
        RECT  2.110 0.980 2.230 1.375 ;
        RECT  1.825 1.145 2.110 1.375 ;
        RECT  1.755 0.875 1.825 1.375 ;
        RECT  1.645 1.145 1.755 1.375 ;
        RECT  1.575 0.875 1.645 1.375 ;
        RECT  1.295 1.145 1.575 1.375 ;
        RECT  1.165 1.120 1.295 1.375 ;
        RECT  0.145 1.145 1.165 1.375 ;
        RECT  0.040 0.990 0.145 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.225 2.395 0.535 ;
        RECT  2.345 0.760 2.395 1.075 ;
        RECT  1.945 0.225 1.995 0.535 ;
        RECT  1.945 0.760 1.995 1.075 ;
        RECT  1.785 0.350 1.855 0.775 ;
        RECT  0.220 0.350 1.785 0.420 ;
        RECT  1.455 0.705 1.785 0.775 ;
        RECT  0.125 0.210 1.670 0.280 ;
        RECT  1.385 0.705 1.455 1.050 ;
        RECT  0.600 0.980 1.385 1.050 ;
        RECT  0.055 0.210 0.125 0.380 ;
    END
END OA31D4BWP40

MACRO OA32D0BWP40
    CLASS CORE ;
    FOREIGN OA32D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.070000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.215 1.645 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 1.145 1.680 1.375 ;
        RECT  1.285 1.025 1.395 1.375 ;
        RECT  1.175 1.145 1.285 1.375 ;
        RECT  1.065 1.025 1.175 1.375 ;
        RECT  0.140 1.145 1.065 1.375 ;
        RECT  0.040 0.920 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.195 1.440 0.955 ;
        RECT  0.035 0.195 1.350 0.265 ;
        RECT  0.740 0.885 1.350 0.955 ;
        RECT  0.220 0.345 1.180 0.415 ;
        RECT  0.640 0.885 0.740 1.045 ;
    END
END OA32D0BWP40

MACRO OA32D1BWP40
    CLASS CORE ;
    FOREIGN OA32D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.138250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.215 1.645 1.075 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.115 1.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 1.145 1.680 1.375 ;
        RECT  1.285 1.025 1.395 1.375 ;
        RECT  1.175 1.145 1.285 1.375 ;
        RECT  1.065 1.025 1.175 1.375 ;
        RECT  0.140 1.145 1.065 1.375 ;
        RECT  0.040 0.845 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.195 1.440 0.920 ;
        RECT  0.035 0.195 1.350 0.265 ;
        RECT  0.740 0.850 1.350 0.920 ;
        RECT  0.220 0.345 1.180 0.415 ;
        RECT  0.635 0.850 0.740 1.075 ;
    END
END OA32D1BWP40

MACRO OA32D2BWP40
    CLASS CORE ;
    FOREIGN OA32D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.605 0.485 1.690 0.805 ;
        RECT  1.500 0.205 1.605 1.070 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.665 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.225 0.665 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.665 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.945 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.115 1.820 0.115 ;
        RECT  1.690 -0.115 1.760 0.365 ;
        RECT  1.405 -0.115 1.690 0.115 ;
        RECT  1.285 -0.115 1.405 0.255 ;
        RECT  0.980 -0.115 1.285 0.115 ;
        RECT  0.860 -0.115 0.980 0.135 ;
        RECT  0.000 -0.115 0.860 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.145 1.820 1.375 ;
        RECT  1.690 0.890 1.760 1.375 ;
        RECT  1.385 1.145 1.690 1.375 ;
        RECT  1.305 0.945 1.385 1.375 ;
        RECT  1.160 1.145 1.305 1.375 ;
        RECT  1.090 0.945 1.160 1.375 ;
        RECT  0.130 1.145 1.090 1.375 ;
        RECT  0.050 0.810 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.345 1.420 0.865 ;
        RECT  0.125 0.345 1.350 0.415 ;
        RECT  0.750 0.795 1.350 0.865 ;
        RECT  0.230 0.205 1.180 0.275 ;
        RECT  0.650 0.795 0.750 1.050 ;
        RECT  0.055 0.255 0.125 0.415 ;
    END
END OA32D2BWP40

MACRO OA32D4BWP40
    CLASS CORE ;
    FOREIGN OA32D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.185 2.835 0.465 ;
        RECT  2.825 0.695 2.835 1.035 ;
        RECT  2.765 0.185 2.825 1.035 ;
        RECT  2.625 0.355 2.765 0.815 ;
        RECT  2.455 0.355 2.625 0.465 ;
        RECT  2.455 0.695 2.625 0.815 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.695 2.455 1.035 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.495 1.785 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.495 2.075 0.775 ;
        RECT  1.375 0.705 1.855 0.775 ;
        RECT  1.295 0.495 1.375 0.775 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.835 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.495 0.995 0.765 ;
        RECT  0.525 0.695 0.915 0.765 ;
        RECT  0.445 0.495 0.525 0.765 ;
        RECT  0.315 0.495 0.445 0.615 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.225 0.905 ;
        RECT  0.245 0.835 1.125 0.905 ;
        RECT  0.155 0.495 0.245 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 -0.115 3.080 0.115 ;
        RECT  2.950 -0.115 3.030 0.475 ;
        RECT  2.670 -0.115 2.950 0.115 ;
        RECT  2.550 -0.115 2.670 0.280 ;
        RECT  2.280 -0.115 2.550 0.115 ;
        RECT  2.180 -0.115 2.280 0.275 ;
        RECT  1.890 -0.115 2.180 0.115 ;
        RECT  1.770 -0.115 1.890 0.135 ;
        RECT  1.490 -0.115 1.770 0.115 ;
        RECT  1.370 -0.115 1.490 0.135 ;
        RECT  0.000 -0.115 1.370 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.145 3.080 1.375 ;
        RECT  2.950 0.675 3.030 1.375 ;
        RECT  2.670 1.145 2.950 1.375 ;
        RECT  2.550 0.885 2.670 1.375 ;
        RECT  2.270 1.145 2.550 1.375 ;
        RECT  2.150 0.995 2.270 1.375 ;
        RECT  2.080 1.145 2.150 1.375 ;
        RECT  1.960 0.995 2.080 1.375 ;
        RECT  1.290 1.145 1.960 1.375 ;
        RECT  1.170 1.125 1.290 1.375 ;
        RECT  0.140 1.145 1.170 1.375 ;
        RECT  0.040 0.985 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.455 0.355 2.555 0.465 ;
        RECT  2.455 0.695 2.555 0.815 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.385 0.695 2.455 1.035 ;
        RECT  2.295 0.540 2.430 0.620 ;
        RECT  2.225 0.345 2.295 0.915 ;
        RECT  0.220 0.345 2.225 0.415 ;
        RECT  1.685 0.845 2.225 0.915 ;
        RECT  0.130 0.205 2.090 0.275 ;
        RECT  1.575 0.845 1.685 1.055 ;
        RECT  0.600 0.985 1.575 1.055 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA32D4BWP40

MACRO OA33D0BWP40
    CLASS CORE ;
    FOREIGN OA33D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.060000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.295 1.645 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.825 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 -0.115 1.680 0.115 ;
        RECT  1.305 -0.115 1.425 0.235 ;
        RECT  0.930 -0.115 1.305 0.115 ;
        RECT  0.810 -0.115 0.930 0.120 ;
        RECT  0.000 -0.115 0.810 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.145 1.680 1.375 ;
        RECT  1.280 1.045 1.405 1.375 ;
        RECT  0.140 1.145 1.280 1.375 ;
        RECT  0.040 0.945 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.345 1.475 0.975 ;
        RECT  0.035 0.345 1.405 0.415 ;
        RECT  0.710 0.905 1.405 0.975 ;
        RECT  0.220 0.195 1.165 0.265 ;
        RECT  0.605 0.905 0.710 1.045 ;
    END
END OA33D0BWP40

MACRO OA33D1BWP40
    CLASS CORE ;
    FOREIGN OA33D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 0.215 1.645 1.075 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.825 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 -0.115 1.680 0.115 ;
        RECT  1.305 -0.115 1.425 0.265 ;
        RECT  0.930 -0.115 1.305 0.115 ;
        RECT  0.810 -0.115 0.930 0.120 ;
        RECT  0.000 -0.115 0.810 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.145 1.680 1.375 ;
        RECT  1.280 1.045 1.405 1.375 ;
        RECT  0.140 1.145 1.280 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.345 1.475 0.975 ;
        RECT  0.035 0.345 1.405 0.415 ;
        RECT  0.600 0.905 1.405 0.975 ;
        RECT  0.220 0.195 1.165 0.265 ;
    END
END OA33D1BWP40

MACRO OA33D2BWP40
    CLASS CORE ;
    FOREIGN OA33D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 0.470 1.645 0.800 ;
        RECT  1.510 0.210 1.615 1.065 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.835 0.770 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.770 ;
        RECT  0.905 0.545 1.015 0.615 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.265 0.630 ;
        RECT  1.155 0.495 1.225 0.770 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.580 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.770 -0.115 1.820 0.115 ;
        RECT  1.695 -0.115 1.770 0.370 ;
        RECT  1.395 -0.115 1.695 0.115 ;
        RECT  1.275 -0.115 1.395 0.275 ;
        RECT  0.940 -0.115 1.275 0.115 ;
        RECT  0.820 -0.115 0.940 0.135 ;
        RECT  0.000 -0.115 0.820 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 1.145 1.820 1.375 ;
        RECT  1.695 0.925 1.765 1.375 ;
        RECT  1.395 1.145 1.695 1.375 ;
        RECT  1.275 1.050 1.395 1.375 ;
        RECT  0.130 1.145 1.275 1.375 ;
        RECT  0.050 0.860 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.355 0.345 1.425 0.975 ;
        RECT  0.130 0.345 1.355 0.415 ;
        RECT  0.610 0.905 1.355 0.975 ;
        RECT  0.220 0.205 1.150 0.275 ;
        RECT  0.050 0.265 0.130 0.415 ;
    END
END OA33D2BWP40

MACRO OA33D4BWP40
    CLASS CORE ;
    FOREIGN OA33D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.245 0.185 3.255 0.465 ;
        RECT  3.245 0.695 3.255 1.045 ;
        RECT  3.185 0.185 3.245 1.045 ;
        RECT  3.045 0.350 3.185 0.815 ;
        RECT  2.875 0.350 3.045 0.465 ;
        RECT  2.855 0.695 3.045 0.815 ;
        RECT  2.805 0.185 2.875 0.465 ;
        RECT  2.785 0.695 2.855 1.045 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 2.005 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.100 0.495 2.205 0.775 ;
        RECT  1.590 0.705 2.100 0.775 ;
        RECT  1.485 0.495 1.590 0.775 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 0.495 2.485 0.915 ;
        RECT  1.385 0.845 2.370 0.915 ;
        RECT  1.295 0.495 1.385 0.915 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.475 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.010 0.775 ;
        RECT  0.395 0.705 0.875 0.775 ;
        RECT  0.315 0.495 0.395 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.495 1.225 0.915 ;
        RECT  0.245 0.845 1.125 0.915 ;
        RECT  0.175 0.495 0.245 0.915 ;
        RECT  0.130 0.495 0.175 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.475 ;
        RECT  3.090 -0.115 3.370 0.115 ;
        RECT  2.970 -0.115 3.090 0.280 ;
        RECT  2.690 -0.115 2.970 0.115 ;
        RECT  2.610 -0.115 2.690 0.275 ;
        RECT  2.340 -0.115 2.610 0.115 ;
        RECT  2.210 -0.115 2.340 0.135 ;
        RECT  1.930 -0.115 2.210 0.115 ;
        RECT  1.810 -0.115 1.930 0.135 ;
        RECT  1.545 -0.115 1.810 0.115 ;
        RECT  1.415 -0.115 1.545 0.135 ;
        RECT  0.000 -0.115 1.415 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.675 3.450 1.375 ;
        RECT  3.080 1.145 3.370 1.375 ;
        RECT  2.960 0.885 3.080 1.375 ;
        RECT  2.690 1.145 2.960 1.375 ;
        RECT  2.570 1.125 2.690 1.375 ;
        RECT  2.480 1.145 2.570 1.375 ;
        RECT  2.360 1.125 2.480 1.375 ;
        RECT  1.335 1.145 2.360 1.375 ;
        RECT  1.210 1.125 1.335 1.375 ;
        RECT  0.140 1.145 1.210 1.375 ;
        RECT  0.040 0.985 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.875 0.350 2.975 0.465 ;
        RECT  2.855 0.695 2.975 0.815 ;
        RECT  2.805 0.185 2.875 0.465 ;
        RECT  2.785 0.695 2.855 1.045 ;
        RECT  2.705 0.545 2.915 0.615 ;
        RECT  2.635 0.345 2.705 1.055 ;
        RECT  0.230 0.345 2.635 0.415 ;
        RECT  0.640 0.985 2.635 1.055 ;
        RECT  0.130 0.205 2.530 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OA33D4BWP40

MACRO OAI211D0BWP40
    CLASS CORE ;
    FOREIGN OAI211D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.095875 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.895 0.735 1.065 ;
        RECT  0.525 0.895 0.665 0.965 ;
        RECT  0.455 0.345 0.525 0.965 ;
        RECT  0.220 0.345 0.455 0.415 ;
        RECT  0.125 0.895 0.455 0.965 ;
        RECT  0.035 0.895 0.125 1.050 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.695 0.685 0.825 ;
        RECT  0.595 0.330 0.665 0.825 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.820 ;
        RECT  0.295 0.695 0.315 0.820 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.940 0.300 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.840 0.935 0.940 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.045 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.150 0.205 0.550 0.275 ;
        RECT  0.035 0.205 0.150 0.295 ;
    END
END OAI211D0BWP40

MACRO OAI211D1BWP40
    CLASS CORE ;
    FOREIGN OAI211D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.171750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.720 0.735 0.970 ;
        RECT  0.525 0.895 0.665 0.970 ;
        RECT  0.455 0.345 0.525 0.970 ;
        RECT  0.220 0.345 0.455 0.415 ;
        RECT  0.125 0.895 0.455 0.970 ;
        RECT  0.035 0.895 0.125 1.050 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.945 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.330 0.665 0.640 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.820 ;
        RECT  0.295 0.695 0.315 0.820 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 -0.115 0.980 0.115 ;
        RECT  0.840 -0.115 0.940 0.415 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.940 1.145 0.980 1.375 ;
        RECT  0.840 0.775 0.940 1.375 ;
        RECT  0.560 1.145 0.840 1.375 ;
        RECT  0.440 1.045 0.560 1.375 ;
        RECT  0.000 1.145 0.440 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.205 0.550 0.275 ;
        RECT  0.050 0.205 0.130 0.395 ;
    END
END OAI211D1BWP40

MACRO OAI211D2BWP40
    CLASS CORE ;
    FOREIGN OAI211D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.292500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.345 1.540 0.415 ;
        RECT  0.945 0.985 1.350 1.055 ;
        RECT  0.915 0.715 0.945 1.055 ;
        RECT  0.875 0.345 0.915 1.055 ;
        RECT  0.845 0.345 0.875 0.785 ;
        RECT  0.700 0.985 0.875 1.055 ;
        RECT  0.620 0.835 0.700 1.055 ;
        RECT  0.330 0.835 0.620 0.905 ;
        RECT  0.230 0.835 0.330 1.075 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.520 0.765 0.640 ;
        RECT  0.625 0.520 0.695 0.765 ;
        RECT  0.245 0.695 0.625 0.765 ;
        RECT  0.155 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.275 0.495 1.375 0.765 ;
        RECT  1.195 0.495 1.275 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.495 1.585 0.905 ;
        RECT  1.085 0.835 1.505 0.905 ;
        RECT  1.015 0.495 1.085 0.905 ;
        RECT  0.985 0.495 1.015 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.530 -0.115 1.820 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.000 -0.115 0.410 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 1.145 1.820 1.375 ;
        RECT  1.695 0.705 1.765 1.375 ;
        RECT  0.940 1.145 1.695 1.375 ;
        RECT  0.820 1.125 0.940 1.375 ;
        RECT  0.520 1.145 0.820 1.375 ;
        RECT  0.420 0.985 0.520 1.375 ;
        RECT  0.140 1.145 0.420 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.205 1.770 0.455 ;
        RECT  0.700 0.205 1.690 0.275 ;
        RECT  0.630 0.205 0.700 0.415 ;
        RECT  0.130 0.345 0.630 0.415 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OAI211D2BWP40

MACRO OAI211D3BWP40
    CLASS CORE ;
    FOREIGN OAI211D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.484300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.775 2.255 1.045 ;
        RECT  1.845 0.785 2.135 0.855 ;
        RECT  1.775 0.785 1.845 1.050 ;
        RECT  1.465 0.785 1.775 0.855 ;
        RECT  1.395 0.785 1.465 1.050 ;
        RECT  1.085 0.785 1.395 0.855 ;
        RECT  1.085 0.335 1.125 0.415 ;
        RECT  1.015 0.335 1.085 0.855 ;
        RECT  0.215 0.335 1.015 0.415 ;
        RECT  0.145 0.785 1.015 0.855 ;
        RECT  0.035 0.785 0.145 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.965 0.495 2.235 0.705 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.535 0.705 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.095200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.495 0.450 0.705 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.093600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.945 0.705 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.445 -0.115 2.520 0.115 ;
        RECT  2.365 -0.115 2.445 0.420 ;
        RECT  2.045 -0.115 2.365 0.115 ;
        RECT  1.965 -0.115 2.045 0.270 ;
        RECT  0.000 -0.115 1.965 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.145 2.520 1.375 ;
        RECT  2.360 0.745 2.440 1.375 ;
        RECT  2.065 1.145 2.360 1.375 ;
        RECT  1.940 0.935 2.065 1.375 ;
        RECT  1.685 1.145 1.940 1.375 ;
        RECT  1.555 0.935 1.685 1.375 ;
        RECT  1.300 1.145 1.555 1.375 ;
        RECT  1.180 0.935 1.300 1.375 ;
        RECT  0.920 1.145 1.180 1.375 ;
        RECT  0.800 1.125 0.920 1.375 ;
        RECT  0.000 1.145 0.800 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.370 0.340 2.265 0.410 ;
        RECT  0.125 0.195 1.690 0.265 ;
        RECT  0.220 0.985 1.110 1.055 ;
        RECT  0.055 0.195 0.125 0.345 ;
    END
END OAI211D3BWP40

MACRO OAI211D4BWP40
    CLASS CORE ;
    FOREIGN OAI211D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.661000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 0.705 3.250 1.035 ;
        RECT  2.840 0.705 3.170 0.820 ;
        RECT  2.760 0.705 2.840 1.035 ;
        RECT  2.430 0.705 2.760 0.820 ;
        RECT  2.350 0.705 2.430 1.035 ;
        RECT  2.020 0.705 2.350 0.820 ;
        RECT  1.940 0.705 2.020 1.035 ;
        RECT  0.735 0.705 1.940 0.820 ;
        RECT  0.735 0.345 1.670 0.415 ;
        RECT  0.525 0.345 0.735 0.820 ;
        RECT  0.130 0.345 0.525 0.415 ;
        RECT  0.220 0.700 0.525 0.820 ;
        RECT  0.050 0.255 0.130 0.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.495 3.315 0.625 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.495 2.455 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.410 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.495 1.435 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.280 -0.115 3.500 0.115 ;
        RECT  3.140 -0.115 3.280 0.275 ;
        RECT  2.860 -0.115 3.140 0.115 ;
        RECT  2.740 -0.115 2.860 0.275 ;
        RECT  0.000 -0.115 2.740 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 1.145 3.500 1.375 ;
        RECT  3.360 0.705 3.460 1.375 ;
        RECT  3.060 1.145 3.360 1.375 ;
        RECT  2.940 0.890 3.060 1.375 ;
        RECT  2.660 1.145 2.940 1.375 ;
        RECT  2.540 0.890 2.660 1.375 ;
        RECT  2.240 1.145 2.540 1.375 ;
        RECT  2.120 0.890 2.240 1.375 ;
        RECT  1.825 1.145 2.120 1.375 ;
        RECT  1.755 0.895 1.825 1.375 ;
        RECT  1.480 1.145 1.755 1.375 ;
        RECT  1.360 1.030 1.480 1.375 ;
        RECT  1.100 1.145 1.360 1.375 ;
        RECT  0.980 1.030 1.100 1.375 ;
        RECT  0.000 1.145 0.980 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.170 0.705 3.250 1.035 ;
        RECT  2.840 0.705 3.170 0.820 ;
        RECT  2.760 0.705 2.840 1.035 ;
        RECT  2.430 0.705 2.760 0.820 ;
        RECT  2.350 0.705 2.430 1.035 ;
        RECT  2.020 0.705 2.350 0.820 ;
        RECT  1.940 0.705 2.020 1.035 ;
        RECT  0.805 0.705 1.940 0.820 ;
        RECT  0.805 0.345 1.670 0.415 ;
        RECT  0.130 0.345 0.455 0.415 ;
        RECT  0.220 0.700 0.455 0.820 ;
        RECT  0.050 0.255 0.130 0.415 ;
        RECT  3.370 0.255 3.450 0.415 ;
        RECT  3.040 0.345 3.370 0.415 ;
        RECT  2.960 0.185 3.040 0.415 ;
        RECT  2.640 0.345 2.960 0.415 ;
        RECT  2.560 0.185 2.640 0.415 ;
        RECT  1.830 0.345 2.560 0.415 ;
        RECT  0.220 0.205 2.450 0.275 ;
        RECT  1.750 0.345 1.830 0.475 ;
        RECT  0.130 0.890 1.670 0.960 ;
        RECT  0.055 0.735 0.130 1.035 ;
    END
END OAI211D4BWP40

MACRO OAI211D6BWP40
    CLASS CORE ;
    FOREIGN OAI211D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.963500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 0.770 4.820 1.070 ;
        RECT  4.410 0.770 4.700 0.840 ;
        RECT  4.290 0.770 4.410 1.070 ;
        RECT  4.010 0.770 4.290 0.840 ;
        RECT  3.890 0.770 4.010 1.070 ;
        RECT  3.630 0.770 3.890 0.840 ;
        RECT  3.510 0.770 3.630 1.070 ;
        RECT  3.250 0.770 3.510 0.840 ;
        RECT  3.130 0.770 3.250 1.070 ;
        RECT  2.870 0.770 3.130 0.840 ;
        RECT  2.750 0.770 2.870 1.070 ;
        RECT  1.435 0.770 2.750 0.840 ;
        RECT  2.365 0.355 2.475 0.525 ;
        RECT  1.435 0.355 2.365 0.430 ;
        RECT  1.225 0.355 1.435 0.840 ;
        RECT  0.125 0.355 1.225 0.430 ;
        RECT  0.220 0.770 1.225 0.840 ;
        RECT  0.055 0.275 0.125 0.430 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.525 4.790 0.665 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.525 3.225 0.665 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.525 0.855 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.525 2.100 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.800 -0.115 5.040 0.115 ;
        RECT  4.720 -0.115 4.800 0.280 ;
        RECT  4.390 -0.115 4.720 0.115 ;
        RECT  4.310 -0.115 4.390 0.280 ;
        RECT  3.990 -0.115 4.310 0.115 ;
        RECT  3.910 -0.115 3.990 0.280 ;
        RECT  0.000 -0.115 3.910 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.720 4.990 1.375 ;
        RECT  4.620 1.145 4.910 1.375 ;
        RECT  4.500 0.910 4.620 1.375 ;
        RECT  4.210 1.145 4.500 1.375 ;
        RECT  4.090 0.910 4.210 1.375 ;
        RECT  3.820 1.145 4.090 1.375 ;
        RECT  3.700 0.910 3.820 1.375 ;
        RECT  3.440 1.145 3.700 1.375 ;
        RECT  3.320 0.910 3.440 1.375 ;
        RECT  3.060 1.145 3.320 1.375 ;
        RECT  2.940 0.910 3.060 1.375 ;
        RECT  2.660 1.145 2.940 1.375 ;
        RECT  2.580 0.985 2.660 1.375 ;
        RECT  2.280 1.145 2.580 1.375 ;
        RECT  2.160 1.050 2.280 1.375 ;
        RECT  1.880 1.145 2.160 1.375 ;
        RECT  1.760 1.050 1.880 1.375 ;
        RECT  1.495 1.145 1.760 1.375 ;
        RECT  1.365 1.050 1.495 1.375 ;
        RECT  0.000 1.145 1.365 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.700 0.770 4.820 1.070 ;
        RECT  4.410 0.770 4.700 0.840 ;
        RECT  4.290 0.770 4.410 1.070 ;
        RECT  4.010 0.770 4.290 0.840 ;
        RECT  3.890 0.770 4.010 1.070 ;
        RECT  3.630 0.770 3.890 0.840 ;
        RECT  3.510 0.770 3.630 1.070 ;
        RECT  3.250 0.770 3.510 0.840 ;
        RECT  3.130 0.770 3.250 1.070 ;
        RECT  2.870 0.770 3.130 0.840 ;
        RECT  2.750 0.770 2.870 1.070 ;
        RECT  1.505 0.770 2.750 0.840 ;
        RECT  2.365 0.355 2.475 0.525 ;
        RECT  1.505 0.355 2.365 0.430 ;
        RECT  0.125 0.355 1.155 0.430 ;
        RECT  0.220 0.770 1.155 0.840 ;
        RECT  0.055 0.275 0.125 0.430 ;
        RECT  2.560 0.360 5.005 0.430 ;
        RECT  0.220 0.195 3.635 0.265 ;
        RECT  0.130 0.910 2.480 0.980 ;
        RECT  0.050 0.815 0.130 0.980 ;
    END
END OAI211D6BWP40

MACRO OAI211D8BWP40
    CLASS CORE ;
    FOREIGN OAI211D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.271000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.240 0.770 6.360 1.070 ;
        RECT  5.950 0.770 6.240 0.840 ;
        RECT  5.830 0.770 5.950 1.070 ;
        RECT  5.550 0.770 5.830 0.840 ;
        RECT  5.430 0.770 5.550 1.070 ;
        RECT  5.150 0.770 5.430 0.840 ;
        RECT  5.035 0.770 5.150 1.070 ;
        RECT  4.770 0.770 5.035 0.840 ;
        RECT  4.650 0.770 4.770 1.070 ;
        RECT  4.390 0.770 4.650 0.840 ;
        RECT  4.270 0.770 4.390 1.070 ;
        RECT  4.010 0.770 4.270 0.840 ;
        RECT  3.890 0.770 4.010 1.070 ;
        RECT  3.630 0.770 3.890 0.840 ;
        RECT  3.510 0.770 3.630 1.070 ;
        RECT  1.575 0.770 3.510 0.840 ;
        RECT  1.575 0.355 3.240 0.430 ;
        RECT  1.365 0.355 1.575 0.840 ;
        RECT  0.125 0.355 1.365 0.425 ;
        RECT  0.220 0.770 1.365 0.840 ;
        RECT  0.055 0.285 0.125 0.425 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.755 0.525 6.330 0.665 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.525 3.985 0.665 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.495 0.855 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.525 2.965 0.665 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.340 -0.115 6.580 0.115 ;
        RECT  6.260 -0.115 6.340 0.275 ;
        RECT  5.930 -0.115 6.260 0.115 ;
        RECT  5.850 -0.115 5.930 0.275 ;
        RECT  5.530 -0.115 5.850 0.115 ;
        RECT  5.450 -0.115 5.530 0.275 ;
        RECT  5.130 -0.115 5.450 0.115 ;
        RECT  5.050 -0.115 5.130 0.275 ;
        RECT  0.000 -0.115 5.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.580 1.375 ;
        RECT  6.450 0.720 6.530 1.375 ;
        RECT  6.160 1.145 6.450 1.375 ;
        RECT  6.040 0.910 6.160 1.375 ;
        RECT  5.750 1.145 6.040 1.375 ;
        RECT  5.630 0.910 5.750 1.375 ;
        RECT  5.350 1.145 5.630 1.375 ;
        RECT  5.230 0.910 5.350 1.375 ;
        RECT  4.960 1.145 5.230 1.375 ;
        RECT  4.840 0.910 4.960 1.375 ;
        RECT  4.580 1.145 4.840 1.375 ;
        RECT  4.460 0.910 4.580 1.375 ;
        RECT  4.200 1.145 4.460 1.375 ;
        RECT  4.080 0.910 4.200 1.375 ;
        RECT  3.820 1.145 4.080 1.375 ;
        RECT  3.700 0.910 3.820 1.375 ;
        RECT  3.420 1.145 3.700 1.375 ;
        RECT  3.340 0.985 3.420 1.375 ;
        RECT  3.040 1.145 3.340 1.375 ;
        RECT  2.920 1.050 3.040 1.375 ;
        RECT  2.640 1.145 2.920 1.375 ;
        RECT  2.520 1.050 2.640 1.375 ;
        RECT  2.255 1.145 2.520 1.375 ;
        RECT  2.125 1.050 2.255 1.375 ;
        RECT  1.875 1.145 2.125 1.375 ;
        RECT  1.745 1.050 1.875 1.375 ;
        RECT  0.000 1.145 1.745 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.240 0.770 6.360 1.070 ;
        RECT  5.950 0.770 6.240 0.840 ;
        RECT  5.830 0.770 5.950 1.070 ;
        RECT  5.550 0.770 5.830 0.840 ;
        RECT  5.430 0.770 5.550 1.070 ;
        RECT  5.150 0.770 5.430 0.840 ;
        RECT  5.035 0.770 5.150 1.070 ;
        RECT  4.770 0.770 5.035 0.840 ;
        RECT  4.650 0.770 4.770 1.070 ;
        RECT  4.390 0.770 4.650 0.840 ;
        RECT  4.270 0.770 4.390 1.070 ;
        RECT  4.010 0.770 4.270 0.840 ;
        RECT  3.890 0.770 4.010 1.070 ;
        RECT  3.630 0.770 3.890 0.840 ;
        RECT  3.510 0.770 3.630 1.070 ;
        RECT  1.645 0.770 3.510 0.840 ;
        RECT  1.645 0.355 3.240 0.430 ;
        RECT  0.125 0.355 1.295 0.425 ;
        RECT  0.220 0.770 1.295 0.840 ;
        RECT  0.055 0.285 0.125 0.425 ;
        RECT  3.320 0.360 6.545 0.430 ;
        RECT  0.220 0.195 4.780 0.265 ;
        RECT  0.130 0.910 3.240 0.980 ;
        RECT  0.050 0.815 0.130 0.980 ;
    END
END OAI211D8BWP40

MACRO OAI21D0BWP40
    CLASS CORE ;
    FOREIGN OAI21D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.078625 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.345 0.525 1.065 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.115 0.840 0.115 ;
        RECT  0.675 -0.115 0.745 0.275 ;
        RECT  0.000 -0.115 0.675 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.650 0.925 0.740 1.375 ;
        RECT  0.140 1.145 0.650 1.375 ;
        RECT  0.040 0.960 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.140 0.205 0.565 0.275 ;
        RECT  0.040 0.185 0.140 0.285 ;
    END
END OAI21D0BWP40

MACRO OAI21D1BWP40
    CLASS CORE ;
    FOREIGN OAI21D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.134750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.745 0.545 1.075 ;
        RECT  0.455 0.345 0.525 1.075 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.745 -0.115 0.840 0.115 ;
        RECT  0.675 -0.115 0.745 0.415 ;
        RECT  0.000 -0.115 0.675 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.840 1.375 ;
        RECT  0.665 0.855 0.740 1.375 ;
        RECT  0.140 1.145 0.665 1.375 ;
        RECT  0.040 0.850 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.205 0.565 0.275 ;
        RECT  0.050 0.205 0.130 0.375 ;
    END
END OAI21D1BWP40

MACRO OAI21D2BWP40
    CLASS CORE ;
    FOREIGN OAI21D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.300000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.845 1.365 1.065 ;
        RECT  0.410 0.845 1.240 0.915 ;
        RECT  0.410 0.345 1.100 0.415 ;
        RECT  0.315 0.345 0.410 0.915 ;
        RECT  0.125 0.845 0.315 0.915 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.765 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.495 1.085 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.280 0.765 ;
        RECT  0.750 0.695 1.155 0.765 ;
        RECT  0.680 0.495 0.750 0.765 ;
        RECT  0.550 0.495 0.680 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 1.400 0.115 ;
        RECT  0.220 -0.115 0.340 0.130 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.145 1.400 1.375 ;
        RECT  0.785 1.050 0.915 1.375 ;
        RECT  0.340 1.145 0.785 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.270 0.205 1.340 0.345 ;
        RECT  0.130 0.205 1.270 0.275 ;
        RECT  0.055 0.205 0.130 0.390 ;
    END
END OAI21D2BWP40

MACRO OAI21D3BWP40
    CLASS CORE ;
    FOREIGN OAI21D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.725 1.680 0.800 ;
        RECT  0.665 0.335 1.105 0.415 ;
        RECT  0.595 0.335 0.665 0.800 ;
        RECT  0.215 0.335 0.595 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.475 0.495 1.845 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.135 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 0.495 1.225 0.645 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 -0.115 1.960 0.115 ;
        RECT  1.800 -0.115 1.880 0.415 ;
        RECT  1.485 -0.115 1.800 0.115 ;
        RECT  1.355 -0.115 1.485 0.210 ;
        RECT  0.000 -0.115 1.355 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.145 1.960 1.375 ;
        RECT  1.800 0.715 1.880 1.375 ;
        RECT  1.465 1.145 1.800 1.375 ;
        RECT  1.380 0.870 1.465 1.375 ;
        RECT  0.530 1.145 1.380 1.375 ;
        RECT  0.410 1.050 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.715 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.265 0.300 1.675 0.370 ;
        RECT  1.195 0.195 1.265 0.370 ;
        RECT  0.125 0.195 1.195 0.265 ;
        RECT  0.215 0.900 1.130 0.970 ;
        RECT  0.055 0.195 0.125 0.365 ;
    END
END OAI21D3BWP40

MACRO OAI21D4BWP40
    CLASS CORE ;
    FOREIGN OAI21D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.508000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 0.705 2.420 1.060 ;
        RECT  1.645 0.705 2.300 0.775 ;
        RECT  1.575 0.355 1.645 0.775 ;
        RECT  0.735 0.355 1.575 0.425 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.035 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.495 2.315 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.885 0.495 1.440 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.435 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 -0.115 2.660 0.115 ;
        RECT  2.510 -0.115 2.590 0.425 ;
        RECT  2.210 -0.115 2.510 0.115 ;
        RECT  2.130 -0.115 2.210 0.270 ;
        RECT  1.850 -0.115 2.130 0.115 ;
        RECT  1.730 -0.115 1.850 0.130 ;
        RECT  0.000 -0.115 1.730 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.710 2.590 1.375 ;
        RECT  2.210 1.145 2.510 1.375 ;
        RECT  2.130 0.855 2.210 1.375 ;
        RECT  1.840 1.145 2.130 1.375 ;
        RECT  1.740 0.855 1.840 1.375 ;
        RECT  1.460 1.145 1.740 1.375 ;
        RECT  1.380 0.995 1.460 1.375 ;
        RECT  1.075 1.145 1.380 1.375 ;
        RECT  1.005 0.995 1.075 1.375 ;
        RECT  0.000 1.145 1.005 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.705 2.300 0.775 ;
        RECT  1.575 0.355 1.645 0.775 ;
        RECT  0.805 0.355 1.575 0.425 ;
        RECT  0.035 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  2.305 0.300 2.420 0.420 ;
        RECT  2.015 0.350 2.305 0.420 ;
        RECT  1.945 0.215 2.015 0.420 ;
        RECT  0.220 0.215 1.945 0.285 ;
        RECT  1.570 0.845 1.650 0.970 ;
        RECT  1.290 0.845 1.570 0.915 ;
        RECT  1.170 0.845 1.290 1.055 ;
        RECT  0.925 0.845 1.170 0.915 ;
        RECT  0.855 0.845 0.925 1.055 ;
        RECT  0.130 0.980 0.855 1.055 ;
        RECT  0.050 0.785 0.130 1.055 ;
        RECT  2.300 0.705 2.420 1.060 ;
    END
END OAI21D4BWP40

MACRO OAI21D6BWP40
    CLASS CORE ;
    FOREIGN OAI21D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.748000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.705 3.560 1.060 ;
        RECT  3.155 0.705 3.440 0.775 ;
        RECT  3.085 0.705 3.155 0.990 ;
        RECT  2.775 0.705 3.085 0.775 ;
        RECT  2.705 0.705 2.775 0.990 ;
        RECT  2.405 0.705 2.705 0.775 ;
        RECT  2.335 0.355 2.405 0.775 ;
        RECT  0.735 0.355 2.335 0.425 ;
        RECT  0.735 0.840 1.115 0.910 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.035 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.085 0.495 3.455 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.495 2.200 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.435 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 -0.115 3.780 0.115 ;
        RECT  3.650 -0.115 3.730 0.420 ;
        RECT  3.350 -0.115 3.650 0.115 ;
        RECT  3.270 -0.115 3.350 0.260 ;
        RECT  2.970 -0.115 3.270 0.115 ;
        RECT  2.900 -0.115 2.970 0.280 ;
        RECT  2.610 -0.115 2.900 0.115 ;
        RECT  2.490 -0.115 2.610 0.130 ;
        RECT  0.000 -0.115 2.490 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.145 3.780 1.375 ;
        RECT  3.650 0.720 3.730 1.375 ;
        RECT  3.360 1.145 3.650 1.375 ;
        RECT  3.260 0.870 3.360 1.375 ;
        RECT  2.980 1.145 3.260 1.375 ;
        RECT  2.880 0.870 2.980 1.375 ;
        RECT  2.600 1.145 2.880 1.375 ;
        RECT  2.500 0.870 2.600 1.375 ;
        RECT  2.220 1.145 2.500 1.375 ;
        RECT  2.140 0.995 2.220 1.375 ;
        RECT  1.835 1.145 2.140 1.375 ;
        RECT  1.765 0.995 1.835 1.375 ;
        RECT  1.455 1.145 1.765 1.375 ;
        RECT  1.385 0.995 1.455 1.375 ;
        RECT  0.000 1.145 1.385 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.440 0.705 3.560 1.060 ;
        RECT  3.155 0.705 3.440 0.775 ;
        RECT  3.085 0.705 3.155 0.990 ;
        RECT  2.775 0.705 3.085 0.775 ;
        RECT  2.705 0.705 2.775 0.990 ;
        RECT  2.405 0.705 2.705 0.775 ;
        RECT  2.335 0.355 2.405 0.775 ;
        RECT  0.805 0.355 2.335 0.425 ;
        RECT  0.805 0.840 1.115 0.910 ;
        RECT  0.035 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  2.330 0.845 2.410 0.970 ;
        RECT  2.050 0.845 2.330 0.915 ;
        RECT  1.930 0.845 2.050 1.055 ;
        RECT  1.670 0.845 1.930 0.915 ;
        RECT  1.550 0.845 1.670 1.055 ;
        RECT  1.305 0.845 1.550 0.915 ;
        RECT  1.235 0.845 1.305 1.055 ;
        RECT  0.130 0.980 1.235 1.055 ;
        RECT  0.050 0.770 0.130 1.055 ;
        RECT  3.450 0.285 3.560 0.420 ;
        RECT  2.775 0.350 3.450 0.420 ;
        RECT  2.705 0.215 2.775 0.420 ;
        RECT  0.220 0.215 2.705 0.285 ;
    END
END OAI21D6BWP40

MACRO OAI21D8BWP40
    CLASS CORE ;
    FOREIGN OAI21D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.008250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 0.705 4.820 1.060 ;
        RECT  4.420 0.705 4.700 0.775 ;
        RECT  4.345 0.705 4.420 0.990 ;
        RECT  4.035 0.705 4.345 0.775 ;
        RECT  3.965 0.705 4.035 0.990 ;
        RECT  3.625 0.705 3.965 0.775 ;
        RECT  3.555 0.705 3.625 0.990 ;
        RECT  3.165 0.705 3.555 0.775 ;
        RECT  3.095 0.355 3.165 0.775 ;
        RECT  1.015 0.355 3.095 0.425 ;
        RECT  1.015 0.840 1.505 0.910 ;
        RECT  0.805 0.355 1.015 0.910 ;
        RECT  0.035 0.355 0.805 0.425 ;
        RECT  0.220 0.840 0.805 0.910 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.254400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.345 0.495 4.715 0.625 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.495 2.960 0.625 ;
        RECT  2.415 0.495 2.485 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.250 0.495 0.455 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.910 -0.115 4.990 0.380 ;
        RECT  4.610 -0.115 4.910 0.115 ;
        RECT  4.530 -0.115 4.610 0.260 ;
        RECT  4.230 -0.115 4.530 0.115 ;
        RECT  4.160 -0.115 4.230 0.280 ;
        RECT  3.845 -0.115 4.160 0.115 ;
        RECT  3.775 -0.115 3.845 0.280 ;
        RECT  3.405 -0.115 3.775 0.115 ;
        RECT  3.260 -0.115 3.405 0.130 ;
        RECT  0.000 -0.115 3.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.910 0.720 4.990 1.375 ;
        RECT  4.620 1.145 4.910 1.375 ;
        RECT  4.520 0.870 4.620 1.375 ;
        RECT  4.240 1.145 4.520 1.375 ;
        RECT  4.140 0.870 4.240 1.375 ;
        RECT  3.860 1.145 4.140 1.375 ;
        RECT  3.760 0.870 3.860 1.375 ;
        RECT  3.415 1.145 3.760 1.375 ;
        RECT  3.315 0.870 3.415 1.375 ;
        RECT  2.980 1.145 3.315 1.375 ;
        RECT  2.900 0.995 2.980 1.375 ;
        RECT  2.595 1.145 2.900 1.375 ;
        RECT  2.525 0.995 2.595 1.375 ;
        RECT  2.215 1.145 2.525 1.375 ;
        RECT  2.145 0.995 2.215 1.375 ;
        RECT  1.835 1.145 2.145 1.375 ;
        RECT  1.765 0.995 1.835 1.375 ;
        RECT  0.000 1.145 1.765 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.700 0.705 4.820 1.060 ;
        RECT  4.420 0.705 4.700 0.775 ;
        RECT  4.345 0.705 4.420 0.990 ;
        RECT  4.035 0.705 4.345 0.775 ;
        RECT  3.965 0.705 4.035 0.990 ;
        RECT  3.625 0.705 3.965 0.775 ;
        RECT  3.555 0.705 3.625 0.990 ;
        RECT  3.165 0.705 3.555 0.775 ;
        RECT  3.095 0.355 3.165 0.775 ;
        RECT  1.085 0.355 3.095 0.425 ;
        RECT  1.085 0.840 1.505 0.910 ;
        RECT  0.035 0.355 0.735 0.425 ;
        RECT  0.220 0.840 0.735 0.910 ;
        RECT  3.620 0.350 4.820 0.420 ;
        RECT  3.550 0.215 3.620 0.420 ;
        RECT  0.220 0.215 3.550 0.285 ;
        RECT  3.090 0.845 3.170 0.970 ;
        RECT  2.810 0.845 3.090 0.915 ;
        RECT  2.690 0.845 2.810 1.055 ;
        RECT  2.430 0.845 2.690 0.915 ;
        RECT  2.310 0.845 2.430 1.055 ;
        RECT  1.930 0.845 2.050 1.055 ;
        RECT  1.685 0.845 1.930 0.915 ;
        RECT  1.615 0.845 1.685 1.055 ;
        RECT  0.130 0.980 1.615 1.055 ;
        RECT  0.050 0.755 0.130 1.055 ;
        RECT  2.050 0.845 2.310 0.915 ;
    END
END OAI21D8BWP40

MACRO OAI221D0BWP40
    CLASS CORE ;
    FOREIGN OAI221D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.118825 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.835 1.150 1.075 ;
        RECT  0.385 0.835 1.050 0.905 ;
        RECT  0.285 0.340 0.385 0.905 ;
        RECT  0.140 0.835 0.285 0.905 ;
        RECT  0.035 0.835 0.140 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.295 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.840 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.495 0.210 0.630 ;
        RECT  0.035 0.495 0.140 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.285 ;
        RECT  0.000 -0.115 1.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.945 1.360 1.375 ;
        RECT  0.770 1.145 1.260 1.375 ;
        RECT  0.670 0.975 0.770 1.375 ;
        RECT  0.590 1.145 0.670 1.375 ;
        RECT  0.490 0.975 0.590 1.375 ;
        RECT  0.000 1.145 0.490 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.185 1.150 0.425 ;
        RECT  0.660 0.355 1.050 0.425 ;
        RECT  0.140 0.195 0.970 0.265 ;
        RECT  0.040 0.195 0.140 0.300 ;
    END
END OAI221D0BWP40

MACRO OAI221D1BWP40
    CLASS CORE ;
    FOREIGN OAI221D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.205250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.835 1.150 1.075 ;
        RECT  0.385 0.835 1.050 0.905 ;
        RECT  0.285 0.340 0.385 0.905 ;
        RECT  0.140 0.835 0.285 0.905 ;
        RECT  0.035 0.835 0.140 1.075 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.295 0.625 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.495 1.085 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.840 0.765 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.665 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.495 0.210 0.630 ;
        RECT  0.035 0.495 0.140 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.425 ;
        RECT  0.000 -0.115 1.260 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.850 1.360 1.375 ;
        RECT  0.770 1.145 1.260 1.375 ;
        RECT  0.670 0.975 0.770 1.375 ;
        RECT  0.590 1.145 0.670 1.375 ;
        RECT  0.490 0.975 0.590 1.375 ;
        RECT  0.000 1.145 0.490 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.185 1.150 0.425 ;
        RECT  0.660 0.355 1.050 0.425 ;
        RECT  0.140 0.195 0.970 0.265 ;
        RECT  0.040 0.195 0.140 0.345 ;
    END
END OAI221D1BWP40

MACRO OAI221D2BWP40
    CLASS CORE ;
    FOREIGN OAI221D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.398500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.845 2.120 1.070 ;
        RECT  0.125 0.845 1.995 0.915 ;
        RECT  0.130 0.345 0.925 0.415 ;
        RECT  0.105 0.215 0.130 0.415 ;
        RECT  0.105 0.845 0.125 1.045 ;
        RECT  0.035 0.215 0.105 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.135 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.645 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.835 0.775 ;
        RECT  1.240 0.705 1.715 0.775 ;
        RECT  1.165 0.495 1.240 0.775 ;
        RECT  1.100 0.495 1.165 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.695 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.765 0.495 0.845 0.775 ;
        RECT  0.255 0.705 0.765 0.775 ;
        RECT  0.175 0.495 0.255 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.105 -0.115 2.380 0.115 ;
        RECT  2.025 -0.115 2.105 0.260 ;
        RECT  0.000 -0.115 2.025 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 1.145 2.380 1.375 ;
        RECT  2.235 0.720 2.315 1.375 ;
        RECT  1.845 1.145 2.235 1.375 ;
        RECT  1.775 0.995 1.845 1.375 ;
        RECT  1.110 1.145 1.775 1.375 ;
        RECT  0.990 0.985 1.110 1.375 ;
        RECT  0.550 1.145 0.990 1.375 ;
        RECT  0.430 1.040 0.550 1.375 ;
        RECT  0.000 1.145 0.430 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.225 0.245 2.325 0.415 ;
        RECT  0.995 0.345 2.225 0.415 ;
        RECT  0.220 0.195 1.680 0.265 ;
        RECT  1.180 0.995 1.680 1.065 ;
    END
END OAI221D2BWP40

MACRO OAI221D4BWP40
    CLASS CORE ;
    FOREIGN OAI221D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.670700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.835 3.970 0.905 ;
        RECT  1.575 0.345 1.670 0.415 ;
        RECT  1.365 0.345 1.575 0.905 ;
        RECT  0.130 0.345 1.365 0.415 ;
        RECT  0.125 0.835 1.365 0.905 ;
        RECT  0.035 0.215 0.130 0.415 ;
        RECT  0.035 0.835 0.125 1.045 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.495 3.745 0.765 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 0.495 2.870 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.220 0.495 3.340 0.765 ;
        RECT  2.135 0.695 3.220 0.765 ;
        RECT  2.060 0.535 2.135 0.765 ;
        RECT  1.995 0.535 2.060 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.495 0.855 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.245 0.765 ;
        RECT  0.255 0.695 1.155 0.765 ;
        RECT  0.175 0.495 0.255 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 -0.115 4.200 0.115 ;
        RECT  3.870 -0.115 3.950 0.260 ;
        RECT  3.570 -0.115 3.870 0.115 ;
        RECT  3.490 -0.115 3.570 0.260 ;
        RECT  0.000 -0.115 3.490 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.140 1.145 4.200 1.375 ;
        RECT  4.060 0.720 4.140 1.375 ;
        RECT  3.760 1.145 4.060 1.375 ;
        RECT  3.680 0.980 3.760 1.375 ;
        RECT  3.350 1.145 3.680 1.375 ;
        RECT  3.280 1.000 3.350 1.375 ;
        RECT  2.235 1.145 3.280 1.375 ;
        RECT  2.105 1.120 2.235 1.375 ;
        RECT  1.845 1.145 2.105 1.375 ;
        RECT  1.730 0.985 1.845 1.375 ;
        RECT  0.910 1.145 1.730 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 1.120 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.835 3.970 0.905 ;
        RECT  1.645 0.345 1.670 0.415 ;
        RECT  0.130 0.345 1.295 0.415 ;
        RECT  0.125 0.835 1.295 0.905 ;
        RECT  0.035 0.215 0.130 0.415 ;
        RECT  0.035 0.835 0.125 1.045 ;
        RECT  1.825 0.345 4.155 0.415 ;
        RECT  1.925 0.975 3.200 1.045 ;
        RECT  0.220 0.205 3.185 0.275 ;
        RECT  1.755 0.345 1.825 0.485 ;
        RECT  0.220 0.975 1.505 1.045 ;
    END
END OAI221D4BWP40

MACRO OAI222D0BWP40
    CLASS CORE ;
    FOREIGN OAI222D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.100375 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.870 1.115 1.075 ;
        RECT  0.525 0.870 1.035 0.940 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.225 0.625 ;
        RECT  1.015 0.495 1.085 0.765 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 1.505 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.485 0.685 0.795 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.775 0.495 0.875 0.645 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.275 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.020 -0.115 1.120 0.275 ;
        RECT  0.000 -0.115 1.020 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.985 1.500 1.375 ;
        RECT  0.950 1.145 1.400 1.375 ;
        RECT  0.830 1.010 0.950 1.375 ;
        RECT  0.140 1.145 0.830 1.375 ;
        RECT  0.040 0.975 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.205 1.320 0.415 ;
        RECT  0.620 0.345 1.200 0.415 ;
        RECT  0.130 0.195 0.945 0.265 ;
        RECT  0.050 0.195 0.130 0.325 ;
    END
END OAI222D0BWP40

MACRO OAI222D1BWP40
    CLASS CORE ;
    FOREIGN OAI222D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.180750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.870 1.115 1.075 ;
        RECT  0.525 0.870 1.035 0.940 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.220 0.345 0.455 0.415 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.155 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.765 ;
        RECT  1.295 0.495 1.435 0.625 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.485 0.685 0.795 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.775 0.495 0.875 0.645 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 -0.115 1.540 0.115 ;
        RECT  1.400 -0.115 1.500 0.360 ;
        RECT  1.120 -0.115 1.400 0.115 ;
        RECT  1.020 -0.115 1.120 0.275 ;
        RECT  0.000 -0.115 1.020 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.145 1.540 1.375 ;
        RECT  1.400 0.845 1.500 1.375 ;
        RECT  0.950 1.145 1.400 1.375 ;
        RECT  0.830 1.010 0.950 1.375 ;
        RECT  0.140 1.145 0.830 1.375 ;
        RECT  0.040 0.870 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 0.205 1.320 0.415 ;
        RECT  0.620 0.345 1.200 0.415 ;
        RECT  0.130 0.195 0.945 0.265 ;
        RECT  0.050 0.195 0.130 0.395 ;
    END
END OAI222D1BWP40

MACRO OAI222D2BWP40
    CLASS CORE ;
    FOREIGN OAI222D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.371500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.845 2.230 0.915 ;
        RECT  0.905 0.485 0.945 0.915 ;
        RECT  0.875 0.345 0.905 0.915 ;
        RECT  0.835 0.345 0.875 0.555 ;
        RECT  0.125 0.845 0.875 0.915 ;
        RECT  0.130 0.345 0.835 0.415 ;
        RECT  0.035 0.215 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.485 2.235 0.625 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.495 2.510 0.765 ;
        RECT  1.925 0.695 2.385 0.765 ;
        RECT  1.845 0.495 1.925 0.765 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.495 1.505 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.705 0.775 ;
        RECT  1.175 0.705 1.575 0.775 ;
        RECT  1.105 0.510 1.175 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.765 0.695 0.805 0.765 ;
        RECT  0.695 0.500 0.765 0.765 ;
        RECT  0.245 0.695 0.695 0.765 ;
        RECT  0.170 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.115 2.660 0.115 ;
        RECT  2.320 -0.115 2.400 0.275 ;
        RECT  2.020 -0.115 2.320 0.115 ;
        RECT  1.940 -0.115 2.020 0.275 ;
        RECT  0.000 -0.115 1.940 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 2.660 1.375 ;
        RECT  2.510 0.840 2.590 1.375 ;
        RECT  1.825 1.145 2.510 1.375 ;
        RECT  1.755 0.985 1.825 1.375 ;
        RECT  1.090 1.145 1.755 1.375 ;
        RECT  0.970 0.985 1.090 1.375 ;
        RECT  0.530 1.145 0.970 1.375 ;
        RECT  0.410 1.040 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.510 0.255 2.590 0.415 ;
        RECT  2.230 0.345 2.510 0.415 ;
        RECT  1.920 0.995 2.420 1.065 ;
        RECT  2.110 0.205 2.230 0.415 ;
        RECT  1.840 0.345 2.110 0.415 ;
        RECT  1.740 0.190 1.840 0.415 ;
        RECT  0.975 0.345 1.740 0.415 ;
        RECT  0.220 0.195 1.660 0.265 ;
        RECT  1.160 0.995 1.660 1.065 ;
    END
END OAI222D2BWP40

MACRO OAI222D4BWP40
    CLASS CORE ;
    FOREIGN OAI222D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.672850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.845 4.610 0.915 ;
        RECT  1.575 0.345 1.650 0.475 ;
        RECT  1.365 0.345 1.575 0.915 ;
        RECT  0.130 0.345 1.365 0.415 ;
        RECT  0.125 0.845 1.365 0.915 ;
        RECT  0.035 0.215 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.045 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.495 4.585 0.630 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.765 0.495 4.890 0.775 ;
        RECT  3.620 0.705 4.765 0.775 ;
        RECT  3.530 0.495 3.620 0.775 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.127200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.495 3.045 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.125600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.250 0.775 ;
        RECT  2.090 0.705 3.115 0.775 ;
        RECT  1.975 0.495 2.090 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.730 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.545 1.235 0.615 ;
        RECT  1.015 0.545 1.130 0.775 ;
        RECT  0.245 0.705 1.015 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.780 -0.115 5.040 0.115 ;
        RECT  4.700 -0.115 4.780 0.275 ;
        RECT  4.400 -0.115 4.700 0.115 ;
        RECT  4.320 -0.115 4.400 0.275 ;
        RECT  3.960 -0.115 4.320 0.115 ;
        RECT  3.870 -0.115 3.960 0.275 ;
        RECT  3.560 -0.115 3.870 0.115 ;
        RECT  3.445 -0.115 3.560 0.275 ;
        RECT  0.000 -0.115 3.445 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 1.145 5.040 1.375 ;
        RECT  4.890 0.860 4.970 1.375 ;
        RECT  3.750 1.145 4.890 1.375 ;
        RECT  3.625 1.125 3.750 1.375 ;
        RECT  3.345 1.145 3.625 1.375 ;
        RECT  3.275 0.985 3.345 1.375 ;
        RECT  2.235 1.145 3.275 1.375 ;
        RECT  2.105 1.125 2.235 1.375 ;
        RECT  1.845 1.145 2.105 1.375 ;
        RECT  1.730 0.985 1.845 1.375 ;
        RECT  0.915 1.145 1.730 1.375 ;
        RECT  0.785 1.125 0.915 1.375 ;
        RECT  0.530 1.145 0.785 1.375 ;
        RECT  0.410 1.125 0.530 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.645 0.845 4.610 0.915 ;
        RECT  1.645 0.345 1.650 0.475 ;
        RECT  0.130 0.345 1.295 0.415 ;
        RECT  0.125 0.845 1.295 0.915 ;
        RECT  0.035 0.215 0.130 0.415 ;
        RECT  0.035 0.845 0.125 1.045 ;
        RECT  4.890 0.255 4.970 0.415 ;
        RECT  4.610 0.345 4.890 0.415 ;
        RECT  3.440 0.985 4.800 1.055 ;
        RECT  4.490 0.205 4.610 0.415 ;
        RECT  4.175 0.345 4.490 0.415 ;
        RECT  4.070 0.190 4.175 0.415 ;
        RECT  3.740 0.345 4.070 0.415 ;
        RECT  3.635 0.190 3.740 0.415 ;
        RECT  3.360 0.345 3.635 0.415 ;
        RECT  3.260 0.190 3.360 0.415 ;
        RECT  1.730 0.345 3.260 0.415 ;
        RECT  0.220 0.195 3.180 0.265 ;
        RECT  1.925 0.985 3.180 1.055 ;
        RECT  0.215 0.985 1.495 1.055 ;
    END
END OAI222D4BWP40

MACRO OAI22D0BWP40
    CLASS CORE ;
    FOREIGN OAI22D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.079600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.335 0.915 0.545 1.045 ;
        RECT  0.335 0.345 0.360 0.430 ;
        RECT  0.265 0.345 0.335 1.045 ;
        RECT  0.240 0.345 0.265 0.430 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.835 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.405 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.250 ;
        RECT  0.000 -0.115 0.640 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 1.145 0.980 1.375 ;
        RECT  0.855 0.945 0.925 1.375 ;
        RECT  0.130 1.145 0.855 1.375 ;
        RECT  0.055 0.945 0.130 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.840 0.195 0.940 0.415 ;
        RECT  0.570 0.345 0.840 0.415 ;
        RECT  0.500 0.205 0.570 0.415 ;
        RECT  0.035 0.205 0.500 0.275 ;
    END
END OAI22D0BWP40

MACRO OAI22D1BWP40
    CLASS CORE ;
    FOREIGN OAI22D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.134000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.335 0.915 0.545 1.045 ;
        RECT  0.335 0.345 0.360 0.430 ;
        RECT  0.265 0.345 0.335 1.045 ;
        RECT  0.240 0.345 0.265 0.430 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.765 ;
        RECT  0.735 0.495 0.875 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.835 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.195 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.405 0.495 0.455 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.250 ;
        RECT  0.000 -0.115 0.640 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 1.145 0.980 1.375 ;
        RECT  0.855 0.855 0.925 1.375 ;
        RECT  0.130 1.145 0.855 1.375 ;
        RECT  0.055 0.845 0.130 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.850 0.265 0.925 0.415 ;
        RECT  0.570 0.345 0.850 0.415 ;
        RECT  0.500 0.205 0.570 0.415 ;
        RECT  0.035 0.205 0.500 0.275 ;
    END
END OAI22D1BWP40

MACRO OAI22D2BWP40
    CLASS CORE ;
    FOREIGN OAI22D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.301200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.345 1.785 1.055 ;
        RECT  1.015 0.345 1.715 0.415 ;
        RECT  0.130 0.985 1.715 1.055 ;
        RECT  0.035 0.855 0.130 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.570 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.495 0.805 0.775 ;
        RECT  0.245 0.705 0.700 0.775 ;
        RECT  0.170 0.495 0.245 0.775 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.505 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.495 1.645 0.775 ;
        RECT  1.085 0.705 1.575 0.775 ;
        RECT  0.950 0.495 1.085 0.775 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.115 1.820 0.115 ;
        RECT  0.620 -0.115 0.740 0.275 ;
        RECT  0.340 -0.115 0.620 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.820 1.375 ;
        RECT  1.200 1.125 1.320 1.375 ;
        RECT  0.540 1.145 1.200 1.375 ;
        RECT  0.420 1.125 0.540 1.375 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.920 0.205 1.760 0.275 ;
        RECT  1.000 0.845 1.530 0.915 ;
        RECT  0.840 0.205 0.920 0.415 ;
        RECT  0.130 0.345 0.840 0.415 ;
        RECT  0.220 0.845 0.750 0.915 ;
        RECT  0.050 0.255 0.130 0.415 ;
    END
END OAI22D2BWP40

MACRO OAI22D3BWP40
    CLASS CORE ;
    FOREIGN OAI22D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.385000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.335 2.300 0.405 ;
        RECT  1.855 0.335 1.925 0.790 ;
        RECT  1.395 0.335 1.855 0.405 ;
        RECT  0.735 0.720 1.855 0.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.490 0.525 0.765 ;
        RECT  0.165 0.490 0.455 0.640 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.495 1.010 0.640 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.495 2.405 0.625 ;
        RECT  2.135 0.495 2.205 0.765 ;
        RECT  2.005 0.495 2.135 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.785 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.100 -0.115 2.520 0.115 ;
        RECT  0.980 -0.115 1.100 0.215 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.215 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.215 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.720 2.470 1.375 ;
        RECT  2.110 1.145 2.390 1.375 ;
        RECT  1.985 1.025 2.110 1.375 ;
        RECT  0.530 1.145 1.985 1.375 ;
        RECT  0.410 1.040 0.530 1.375 ;
        RECT  0.130 1.145 0.410 1.375 ;
        RECT  0.050 0.720 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.390 0.195 2.470 0.335 ;
        RECT  1.300 0.195 2.390 0.265 ;
        RECT  1.405 0.875 2.310 0.945 ;
        RECT  1.220 0.195 1.300 0.395 ;
        RECT  0.130 0.325 1.220 0.395 ;
        RECT  0.210 0.875 1.115 0.945 ;
        RECT  0.050 0.255 0.130 0.395 ;
    END
END OAI22D3BWP40

MACRO OAI22D4BWP40
    CLASS CORE ;
    FOREIGN OAI22D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.517000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 0.705 3.270 0.775 ;
        RECT  2.570 0.355 2.640 0.775 ;
        RECT  0.735 0.355 2.570 0.425 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.125 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.435 0.625 ;
        RECT  1.925 0.495 1.995 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.495 3.315 0.625 ;
        RECT  2.835 0.355 2.905 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.435 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.115 3.500 0.115 ;
        RECT  3.375 -0.115 3.445 0.420 ;
        RECT  3.060 -0.115 3.375 0.115 ;
        RECT  2.940 -0.115 3.060 0.140 ;
        RECT  2.660 -0.115 2.940 0.115 ;
        RECT  2.540 -0.115 2.660 0.140 ;
        RECT  2.240 -0.115 2.540 0.115 ;
        RECT  2.120 -0.115 2.240 0.140 ;
        RECT  1.850 -0.115 2.120 0.115 ;
        RECT  1.730 -0.115 1.850 0.140 ;
        RECT  0.000 -0.115 1.730 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.145 3.500 1.375 ;
        RECT  2.330 1.005 2.450 1.375 ;
        RECT  2.030 1.145 2.330 1.375 ;
        RECT  1.950 0.985 2.030 1.375 ;
        RECT  1.460 1.145 1.950 1.375 ;
        RECT  1.380 0.995 1.460 1.375 ;
        RECT  1.090 1.145 1.380 1.375 ;
        RECT  1.010 0.995 1.090 1.375 ;
        RECT  0.000 1.145 1.010 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.640 0.705 3.270 0.775 ;
        RECT  2.570 0.355 2.640 0.775 ;
        RECT  0.805 0.355 2.570 0.425 ;
        RECT  0.125 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  3.370 0.755 3.450 1.045 ;
        RECT  1.850 0.845 3.370 0.915 ;
        RECT  0.220 0.215 3.280 0.285 ;
        RECT  1.735 0.845 1.850 1.055 ;
        RECT  1.550 0.845 1.665 1.055 ;
        RECT  0.930 0.845 1.550 0.915 ;
        RECT  0.860 0.845 0.930 1.050 ;
        RECT  0.130 0.980 0.860 1.050 ;
        RECT  0.050 0.890 0.130 1.050 ;
    END
END OAI22D4BWP40

MACRO OAI22D6BWP40
    CLASS CORE ;
    FOREIGN OAI22D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.766000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.785 0.705 4.810 0.775 ;
        RECT  3.715 0.355 3.785 0.775 ;
        RECT  0.735 0.355 3.715 0.425 ;
        RECT  0.735 0.840 1.100 0.910 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.125 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.755 0.495 3.635 0.625 ;
        RECT  2.685 0.495 2.755 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 0.495 4.585 0.625 ;
        RECT  4.095 0.355 4.165 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.495 2.195 0.625 ;
        RECT  1.295 0.495 1.365 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.192000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.985 0.420 ;
        RECT  4.600 -0.115 4.915 0.115 ;
        RECT  4.480 -0.115 4.600 0.140 ;
        RECT  4.210 -0.115 4.480 0.115 ;
        RECT  4.090 -0.115 4.210 0.140 ;
        RECT  3.810 -0.115 4.090 0.115 ;
        RECT  3.690 -0.115 3.810 0.140 ;
        RECT  3.415 -0.115 3.690 0.115 ;
        RECT  3.285 -0.115 3.415 0.140 ;
        RECT  3.000 -0.115 3.285 0.115 ;
        RECT  2.880 -0.115 3.000 0.140 ;
        RECT  2.610 -0.115 2.880 0.115 ;
        RECT  2.490 -0.115 2.610 0.140 ;
        RECT  0.000 -0.115 2.490 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.145 5.040 1.375 ;
        RECT  3.490 1.005 3.610 1.375 ;
        RECT  3.210 1.145 3.490 1.375 ;
        RECT  3.090 1.005 3.210 1.375 ;
        RECT  2.790 1.145 3.090 1.375 ;
        RECT  2.710 0.985 2.790 1.375 ;
        RECT  2.220 1.145 2.710 1.375 ;
        RECT  2.140 0.995 2.220 1.375 ;
        RECT  1.840 1.145 2.140 1.375 ;
        RECT  1.760 0.995 1.840 1.375 ;
        RECT  1.455 1.145 1.760 1.375 ;
        RECT  1.380 0.985 1.455 1.375 ;
        RECT  0.000 1.145 1.380 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.705 4.810 0.775 ;
        RECT  3.715 0.355 3.785 0.775 ;
        RECT  0.805 0.355 3.715 0.425 ;
        RECT  0.805 0.840 1.100 0.910 ;
        RECT  0.125 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  4.910 0.755 4.990 1.050 ;
        RECT  4.585 0.845 4.910 0.915 ;
        RECT  4.700 0.215 4.805 0.445 ;
        RECT  0.220 0.215 4.700 0.285 ;
        RECT  4.500 0.845 4.585 1.075 ;
        RECT  4.195 0.845 4.500 0.915 ;
        RECT  4.110 0.845 4.195 1.075 ;
        RECT  3.790 0.845 4.110 0.915 ;
        RECT  3.710 0.845 3.790 1.075 ;
        RECT  3.390 0.845 3.710 0.915 ;
        RECT  3.310 0.845 3.390 1.075 ;
        RECT  2.990 0.845 3.310 0.915 ;
        RECT  2.915 0.845 2.990 1.075 ;
        RECT  2.610 0.845 2.915 0.915 ;
        RECT  2.495 0.845 2.610 1.055 ;
        RECT  2.310 0.845 2.425 1.055 ;
        RECT  1.265 0.845 2.310 0.915 ;
        RECT  1.195 0.845 1.265 1.050 ;
        RECT  0.130 0.980 1.195 1.050 ;
        RECT  0.050 0.890 0.130 1.050 ;
    END
END OAI22D6BWP40

MACRO OAI22D8BWP40
    CLASS CORE ;
    FOREIGN OAI22D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.580 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 1.006000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.925 0.705 6.350 0.775 ;
        RECT  4.855 0.355 4.925 0.775 ;
        RECT  0.735 0.355 4.855 0.425 ;
        RECT  0.735 0.840 1.480 0.910 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.125 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.249600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.465 0.495 4.765 0.625 ;
        RECT  3.395 0.495 3.465 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.254400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.035 0.495 6.395 0.625 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.780 0.495 2.955 0.625 ;
        RECT  1.710 0.495 1.780 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.256000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.525 -0.115 6.580 0.115 ;
        RECT  6.455 -0.115 6.525 0.400 ;
        RECT  6.140 -0.115 6.455 0.115 ;
        RECT  6.020 -0.115 6.140 0.210 ;
        RECT  5.750 -0.115 6.020 0.115 ;
        RECT  5.630 -0.115 5.750 0.210 ;
        RECT  5.325 -0.115 5.630 0.115 ;
        RECT  5.230 -0.115 5.325 0.260 ;
        RECT  4.950 -0.115 5.230 0.115 ;
        RECT  4.830 -0.115 4.950 0.140 ;
        RECT  4.570 -0.115 4.830 0.115 ;
        RECT  4.450 -0.115 4.570 0.140 ;
        RECT  4.170 -0.115 4.450 0.115 ;
        RECT  4.050 -0.115 4.170 0.140 ;
        RECT  3.760 -0.115 4.050 0.115 ;
        RECT  3.640 -0.115 3.760 0.140 ;
        RECT  3.370 -0.115 3.640 0.115 ;
        RECT  3.250 -0.115 3.370 0.140 ;
        RECT  0.000 -0.115 3.250 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.760 1.145 6.580 1.375 ;
        RECT  4.640 1.005 4.760 1.375 ;
        RECT  4.370 1.145 4.640 1.375 ;
        RECT  4.250 1.005 4.370 1.375 ;
        RECT  3.970 1.145 4.250 1.375 ;
        RECT  3.850 1.005 3.970 1.375 ;
        RECT  3.550 1.145 3.850 1.375 ;
        RECT  3.470 0.985 3.550 1.375 ;
        RECT  2.980 1.145 3.470 1.375 ;
        RECT  2.900 0.995 2.980 1.375 ;
        RECT  2.600 1.145 2.900 1.375 ;
        RECT  2.520 0.995 2.600 1.375 ;
        RECT  2.215 1.145 2.520 1.375 ;
        RECT  2.140 0.985 2.215 1.375 ;
        RECT  1.835 1.145 2.140 1.375 ;
        RECT  1.765 0.985 1.835 1.375 ;
        RECT  0.000 1.145 1.765 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.925 0.705 6.350 0.775 ;
        RECT  4.855 0.355 4.925 0.775 ;
        RECT  0.805 0.355 4.855 0.425 ;
        RECT  0.805 0.840 1.480 0.910 ;
        RECT  0.125 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  6.455 0.755 6.525 1.055 ;
        RECT  6.450 0.755 6.455 0.915 ;
        RECT  6.115 0.845 6.450 0.915 ;
        RECT  5.115 0.335 6.360 0.405 ;
        RECT  6.045 0.845 6.115 1.075 ;
        RECT  5.725 0.845 6.045 0.915 ;
        RECT  5.655 0.845 5.725 1.075 ;
        RECT  5.315 0.845 5.655 0.915 ;
        RECT  5.245 0.845 5.315 1.075 ;
        RECT  4.925 0.845 5.245 0.915 ;
        RECT  5.040 0.215 5.115 0.405 ;
        RECT  0.220 0.215 5.040 0.285 ;
        RECT  4.855 0.845 4.925 1.075 ;
        RECT  4.545 0.845 4.855 0.915 ;
        RECT  4.475 0.845 4.545 1.075 ;
        RECT  4.145 0.845 4.475 0.915 ;
        RECT  4.075 0.845 4.145 1.075 ;
        RECT  3.745 0.845 4.075 0.915 ;
        RECT  3.675 0.845 3.745 1.075 ;
        RECT  3.370 0.845 3.675 0.915 ;
        RECT  3.255 0.845 3.370 1.055 ;
        RECT  3.070 0.845 3.185 1.055 ;
        RECT  1.645 0.845 3.070 0.915 ;
        RECT  1.575 0.845 1.645 1.050 ;
        RECT  0.130 0.980 1.575 1.050 ;
        RECT  0.860 0.495 1.525 0.625 ;
        RECT  0.050 0.890 0.130 1.050 ;
    END
END OAI22D8BWP40

MACRO OAI31D0BWP40
    CLASS CORE ;
    FOREIGN OAI31D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.097250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.970 0.740 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.055 0.200 0.125 0.415 ;
        RECT  0.035 0.200 0.055 0.290 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.635 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 -0.115 0.980 0.115 ;
        RECT  0.835 -0.115 0.935 0.285 ;
        RECT  0.000 -0.115 0.835 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.840 0.940 0.930 1.375 ;
        RECT  0.135 1.145 0.840 1.375 ;
        RECT  0.050 0.940 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.230 0.205 0.740 0.275 ;
    END
END OAI31D0BWP40

MACRO OAI31D1BWP40
    CLASS CORE ;
    FOREIGN OAI31D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.170500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.970 0.740 1.045 ;
        RECT  0.455 0.345 0.525 1.045 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.055 0.215 0.125 0.415 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.495 0.945 0.635 ;
        RECT  0.735 0.495 0.805 0.765 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.810 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 -0.115 0.980 0.115 ;
        RECT  0.835 -0.115 0.935 0.425 ;
        RECT  0.000 -0.115 0.835 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.145 0.980 1.375 ;
        RECT  0.830 0.860 0.930 1.375 ;
        RECT  0.150 1.145 0.830 1.375 ;
        RECT  0.050 0.850 0.150 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 0.205 0.740 0.415 ;
        RECT  0.230 0.205 0.620 0.275 ;
    END
END OAI31D1BWP40

MACRO OAI31D2BWP40
    CLASS CORE ;
    FOREIGN OAI31D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.287900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.365 0.775 1.505 0.905 ;
        RECT  1.285 0.340 1.365 1.055 ;
        RECT  0.220 0.340 1.285 0.410 ;
        RECT  0.595 0.985 1.285 1.055 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.059200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.695 0.495 1.785 0.765 ;
        RECT  1.505 0.495 1.695 0.630 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.059200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.059200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.000 0.770 ;
        RECT  0.435 0.700 0.875 0.770 ;
        RECT  0.345 0.495 0.435 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.059200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.510 1.195 0.915 ;
        RECT  0.255 0.845 1.115 0.915 ;
        RECT  0.170 0.495 0.255 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 -0.115 1.820 0.115 ;
        RECT  1.425 -0.115 1.545 0.130 ;
        RECT  0.000 -0.115 1.425 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.145 1.820 1.375 ;
        RECT  1.670 0.845 1.750 1.375 ;
        RECT  1.310 1.145 1.670 1.375 ;
        RECT  1.190 1.130 1.310 1.375 ;
        RECT  0.125 1.145 1.190 1.375 ;
        RECT  0.050 0.980 0.125 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.675 0.200 1.745 0.370 ;
        RECT  0.130 0.200 1.675 0.270 ;
        RECT  0.050 0.200 0.130 0.380 ;
    END
END OAI31D2BWP40

MACRO OAI31D4BWP40
    CLASS CORE ;
    FOREIGN OAI31D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.605200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.845 3.270 1.055 ;
        RECT  2.850 0.845 3.150 0.915 ;
        RECT  2.730 0.845 2.850 1.055 ;
        RECT  2.685 0.845 2.730 0.915 ;
        RECT  2.575 0.355 2.685 0.915 ;
        RECT  0.735 0.355 2.575 0.425 ;
        RECT  0.525 0.355 0.735 0.910 ;
        RECT  0.125 0.355 0.525 0.425 ;
        RECT  0.220 0.840 0.525 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.185 0.765 ;
        RECT  2.805 0.495 3.115 0.625 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.445 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.435 0.625 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.121600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.495 2.485 0.765 ;
        RECT  1.945 0.495 2.415 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.270 -0.115 3.500 0.115 ;
        RECT  3.150 -0.115 3.270 0.230 ;
        RECT  2.850 -0.115 3.150 0.115 ;
        RECT  2.730 -0.115 2.850 0.145 ;
        RECT  0.000 -0.115 2.730 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.710 3.450 1.375 ;
        RECT  3.040 1.145 3.370 1.375 ;
        RECT  2.960 0.985 3.040 1.375 ;
        RECT  2.630 1.145 2.960 1.375 ;
        RECT  2.550 0.985 2.630 1.375 ;
        RECT  2.220 1.145 2.550 1.375 ;
        RECT  2.140 0.985 2.220 1.375 ;
        RECT  1.825 1.145 2.140 1.375 ;
        RECT  1.755 0.990 1.825 1.375 ;
        RECT  0.000 1.145 1.755 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.845 3.270 1.055 ;
        RECT  2.850 0.845 3.150 0.915 ;
        RECT  2.730 0.845 2.850 1.055 ;
        RECT  2.685 0.845 2.730 0.915 ;
        RECT  2.575 0.355 2.685 0.915 ;
        RECT  0.805 0.355 2.575 0.425 ;
        RECT  0.125 0.355 0.455 0.425 ;
        RECT  0.220 0.840 0.455 0.910 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  3.370 0.230 3.450 0.400 ;
        RECT  3.040 0.330 3.370 0.400 ;
        RECT  2.965 0.215 3.040 0.400 ;
        RECT  0.220 0.215 2.965 0.285 ;
        RECT  2.325 0.845 2.445 1.055 ;
        RECT  2.040 0.845 2.325 0.915 ;
        RECT  1.920 0.845 2.040 1.055 ;
        RECT  0.980 0.845 1.920 0.915 ;
        RECT  0.130 0.985 1.670 1.055 ;
        RECT  0.050 0.890 0.130 1.055 ;
    END
END OAI31D4BWP40

MACRO OAI32D0BWP40
    CLASS CORE ;
    FOREIGN OAI32D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.109750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.890 0.805 1.045 ;
        RECT  0.105 0.890 0.700 0.960 ;
        RECT  0.140 0.345 0.600 0.415 ;
        RECT  0.105 0.205 0.140 0.415 ;
        RECT  0.035 0.205 0.105 0.960 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.810 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.155 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.495 0.805 0.630 ;
        RECT  0.595 0.495 0.665 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.115 1.260 0.115 ;
        RECT  0.915 -0.115 1.015 0.275 ;
        RECT  0.000 -0.115 0.915 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.950 1.210 1.375 ;
        RECT  0.165 1.145 1.130 1.375 ;
        RECT  0.045 1.030 0.165 1.375 ;
        RECT  0.000 1.145 0.045 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.185 1.205 0.415 ;
        RECT  0.820 0.345 1.135 0.415 ;
        RECT  0.750 0.205 0.820 0.415 ;
        RECT  0.250 0.205 0.750 0.275 ;
    END
END OAI32D0BWP40

MACRO OAI32D1BWP40
    CLASS CORE ;
    FOREIGN OAI32D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.194500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.890 0.805 0.960 ;
        RECT  0.130 0.345 0.600 0.415 ;
        RECT  0.105 0.215 0.130 0.415 ;
        RECT  0.035 0.215 0.105 0.960 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 0.945 0.810 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.225 0.765 ;
        RECT  1.015 0.495 1.155 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.805 0.765 ;
        RECT  0.595 0.495 0.735 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.525 0.765 ;
        RECT  0.315 0.495 0.455 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.245 0.810 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.115 1.260 0.115 ;
        RECT  0.915 -0.115 1.015 0.275 ;
        RECT  0.000 -0.115 0.915 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.145 1.260 1.375 ;
        RECT  1.130 0.860 1.210 1.375 ;
        RECT  0.165 1.145 1.130 1.375 ;
        RECT  0.045 1.030 0.165 1.375 ;
        RECT  0.000 1.145 0.045 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.135 0.255 1.205 0.415 ;
        RECT  0.775 0.345 1.135 0.415 ;
        RECT  0.705 0.205 0.775 0.415 ;
        RECT  0.250 0.205 0.705 0.275 ;
    END
END OAI32D1BWP40

MACRO OAI32D2BWP40
    CLASS CORE ;
    FOREIGN OAI32D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.284100 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.985 1.785 1.055 ;
        RECT  1.330 0.915 1.575 1.055 ;
        RECT  1.260 0.340 1.330 1.055 ;
        RECT  0.220 0.340 1.260 0.410 ;
        RECT  0.595 0.985 1.260 1.055 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.495 1.785 0.770 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.355 2.065 0.640 ;
        RECT  1.575 0.355 1.945 0.425 ;
        RECT  1.505 0.355 1.575 0.640 ;
        RECT  1.400 0.495 1.505 0.640 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.015 0.765 ;
        RECT  0.435 0.695 0.875 0.765 ;
        RECT  0.325 0.495 0.435 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 0.495 1.190 0.915 ;
        RECT  0.255 0.845 1.110 0.915 ;
        RECT  0.170 0.495 0.255 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.970 -0.115 2.240 0.115 ;
        RECT  1.850 -0.115 1.970 0.130 ;
        RECT  1.570 -0.115 1.850 0.115 ;
        RECT  1.450 -0.115 1.570 0.130 ;
        RECT  0.000 -0.115 1.450 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.145 2.240 1.375 ;
        RECT  2.110 0.770 2.190 1.375 ;
        RECT  1.360 1.145 2.110 1.375 ;
        RECT  1.240 1.125 1.360 1.375 ;
        RECT  0.130 1.145 1.240 1.375 ;
        RECT  0.050 0.980 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.130 0.200 2.180 0.270 ;
        RECT  0.050 0.200 0.130 0.385 ;
    END
END OAI32D2BWP40

MACRO OAI32D4BWP40
    CLASS CORE ;
    FOREIGN OAI32D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.621000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.995 3.370 1.065 ;
        RECT  2.555 0.845 2.560 1.065 ;
        RECT  2.490 0.455 2.555 1.065 ;
        RECT  2.420 0.455 2.490 0.915 ;
        RECT  2.345 0.345 2.420 0.915 ;
        RECT  0.220 0.345 2.345 0.415 ;
        RECT  1.735 0.845 2.345 0.915 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.495 3.185 0.765 ;
        RECT  2.780 0.495 3.115 0.630 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.495 4.165 0.630 ;
        RECT  3.675 0.495 3.745 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.135 0.495 2.205 0.765 ;
        RECT  1.865 0.495 2.135 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.495 1.505 0.765 ;
        RECT  0.940 0.495 1.435 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.805 0.640 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.125 -0.115 4.340 0.115 ;
        RECT  3.995 -0.115 4.125 0.230 ;
        RECT  3.740 -0.115 3.995 0.115 ;
        RECT  3.615 -0.115 3.740 0.235 ;
        RECT  3.180 -0.115 3.615 0.115 ;
        RECT  3.060 -0.115 3.180 0.235 ;
        RECT  2.800 -0.115 3.060 0.115 ;
        RECT  2.680 -0.115 2.800 0.235 ;
        RECT  0.000 -0.115 2.680 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.290 1.145 4.340 1.375 ;
        RECT  4.210 0.720 4.290 1.375 ;
        RECT  3.935 1.145 4.210 1.375 ;
        RECT  3.810 1.005 3.935 1.375 ;
        RECT  3.530 1.145 3.810 1.375 ;
        RECT  3.450 0.995 3.530 1.375 ;
        RECT  0.725 1.145 3.450 1.375 ;
        RECT  0.595 1.030 0.725 1.375 ;
        RECT  0.345 1.145 0.595 1.375 ;
        RECT  0.215 1.030 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.625 0.995 3.370 1.065 ;
        RECT  0.220 0.345 2.275 0.415 ;
        RECT  1.735 0.845 2.275 0.915 ;
        RECT  4.210 0.205 4.290 0.375 ;
        RECT  2.590 0.305 4.210 0.375 ;
        RECT  2.665 0.845 4.125 0.915 ;
        RECT  2.510 0.195 2.590 0.375 ;
        RECT  0.130 0.195 2.510 0.265 ;
        RECT  0.975 0.995 2.420 1.065 ;
        RECT  0.035 0.845 1.665 0.915 ;
        RECT  0.050 0.195 0.130 0.455 ;
    END
END OAI32D4BWP40

MACRO OAI33D0BWP40
    CLASS CORE ;
    FOREIGN OAI33D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.100325 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.935 0.760 1.025 ;
        RECT  0.455 0.345 0.525 1.025 ;
        RECT  0.150 0.345 0.455 0.415 ;
        RECT  0.035 0.215 0.150 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.810 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.820 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.495 1.365 0.765 ;
        RECT  1.155 0.495 1.290 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.820 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.110 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.275 ;
        RECT  0.960 -0.115 1.260 0.115 ;
        RECT  0.840 -0.115 0.960 0.270 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.960 1.360 1.375 ;
        RECT  0.140 1.145 1.260 1.375 ;
        RECT  0.040 0.930 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.200 1.170 0.410 ;
        RECT  0.735 0.340 1.050 0.410 ;
        RECT  0.665 0.195 0.735 0.410 ;
        RECT  0.220 0.195 0.665 0.265 ;
    END
END OAI33D0BWP40

MACRO OAI33D1BWP40
    CLASS CORE ;
    FOREIGN OAI33D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.172750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.935 0.760 1.025 ;
        RECT  0.455 0.345 0.525 1.025 ;
        RECT  0.125 0.345 0.455 0.415 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.495 0.945 0.625 ;
        RECT  0.735 0.495 0.810 0.765 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.820 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.495 1.365 0.625 ;
        RECT  1.155 0.495 1.230 0.765 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.820 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.905 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.110 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 -0.115 1.400 0.115 ;
        RECT  1.260 -0.115 1.360 0.275 ;
        RECT  0.960 -0.115 1.260 0.115 ;
        RECT  0.840 -0.115 0.960 0.270 ;
        RECT  0.000 -0.115 0.840 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.145 1.400 1.375 ;
        RECT  1.260 0.870 1.360 1.375 ;
        RECT  0.140 1.145 1.260 1.375 ;
        RECT  0.040 0.870 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 0.200 1.170 0.410 ;
        RECT  0.735 0.340 1.050 0.410 ;
        RECT  0.665 0.195 0.735 0.410 ;
        RECT  0.220 0.195 0.665 0.265 ;
    END
END OAI33D1BWP40

MACRO OAI33D2BWP40
    CLASS CORE ;
    FOREIGN OAI33D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.300500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.335 2.485 1.060 ;
        RECT  1.365 0.335 2.415 0.405 ;
        RECT  0.595 0.990 2.415 1.060 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.495 0.845 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 0.485 1.015 0.765 ;
        RECT  0.405 0.695 0.915 0.765 ;
        RECT  0.315 0.485 0.405 0.765 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.515 1.225 0.645 ;
        RECT  1.085 0.515 1.155 0.920 ;
        RECT  0.245 0.850 1.085 0.920 ;
        RECT  0.130 0.495 0.245 0.920 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 0.495 1.925 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 0.495 2.125 0.765 ;
        RECT  1.585 0.695 1.995 0.765 ;
        RECT  1.435 0.485 1.585 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 0.490 2.345 0.920 ;
        RECT  1.365 0.850 2.245 0.920 ;
        RECT  1.295 0.515 1.365 0.920 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.100 -0.115 2.520 0.115 ;
        RECT  0.980 -0.115 1.100 0.275 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.275 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.145 2.520 1.375 ;
        RECT  2.315 1.130 2.450 1.375 ;
        RECT  1.300 1.145 2.315 1.375 ;
        RECT  1.180 1.130 1.300 1.375 ;
        RECT  0.130 1.145 1.180 1.375 ;
        RECT  0.050 1.060 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.265 0.195 2.475 0.265 ;
        RECT  1.195 0.195 1.265 0.415 ;
        RECT  0.885 0.345 1.195 0.415 ;
        RECT  0.815 0.185 0.885 0.415 ;
        RECT  0.505 0.345 0.815 0.415 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.125 0.345 0.435 0.415 ;
        RECT  0.055 0.255 0.125 0.415 ;
    END
END OAI33D2BWP40

MACRO OAI33D3BWP40
    CLASS CORE ;
    FOREIGN OAI33D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.452750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.770 2.250 0.850 ;
        RECT  1.735 0.495 1.850 0.850 ;
        RECT  1.665 0.345 1.735 0.850 ;
        RECT  0.125 0.345 1.665 0.415 ;
        RECT  1.350 0.770 1.665 0.850 ;
        RECT  0.035 0.215 0.125 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.495 2.220 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.495 2.830 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 0.495 3.365 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.520 0.650 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.495 1.085 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.425 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.565 -0.115 3.640 0.115 ;
        RECT  3.465 -0.115 3.565 0.405 ;
        RECT  3.200 -0.115 3.465 0.115 ;
        RECT  3.070 -0.115 3.200 0.275 ;
        RECT  2.820 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.820 0.275 ;
        RECT  2.440 -0.115 2.690 0.115 ;
        RECT  2.305 -0.115 2.440 0.275 ;
        RECT  2.025 -0.115 2.305 0.115 ;
        RECT  1.955 -0.115 2.025 0.275 ;
        RECT  0.000 -0.115 1.955 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.565 1.145 3.640 1.375 ;
        RECT  3.465 0.705 3.565 1.375 ;
        RECT  3.195 1.145 3.465 1.375 ;
        RECT  3.075 0.905 3.195 1.375 ;
        RECT  0.530 1.145 3.075 1.375 ;
        RECT  0.410 0.905 0.530 1.375 ;
        RECT  0.140 1.145 0.410 1.375 ;
        RECT  0.040 0.725 0.140 1.375 ;
        RECT  0.000 1.145 0.040 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.905 0.770 2.250 0.850 ;
        RECT  0.125 0.345 1.660 0.415 ;
        RECT  1.350 0.770 1.660 0.850 ;
        RECT  0.035 0.215 0.125 0.415 ;
        RECT  3.290 0.760 3.390 1.025 ;
        RECT  3.290 0.195 3.380 0.425 ;
        RECT  2.980 0.355 3.290 0.425 ;
        RECT  2.985 0.760 3.290 0.830 ;
        RECT  2.910 0.760 2.985 1.020 ;
        RECT  2.910 0.195 2.980 0.425 ;
        RECT  2.600 0.355 2.910 0.425 ;
        RECT  2.505 0.760 2.910 0.830 ;
        RECT  1.930 0.955 2.820 1.025 ;
        RECT  2.530 0.195 2.600 0.425 ;
        RECT  2.215 0.355 2.530 0.425 ;
        RECT  2.145 0.195 2.215 0.425 ;
        RECT  1.885 0.355 2.145 0.425 ;
        RECT  1.815 0.195 1.885 0.425 ;
        RECT  0.215 0.195 1.815 0.265 ;
        RECT  0.790 0.955 1.675 1.025 ;
        RECT  0.215 0.760 1.100 0.835 ;
    END
END OAI33D3BWP40

MACRO OAI33D4BWP40
    CLASS CORE ;
    FOREIGN OAI33D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.623250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.770 3.370 0.850 ;
        RECT  2.490 0.495 2.695 0.850 ;
        RECT  2.485 0.345 2.490 0.850 ;
        RECT  2.420 0.345 2.485 0.565 ;
        RECT  1.740 0.770 2.485 0.850 ;
        RECT  0.210 0.345 2.420 0.415 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 0.495 3.200 0.625 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.780 0.495 4.140 0.625 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.370 0.495 4.675 0.625 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.495 2.275 0.650 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.495 1.245 0.650 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 0.495 0.615 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.890 -0.115 5.180 0.115 ;
        RECT  4.760 -0.115 4.890 0.275 ;
        RECT  4.510 -0.115 4.760 0.115 ;
        RECT  4.380 -0.115 4.510 0.275 ;
        RECT  4.130 -0.115 4.380 0.115 ;
        RECT  4.000 -0.115 4.130 0.275 ;
        RECT  3.750 -0.115 4.000 0.115 ;
        RECT  3.620 -0.115 3.750 0.275 ;
        RECT  3.195 -0.115 3.620 0.115 ;
        RECT  3.060 -0.115 3.195 0.275 ;
        RECT  2.780 -0.115 3.060 0.115 ;
        RECT  2.710 -0.115 2.780 0.275 ;
        RECT  0.000 -0.115 2.710 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.145 5.180 1.375 ;
        RECT  4.760 0.905 4.890 1.375 ;
        RECT  4.510 1.145 4.760 1.375 ;
        RECT  4.380 0.905 4.510 1.375 ;
        RECT  0.725 1.145 4.380 1.375 ;
        RECT  0.595 0.905 0.725 1.375 ;
        RECT  0.345 1.145 0.595 1.375 ;
        RECT  0.215 0.905 0.345 1.375 ;
        RECT  0.000 1.145 0.215 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.765 0.770 3.370 0.850 ;
        RECT  0.210 0.345 2.415 0.415 ;
        RECT  1.740 0.770 2.415 0.850 ;
        RECT  5.030 0.195 5.120 0.425 ;
        RECT  5.030 0.755 5.100 1.055 ;
        RECT  4.670 0.355 5.030 0.425 ;
        RECT  4.670 0.755 5.030 0.825 ;
        RECT  4.600 0.195 4.670 0.425 ;
        RECT  4.600 0.755 4.670 1.015 ;
        RECT  4.290 0.355 4.600 0.425 ;
        RECT  4.290 0.755 4.600 0.825 ;
        RECT  4.220 0.195 4.290 0.425 ;
        RECT  4.220 0.755 4.290 1.015 ;
        RECT  3.910 0.355 4.220 0.425 ;
        RECT  3.440 0.755 4.220 0.825 ;
        RECT  2.685 0.955 4.130 1.025 ;
        RECT  3.840 0.195 3.910 0.425 ;
        RECT  3.530 0.355 3.840 0.425 ;
        RECT  3.460 0.195 3.530 0.425 ;
        RECT  3.350 0.355 3.460 0.425 ;
        RECT  3.280 0.195 3.350 0.425 ;
        RECT  2.970 0.355 3.280 0.425 ;
        RECT  2.900 0.195 2.970 0.425 ;
        RECT  2.640 0.355 2.900 0.425 ;
        RECT  2.570 0.195 2.640 0.425 ;
        RECT  0.035 0.195 2.570 0.265 ;
        RECT  0.980 0.955 2.430 1.025 ;
        RECT  0.035 0.755 1.670 0.830 ;
    END
END OAI33D4BWP40

MACRO OR2D0BWP40
    CLASS CORE ;
    FOREIGN OR2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.075 ;
        RECT  0.715 0.185 0.735 0.305 ;
        RECT  0.695 0.980 0.735 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 -0.115 0.840 0.115 ;
        RECT  0.470 -0.115 0.590 0.275 ;
        RECT  0.140 -0.115 0.470 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.145 0.840 1.375 ;
        RECT  0.470 0.985 0.590 1.375 ;
        RECT  0.000 1.145 0.470 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.915 ;
        RECT  0.350 0.355 0.595 0.425 ;
        RECT  0.130 0.845 0.595 0.915 ;
        RECT  0.270 0.185 0.350 0.425 ;
        RECT  0.050 0.845 0.130 1.060 ;
    END
END OR2D0BWP40

MACRO OR2D12BWP40
    CLASS CORE ;
    FOREIGN OR2D12BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.720000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.700 3.820 1.025 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.415 0.345 3.745 0.465 ;
        RECT  3.415 0.700 3.740 0.820 ;
        RECT  3.345 0.185 3.415 0.465 ;
        RECT  3.340 0.700 3.415 1.045 ;
        RECT  3.045 0.345 3.345 0.465 ;
        RECT  3.045 0.700 3.340 0.820 ;
        RECT  2.975 0.185 3.045 0.465 ;
        RECT  2.975 0.700 3.045 1.045 ;
        RECT  2.945 0.185 2.975 1.045 ;
        RECT  2.940 0.345 2.945 1.045 ;
        RECT  2.765 0.345 2.940 0.820 ;
        RECT  2.635 0.345 2.765 0.465 ;
        RECT  2.640 0.700 2.765 0.820 ;
        RECT  2.560 0.700 2.640 1.025 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.345 2.565 0.465 ;
        RECT  2.260 0.700 2.560 0.820 ;
        RECT  2.180 0.700 2.260 1.025 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.880 0.345 2.185 0.465 ;
        RECT  1.880 0.700 2.180 0.820 ;
        RECT  1.805 0.185 1.880 0.465 ;
        RECT  1.800 0.700 1.880 1.025 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.495 1.555 0.625 ;
        RECT  1.110 0.355 1.190 0.625 ;
        RECT  0.275 0.355 1.110 0.425 ;
        RECT  0.205 0.355 0.275 0.625 ;
        RECT  0.110 0.495 0.205 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.940 0.615 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 -0.115 4.060 0.115 ;
        RECT  3.930 -0.115 4.010 0.465 ;
        RECT  3.640 -0.115 3.930 0.115 ;
        RECT  3.520 -0.115 3.640 0.265 ;
        RECT  3.240 -0.115 3.520 0.115 ;
        RECT  3.120 -0.115 3.240 0.265 ;
        RECT  2.850 -0.115 3.120 0.115 ;
        RECT  2.730 -0.115 2.850 0.265 ;
        RECT  2.450 -0.115 2.730 0.115 ;
        RECT  2.370 -0.115 2.450 0.275 ;
        RECT  2.070 -0.115 2.370 0.115 ;
        RECT  1.990 -0.115 2.070 0.275 ;
        RECT  1.690 -0.115 1.990 0.115 ;
        RECT  1.610 -0.115 1.690 0.275 ;
        RECT  1.310 -0.115 1.610 0.115 ;
        RECT  1.190 -0.115 1.310 0.125 ;
        RECT  0.910 -0.115 1.190 0.115 ;
        RECT  0.790 -0.115 0.910 0.145 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.145 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.425 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.145 4.060 1.375 ;
        RECT  3.930 0.705 4.010 1.375 ;
        RECT  3.640 1.145 3.930 1.375 ;
        RECT  3.520 0.890 3.640 1.375 ;
        RECT  3.240 1.145 3.520 1.375 ;
        RECT  3.120 0.890 3.240 1.375 ;
        RECT  2.850 1.145 3.120 1.375 ;
        RECT  2.730 0.890 2.850 1.375 ;
        RECT  2.470 1.145 2.730 1.375 ;
        RECT  2.350 0.890 2.470 1.375 ;
        RECT  2.090 1.145 2.350 1.375 ;
        RECT  1.970 0.890 2.090 1.375 ;
        RECT  1.710 1.145 1.970 1.375 ;
        RECT  1.590 0.995 1.710 1.375 ;
        RECT  1.305 1.145 1.590 1.375 ;
        RECT  1.185 0.995 1.305 1.375 ;
        RECT  0.125 1.145 1.185 1.375 ;
        RECT  0.055 0.720 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.740 0.700 3.820 1.025 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.415 0.345 3.745 0.465 ;
        RECT  3.415 0.700 3.740 0.820 ;
        RECT  3.345 0.185 3.415 0.465 ;
        RECT  3.340 0.700 3.415 1.045 ;
        RECT  3.045 0.345 3.345 0.465 ;
        RECT  3.045 0.700 3.340 0.820 ;
        RECT  2.635 0.345 2.695 0.465 ;
        RECT  2.640 0.700 2.695 0.820 ;
        RECT  2.560 0.700 2.640 1.025 ;
        RECT  2.565 0.185 2.635 0.465 ;
        RECT  2.255 0.345 2.565 0.465 ;
        RECT  2.260 0.700 2.560 0.820 ;
        RECT  2.180 0.700 2.260 1.025 ;
        RECT  2.185 0.185 2.255 0.465 ;
        RECT  1.880 0.345 2.185 0.465 ;
        RECT  1.880 0.700 2.180 0.820 ;
        RECT  1.805 0.185 1.880 0.465 ;
        RECT  1.800 0.700 1.880 1.025 ;
        RECT  1.705 0.545 2.505 0.615 ;
        RECT  1.635 0.355 1.705 0.915 ;
        RECT  1.520 0.355 1.635 0.425 ;
        RECT  0.895 0.845 1.635 0.915 ;
        RECT  1.450 0.215 1.520 0.425 ;
        RECT  0.335 0.695 1.520 0.765 ;
        RECT  0.220 0.215 1.450 0.285 ;
        RECT  0.800 0.845 0.895 1.075 ;
        RECT  0.515 0.845 0.800 0.915 ;
        RECT  0.410 0.845 0.515 1.075 ;
        RECT  0.225 0.695 0.335 1.075 ;
    END
END OR2D12BWP40

MACRO OR2D16BWP40
    CLASS CORE ;
    FOREIGN OR2D16BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.960000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.275 0.185 5.370 0.465 ;
        RECT  5.280 0.700 5.360 1.025 ;
        RECT  4.980 0.700 5.280 0.820 ;
        RECT  4.985 0.345 5.275 0.465 ;
        RECT  4.900 0.185 4.985 0.465 ;
        RECT  4.900 0.700 4.980 1.025 ;
        RECT  4.600 0.345 4.900 0.465 ;
        RECT  4.600 0.700 4.900 0.820 ;
        RECT  4.525 0.185 4.600 0.465 ;
        RECT  4.520 0.700 4.600 1.025 ;
        RECT  4.215 0.345 4.525 0.465 ;
        RECT  4.215 0.700 4.520 0.820 ;
        RECT  4.145 0.185 4.215 0.465 ;
        RECT  4.140 0.700 4.215 1.045 ;
        RECT  4.095 0.345 4.145 0.465 ;
        RECT  4.095 0.700 4.140 0.820 ;
        RECT  3.885 0.345 4.095 0.820 ;
        RECT  3.815 0.345 3.885 0.465 ;
        RECT  3.815 0.700 3.885 0.820 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.740 0.700 3.815 1.025 ;
        RECT  3.435 0.345 3.745 0.465 ;
        RECT  3.440 0.700 3.740 0.820 ;
        RECT  3.360 0.700 3.440 1.025 ;
        RECT  3.365 0.185 3.435 0.465 ;
        RECT  3.055 0.345 3.365 0.465 ;
        RECT  3.060 0.700 3.360 0.820 ;
        RECT  2.980 0.700 3.060 1.025 ;
        RECT  2.985 0.185 3.055 0.465 ;
        RECT  2.680 0.345 2.985 0.465 ;
        RECT  2.680 0.700 2.980 0.820 ;
        RECT  2.605 0.185 2.680 0.465 ;
        RECT  2.600 0.700 2.680 1.025 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.495 2.355 0.625 ;
        RECT  1.435 0.355 1.530 0.625 ;
        RECT  0.245 0.355 1.435 0.425 ;
        RECT  0.135 0.355 0.245 0.645 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.187200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 1.325 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 -0.115 5.600 0.115 ;
        RECT  5.470 -0.115 5.550 0.465 ;
        RECT  5.190 -0.115 5.470 0.115 ;
        RECT  5.070 -0.115 5.190 0.265 ;
        RECT  4.810 -0.115 5.070 0.115 ;
        RECT  4.690 -0.115 4.810 0.265 ;
        RECT  4.430 -0.115 4.690 0.115 ;
        RECT  4.310 -0.115 4.430 0.265 ;
        RECT  4.040 -0.115 4.310 0.115 ;
        RECT  3.920 -0.115 4.040 0.265 ;
        RECT  3.650 -0.115 3.920 0.115 ;
        RECT  3.530 -0.115 3.650 0.265 ;
        RECT  3.250 -0.115 3.530 0.115 ;
        RECT  3.170 -0.115 3.250 0.275 ;
        RECT  2.870 -0.115 3.170 0.115 ;
        RECT  2.790 -0.115 2.870 0.275 ;
        RECT  2.490 -0.115 2.790 0.115 ;
        RECT  2.410 -0.115 2.490 0.275 ;
        RECT  2.090 -0.115 2.410 0.115 ;
        RECT  2.010 -0.115 2.090 0.265 ;
        RECT  1.690 -0.115 2.010 0.115 ;
        RECT  1.570 -0.115 1.690 0.125 ;
        RECT  1.290 -0.115 1.570 0.115 ;
        RECT  1.170 -0.115 1.290 0.145 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.145 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.145 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.280 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 1.145 5.600 1.375 ;
        RECT  5.470 0.720 5.550 1.375 ;
        RECT  5.190 1.145 5.470 1.375 ;
        RECT  5.070 0.890 5.190 1.375 ;
        RECT  4.810 1.145 5.070 1.375 ;
        RECT  4.690 0.890 4.810 1.375 ;
        RECT  4.430 1.145 4.690 1.375 ;
        RECT  4.310 0.890 4.430 1.375 ;
        RECT  4.040 1.145 4.310 1.375 ;
        RECT  3.920 0.890 4.040 1.375 ;
        RECT  3.650 1.145 3.920 1.375 ;
        RECT  3.530 0.890 3.650 1.375 ;
        RECT  3.270 1.145 3.530 1.375 ;
        RECT  3.150 0.890 3.270 1.375 ;
        RECT  2.890 1.145 3.150 1.375 ;
        RECT  2.770 0.890 2.890 1.375 ;
        RECT  2.490 1.145 2.770 1.375 ;
        RECT  2.410 0.880 2.490 1.375 ;
        RECT  2.090 1.145 2.410 1.375 ;
        RECT  2.010 0.985 2.090 1.375 ;
        RECT  1.670 1.145 2.010 1.375 ;
        RECT  1.580 0.985 1.670 1.375 ;
        RECT  0.125 1.145 1.580 1.375 ;
        RECT  0.055 0.725 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.275 0.185 5.370 0.465 ;
        RECT  5.280 0.700 5.360 1.025 ;
        RECT  4.980 0.700 5.280 0.820 ;
        RECT  4.985 0.345 5.275 0.465 ;
        RECT  4.900 0.185 4.985 0.465 ;
        RECT  4.900 0.700 4.980 1.025 ;
        RECT  4.600 0.345 4.900 0.465 ;
        RECT  4.600 0.700 4.900 0.820 ;
        RECT  4.525 0.185 4.600 0.465 ;
        RECT  4.520 0.700 4.600 1.025 ;
        RECT  4.215 0.345 4.525 0.465 ;
        RECT  4.215 0.700 4.520 0.820 ;
        RECT  4.165 0.185 4.215 0.465 ;
        RECT  4.165 0.700 4.215 1.045 ;
        RECT  3.745 0.185 3.815 0.465 ;
        RECT  3.740 0.700 3.815 1.025 ;
        RECT  3.435 0.345 3.745 0.465 ;
        RECT  3.440 0.700 3.740 0.820 ;
        RECT  3.360 0.700 3.440 1.025 ;
        RECT  3.365 0.185 3.435 0.465 ;
        RECT  3.055 0.345 3.365 0.465 ;
        RECT  3.060 0.700 3.360 0.820 ;
        RECT  2.980 0.700 3.060 1.025 ;
        RECT  2.985 0.185 3.055 0.465 ;
        RECT  2.680 0.345 2.985 0.465 ;
        RECT  2.680 0.700 2.980 0.820 ;
        RECT  2.605 0.185 2.680 0.465 ;
        RECT  2.600 0.700 2.680 1.025 ;
        RECT  2.505 0.545 3.735 0.615 ;
        RECT  2.435 0.355 2.505 0.765 ;
        RECT  2.315 0.355 2.435 0.425 ;
        RECT  0.410 0.695 2.435 0.765 ;
        RECT  2.205 0.195 2.315 0.425 ;
        RECT  2.220 0.845 2.315 1.075 ;
        RECT  1.875 0.845 2.220 0.915 ;
        RECT  1.895 0.355 2.205 0.425 ;
        RECT  1.785 0.215 1.895 0.425 ;
        RECT  1.800 0.845 1.875 1.075 ;
        RECT  1.455 0.845 1.800 0.915 ;
        RECT  0.220 0.215 1.785 0.285 ;
        RECT  1.380 0.845 1.455 1.075 ;
        RECT  1.075 0.845 1.380 0.915 ;
        RECT  1.000 0.845 1.075 1.075 ;
        RECT  0.695 0.845 1.000 0.915 ;
        RECT  0.620 0.845 0.695 1.075 ;
        RECT  0.330 0.845 0.620 0.915 ;
        RECT  0.225 0.845 0.330 1.075 ;
    END
END OR2D16BWP40

MACRO OR2D1BWP40
    CLASS CORE ;
    FOREIGN OR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.185 0.805 1.075 ;
        RECT  0.715 0.185 0.735 0.305 ;
        RECT  0.695 0.980 0.735 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.525 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 -0.115 0.840 0.115 ;
        RECT  0.470 -0.115 0.590 0.275 ;
        RECT  0.140 -0.115 0.470 0.115 ;
        RECT  0.040 -0.115 0.140 0.275 ;
        RECT  0.000 -0.115 0.040 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.145 0.840 1.375 ;
        RECT  0.470 0.985 0.590 1.375 ;
        RECT  0.000 1.145 0.470 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.595 0.355 0.665 0.915 ;
        RECT  0.350 0.355 0.595 0.425 ;
        RECT  0.130 0.845 0.595 0.915 ;
        RECT  0.270 0.185 0.350 0.425 ;
        RECT  0.050 0.845 0.130 1.035 ;
    END
END OR2D1BWP40

MACRO OR2D2BWP40
    CLASS CORE ;
    FOREIGN OR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.355 0.815 0.905 ;
        RECT  0.715 0.355 0.735 0.435 ;
        RECT  0.715 0.785 0.735 0.905 ;
        RECT  0.645 0.215 0.715 0.435 ;
        RECT  0.645 0.785 0.715 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.390 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.210 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.115 0.980 0.115 ;
        RECT  0.830 -0.115 0.910 0.280 ;
        RECT  0.540 -0.115 0.830 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.145 0.980 1.375 ;
        RECT  0.830 0.980 0.910 1.375 ;
        RECT  0.550 1.145 0.830 1.375 ;
        RECT  0.410 1.050 0.550 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 0.520 0.620 0.640 ;
        RECT  0.470 0.345 0.540 0.915 ;
        RECT  0.320 0.345 0.470 0.415 ;
        RECT  0.145 0.845 0.470 0.915 ;
        RECT  0.220 0.185 0.320 0.415 ;
        RECT  0.035 0.845 0.145 1.075 ;
    END
END OR2D2BWP40

MACRO OR2D3BWP40
    CLASS CORE ;
    FOREIGN OR2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.268000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.195 1.205 0.475 ;
        RECT  1.135 0.785 1.205 1.075 ;
        RECT  1.015 0.785 1.135 0.905 ;
        RECT  1.015 0.355 1.130 0.475 ;
        RECT  0.805 0.355 1.015 0.905 ;
        RECT  0.755 0.355 0.805 0.475 ;
        RECT  0.745 0.785 0.805 0.905 ;
        RECT  0.665 0.195 0.755 0.475 ;
        RECT  0.675 0.785 0.745 1.075 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.390 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.205 0.640 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.990 -0.115 1.260 0.115 ;
        RECT  0.865 -0.115 0.990 0.280 ;
        RECT  0.540 -0.115 0.865 0.115 ;
        RECT  0.420 -0.115 0.540 0.275 ;
        RECT  0.130 -0.115 0.420 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 1.145 1.260 1.375 ;
        RECT  0.865 0.980 0.985 1.375 ;
        RECT  0.550 1.145 0.865 1.375 ;
        RECT  0.410 1.050 0.550 1.375 ;
        RECT  0.000 1.145 0.410 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.130 0.195 1.205 0.475 ;
        RECT  1.135 0.785 1.205 1.075 ;
        RECT  1.085 0.785 1.135 0.905 ;
        RECT  1.085 0.355 1.130 0.475 ;
        RECT  0.745 0.785 0.775 0.905 ;
        RECT  0.675 0.785 0.745 1.075 ;
        RECT  0.665 0.195 0.735 0.475 ;
        RECT  0.540 0.545 0.700 0.615 ;
        RECT  0.470 0.345 0.540 0.915 ;
        RECT  0.340 0.345 0.470 0.415 ;
        RECT  0.145 0.845 0.470 0.915 ;
        RECT  0.220 0.195 0.340 0.415 ;
        RECT  0.035 0.845 0.145 1.075 ;
    END
END OR2D3BWP40

MACRO OR2D4BWP40
    CLASS CORE ;
    FOREIGN OR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.820 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 0.185 1.515 0.480 ;
        RECT  1.445 0.695 1.515 1.025 ;
        RECT  1.435 0.350 1.445 0.480 ;
        RECT  1.435 0.695 1.445 0.815 ;
        RECT  1.225 0.350 1.435 0.815 ;
        RECT  1.135 0.350 1.225 0.470 ;
        RECT  1.135 0.695 1.225 0.815 ;
        RECT  1.065 0.185 1.135 0.470 ;
        RECT  1.065 0.695 1.135 1.025 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.510 0.780 0.630 ;
        RECT  0.625 0.510 0.695 0.780 ;
        RECT  0.245 0.710 0.625 0.780 ;
        RECT  0.170 0.495 0.245 0.780 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.115 1.820 0.115 ;
        RECT  1.655 -0.115 1.735 0.475 ;
        RECT  1.350 -0.115 1.655 0.115 ;
        RECT  1.230 -0.115 1.350 0.260 ;
        RECT  0.920 -0.115 1.230 0.115 ;
        RECT  0.840 -0.115 0.920 0.260 ;
        RECT  0.510 -0.115 0.840 0.115 ;
        RECT  0.430 -0.115 0.510 0.260 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.145 1.820 1.375 ;
        RECT  1.650 0.720 1.730 1.375 ;
        RECT  1.350 1.145 1.650 1.375 ;
        RECT  1.230 0.895 1.350 1.375 ;
        RECT  0.940 1.145 1.230 1.375 ;
        RECT  0.820 1.020 0.940 1.375 ;
        RECT  0.130 1.145 0.820 1.375 ;
        RECT  0.050 0.840 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.505 0.185 1.515 0.480 ;
        RECT  1.505 0.695 1.515 1.025 ;
        RECT  1.135 0.350 1.155 0.470 ;
        RECT  1.135 0.695 1.155 0.815 ;
        RECT  1.065 0.185 1.135 0.470 ;
        RECT  1.065 0.695 1.135 1.025 ;
        RECT  0.925 0.545 1.145 0.615 ;
        RECT  0.855 0.345 0.925 0.925 ;
        RECT  0.695 0.345 0.855 0.415 ;
        RECT  0.415 0.855 0.855 0.925 ;
        RECT  0.335 0.995 0.720 1.065 ;
        RECT  0.625 0.190 0.695 0.415 ;
        RECT  0.325 0.345 0.625 0.415 ;
        RECT  0.220 0.850 0.335 1.065 ;
        RECT  0.225 0.185 0.325 0.415 ;
    END
END OR2D4BWP40

MACRO OR2D6BWP40
    CLASS CORE ;
    FOREIGN OR2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.100 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.195 1.855 0.465 ;
        RECT  1.785 0.710 1.855 1.040 ;
        RECT  1.575 0.355 1.785 0.465 ;
        RECT  1.575 0.710 1.785 0.830 ;
        RECT  1.475 0.355 1.575 0.830 ;
        RECT  1.405 0.195 1.475 1.040 ;
        RECT  1.365 0.355 1.405 0.830 ;
        RECT  1.095 0.355 1.365 0.475 ;
        RECT  1.095 0.710 1.365 0.830 ;
        RECT  1.025 0.195 1.095 0.475 ;
        RECT  1.025 0.710 1.095 1.040 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.695 0.510 0.780 0.630 ;
        RECT  0.625 0.510 0.695 0.780 ;
        RECT  0.245 0.710 0.625 0.780 ;
        RECT  0.170 0.485 0.245 0.780 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.064000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.545 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.115 2.100 0.115 ;
        RECT  1.970 -0.115 2.050 0.425 ;
        RECT  1.690 -0.115 1.970 0.115 ;
        RECT  1.570 -0.115 1.690 0.270 ;
        RECT  1.310 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.310 0.270 ;
        RECT  0.900 -0.115 1.190 0.115 ;
        RECT  0.820 -0.115 0.900 0.260 ;
        RECT  0.510 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.510 0.260 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.395 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.145 2.100 1.375 ;
        RECT  1.965 0.720 2.045 1.375 ;
        RECT  1.690 1.145 1.965 1.375 ;
        RECT  1.570 0.905 1.690 1.375 ;
        RECT  1.310 1.145 1.570 1.375 ;
        RECT  1.190 0.905 1.310 1.375 ;
        RECT  0.920 1.145 1.190 1.375 ;
        RECT  0.800 1.015 0.920 1.375 ;
        RECT  0.130 1.145 0.800 1.375 ;
        RECT  0.050 0.840 0.130 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.785 0.195 1.855 0.465 ;
        RECT  1.025 0.195 1.095 0.475 ;
        RECT  1.025 0.710 1.095 1.040 ;
        RECT  1.645 0.545 1.985 0.615 ;
        RECT  0.925 0.545 1.255 0.615 ;
        RECT  0.855 0.330 0.925 0.925 ;
        RECT  0.720 0.330 0.855 0.400 ;
        RECT  0.415 0.855 0.855 0.925 ;
        RECT  0.600 0.195 0.720 0.400 ;
        RECT  0.335 0.995 0.720 1.065 ;
        RECT  0.340 0.330 0.600 0.400 ;
        RECT  0.220 0.195 0.340 0.400 ;
        RECT  0.225 0.850 0.335 1.065 ;
        RECT  1.785 0.710 1.855 1.040 ;
        RECT  1.645 0.355 1.785 0.465 ;
        RECT  1.645 0.710 1.785 0.830 ;
        RECT  1.095 0.355 1.295 0.475 ;
        RECT  1.095 0.710 1.295 0.830 ;
    END
END OR2D6BWP40

MACRO OR2D8BWP40
    CLASS CORE ;
    FOREIGN OR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.477000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.135 0.325 2.220 0.445 ;
        RECT  2.135 0.700 2.220 0.820 ;
        RECT  1.925 0.325 2.135 0.820 ;
        RECT  1.900 0.325 1.925 0.445 ;
        RECT  1.900 0.700 1.925 0.820 ;
        RECT  1.805 0.185 1.900 0.445 ;
        RECT  1.805 0.700 1.900 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.420 0.700 1.500 0.990 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.093600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.490 1.160 0.765 ;
        RECT  0.535 0.695 1.090 0.765 ;
        RECT  0.445 0.495 0.535 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.093600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.540 0.915 0.625 ;
        RECT  0.730 0.355 0.815 0.625 ;
        RECT  0.300 0.355 0.730 0.425 ;
        RECT  0.220 0.355 0.300 0.650 ;
        RECT  0.125 0.495 0.220 0.650 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 -0.115 2.940 0.115 ;
        RECT  2.810 -0.115 2.890 0.445 ;
        RECT  2.520 -0.115 2.810 0.115 ;
        RECT  2.400 -0.115 2.520 0.255 ;
        RECT  2.120 -0.115 2.400 0.115 ;
        RECT  2.000 -0.115 2.120 0.255 ;
        RECT  1.720 -0.115 2.000 0.115 ;
        RECT  1.600 -0.115 1.720 0.255 ;
        RECT  1.330 -0.115 1.600 0.115 ;
        RECT  1.190 -0.115 1.330 0.235 ;
        RECT  0.930 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.930 0.145 ;
        RECT  0.550 -0.115 0.810 0.115 ;
        RECT  0.410 -0.115 0.550 0.145 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.145 2.940 1.375 ;
        RECT  2.810 0.720 2.890 1.375 ;
        RECT  2.520 1.145 2.810 1.375 ;
        RECT  2.400 0.890 2.520 1.375 ;
        RECT  2.120 1.145 2.400 1.375 ;
        RECT  2.000 0.890 2.120 1.375 ;
        RECT  1.720 1.145 2.000 1.375 ;
        RECT  1.600 0.890 1.720 1.375 ;
        RECT  1.300 1.145 1.600 1.375 ;
        RECT  1.220 0.995 1.300 1.375 ;
        RECT  0.540 1.145 1.220 1.375 ;
        RECT  0.420 1.000 0.540 1.375 ;
        RECT  0.000 1.145 0.420 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.620 0.185 2.700 0.445 ;
        RECT  2.620 0.700 2.700 0.990 ;
        RECT  2.300 0.325 2.620 0.445 ;
        RECT  2.300 0.700 2.620 0.820 ;
        RECT  2.220 0.185 2.300 0.445 ;
        RECT  2.220 0.700 2.300 0.990 ;
        RECT  2.205 0.325 2.220 0.445 ;
        RECT  2.205 0.700 2.220 0.820 ;
        RECT  1.805 0.185 1.855 0.445 ;
        RECT  1.805 0.700 1.855 1.045 ;
        RECT  1.500 0.325 1.805 0.445 ;
        RECT  1.500 0.700 1.805 0.820 ;
        RECT  1.420 0.185 1.500 0.445 ;
        RECT  1.095 0.340 1.250 0.410 ;
        RECT  0.905 0.845 1.250 0.915 ;
        RECT  1.025 0.215 1.095 0.410 ;
        RECT  0.220 0.215 1.025 0.285 ;
        RECT  0.830 0.845 0.905 1.075 ;
        RECT  0.145 0.845 0.830 0.915 ;
        RECT  0.035 0.845 0.145 1.075 ;
        RECT  1.420 0.700 1.500 0.990 ;
        RECT  2.205 0.545 2.715 0.615 ;
        RECT  1.320 0.545 1.775 0.615 ;
        RECT  1.250 0.340 1.320 0.915 ;
    END
END OR2D8BWP40

MACRO OR3D0BWP40
    CLASS CORE ;
    FOREIGN OR3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.075 ;
        RECT  0.840 0.190 0.875 0.290 ;
        RECT  0.835 0.985 0.875 1.075 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.285 ;
        RECT  0.350 -0.115 0.640 0.115 ;
        RECT  0.230 -0.115 0.350 0.145 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.735 1.145 0.980 1.375 ;
        RECT  0.665 0.995 0.735 1.375 ;
        RECT  0.000 1.145 0.665 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.915 ;
        RECT  0.565 0.355 0.735 0.425 ;
        RECT  0.130 0.845 0.735 0.915 ;
        RECT  0.495 0.215 0.565 0.425 ;
        RECT  0.140 0.215 0.495 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
        RECT  0.060 0.845 0.130 1.040 ;
    END
END OR3D0BWP40

MACRO OR3D1BWP40
    CLASS CORE ;
    FOREIGN OR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.980 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.190 0.945 1.075 ;
        RECT  0.840 0.190 0.875 0.290 ;
        RECT  0.835 0.985 0.875 1.075 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.665 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.455 0.495 0.595 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 -0.115 0.980 0.115 ;
        RECT  0.640 -0.115 0.760 0.285 ;
        RECT  0.350 -0.115 0.640 0.115 ;
        RECT  0.230 -0.115 0.350 0.145 ;
        RECT  0.000 -0.115 0.230 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.145 0.980 1.375 ;
        RECT  0.660 0.995 0.740 1.375 ;
        RECT  0.000 1.145 0.660 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.355 0.805 0.915 ;
        RECT  0.565 0.355 0.735 0.425 ;
        RECT  0.130 0.845 0.735 0.915 ;
        RECT  0.495 0.215 0.565 0.425 ;
        RECT  0.140 0.215 0.495 0.285 ;
        RECT  0.040 0.185 0.140 0.285 ;
        RECT  0.060 0.845 0.130 1.040 ;
    END
END OR3D1BWP40

MACRO OR3D2BWP40
    CLASS CORE ;
    FOREIGN OR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.215 0.965 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.645 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.485 0.385 0.800 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 0.490 0.665 0.625 ;
        RECT  0.455 0.490 0.530 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.195 -0.115 1.260 0.115 ;
        RECT  1.115 -0.115 1.195 0.485 ;
        RECT  0.750 -0.115 1.115 0.115 ;
        RECT  0.630 -0.115 0.750 0.245 ;
        RECT  0.340 -0.115 0.630 0.115 ;
        RECT  0.220 -0.115 0.340 0.245 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.145 1.260 1.375 ;
        RECT  1.110 0.720 1.190 1.375 ;
        RECT  0.750 1.145 1.110 1.375 ;
        RECT  0.630 1.050 0.750 1.375 ;
        RECT  0.000 1.145 0.630 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.735 0.325 0.805 0.980 ;
        RECT  0.130 0.325 0.735 0.395 ;
        RECT  0.140 0.910 0.735 0.980 ;
        RECT  0.050 0.910 0.140 1.060 ;
        RECT  0.050 0.225 0.130 0.395 ;
    END
END OR3D2BWP40

MACRO OR3D3BWP40
    CLASS CORE ;
    FOREIGN OR3D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.236000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.195 1.365 0.475 ;
        RECT  1.295 0.760 1.365 1.055 ;
        RECT  1.270 0.195 1.295 1.055 ;
        RECT  1.265 0.365 1.270 1.055 ;
        RECT  1.085 0.365 1.265 0.915 ;
        RECT  0.955 0.365 1.085 0.475 ;
        RECT  0.955 0.760 1.085 0.915 ;
        RECT  0.885 0.195 0.955 0.475 ;
        RECT  0.885 0.760 0.955 1.055 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 0.495 0.385 0.785 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.545 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 -0.115 1.400 0.115 ;
        RECT  1.060 -0.115 1.180 0.270 ;
        RECT  0.750 -0.115 1.060 0.115 ;
        RECT  0.630 -0.115 0.750 0.270 ;
        RECT  0.340 -0.115 0.630 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.145 1.400 1.375 ;
        RECT  1.060 1.050 1.180 1.375 ;
        RECT  0.750 1.145 1.060 1.375 ;
        RECT  0.630 1.050 0.750 1.375 ;
        RECT  0.000 1.145 0.630 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.955 0.365 0.975 0.475 ;
        RECT  0.955 0.760 0.975 0.915 ;
        RECT  0.885 0.195 0.955 0.475 ;
        RECT  0.885 0.760 0.955 1.055 ;
        RECT  0.805 0.545 0.900 0.615 ;
        RECT  0.735 0.345 0.805 0.980 ;
        RECT  0.515 0.345 0.735 0.415 ;
        RECT  0.140 0.910 0.735 0.980 ;
        RECT  0.420 0.185 0.515 0.415 ;
        RECT  0.130 0.345 0.420 0.415 ;
        RECT  0.050 0.910 0.140 1.060 ;
        RECT  0.035 0.185 0.130 0.415 ;
    END
END OR3D3BWP40

MACRO OR3D4BWP40
    CLASS CORE ;
    FOREIGN OR3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.256000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.185 1.945 0.465 ;
        RECT  1.875 0.785 1.945 1.065 ;
        RECT  1.855 0.335 1.875 0.465 ;
        RECT  1.855 0.785 1.875 0.905 ;
        RECT  1.645 0.335 1.855 0.905 ;
        RECT  1.535 0.335 1.645 0.465 ;
        RECT  1.535 0.785 1.645 0.905 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.785 1.535 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.000 0.640 ;
        RECT  0.430 0.355 0.875 0.425 ;
        RECT  0.350 0.355 0.430 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.495 1.225 0.790 ;
        RECT  0.260 0.720 1.105 0.790 ;
        RECT  0.170 0.495 0.260 0.790 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 -0.115 2.240 0.115 ;
        RECT  2.090 -0.115 2.170 0.475 ;
        RECT  1.760 -0.115 2.090 0.115 ;
        RECT  1.640 -0.115 1.760 0.245 ;
        RECT  1.320 -0.115 1.640 0.115 ;
        RECT  1.240 -0.115 1.320 0.265 ;
        RECT  0.930 -0.115 1.240 0.115 ;
        RECT  0.810 -0.115 0.930 0.145 ;
        RECT  0.530 -0.115 0.810 0.115 ;
        RECT  0.410 -0.115 0.530 0.145 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.145 2.240 1.375 ;
        RECT  2.090 0.720 2.170 1.375 ;
        RECT  1.760 1.145 2.090 1.375 ;
        RECT  1.640 0.985 1.760 1.375 ;
        RECT  1.320 1.145 1.640 1.375 ;
        RECT  1.240 1.010 1.320 1.375 ;
        RECT  0.125 1.145 1.240 1.375 ;
        RECT  0.055 0.860 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.925 0.185 1.945 0.465 ;
        RECT  1.925 0.785 1.945 1.065 ;
        RECT  1.535 0.335 1.575 0.465 ;
        RECT  1.535 0.785 1.575 0.905 ;
        RECT  1.465 0.185 1.535 0.465 ;
        RECT  1.465 0.785 1.535 1.065 ;
        RECT  1.375 0.545 1.550 0.630 ;
        RECT  1.305 0.345 1.375 0.940 ;
        RECT  1.145 0.345 1.305 0.415 ;
        RECT  0.730 0.870 1.305 0.940 ;
        RECT  1.075 0.215 1.145 0.415 ;
        RECT  0.220 0.215 1.075 0.285 ;
        RECT  0.610 0.870 0.730 1.075 ;
    END
END OR3D4BWP40

MACRO OR3D6BWP40
    CLASS CORE ;
    FOREIGN OR3D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.360000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.185 2.275 0.465 ;
        RECT  2.205 0.695 2.275 1.065 ;
        RECT  1.995 0.355 2.205 0.465 ;
        RECT  1.995 0.695 2.205 0.815 ;
        RECT  1.895 0.355 1.995 0.815 ;
        RECT  1.825 0.185 1.895 1.065 ;
        RECT  1.785 0.355 1.825 0.815 ;
        RECT  1.495 0.355 1.785 0.465 ;
        RECT  1.495 0.695 1.785 0.815 ;
        RECT  1.425 0.185 1.495 0.465 ;
        RECT  1.425 0.695 1.495 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.805 0.625 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.355 1.000 0.645 ;
        RECT  0.430 0.355 0.875 0.425 ;
        RECT  0.350 0.355 0.430 0.645 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.105 0.495 1.185 0.790 ;
        RECT  0.260 0.720 1.105 0.790 ;
        RECT  0.170 0.495 0.260 0.790 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 -0.115 2.520 0.115 ;
        RECT  2.390 -0.115 2.470 0.475 ;
        RECT  2.110 -0.115 2.390 0.115 ;
        RECT  1.990 -0.115 2.110 0.275 ;
        RECT  1.720 -0.115 1.990 0.115 ;
        RECT  1.600 -0.115 1.720 0.275 ;
        RECT  1.300 -0.115 1.600 0.115 ;
        RECT  1.220 -0.115 1.300 0.265 ;
        RECT  0.930 -0.115 1.220 0.115 ;
        RECT  0.810 -0.115 0.930 0.145 ;
        RECT  0.530 -0.115 0.810 0.115 ;
        RECT  0.410 -0.115 0.530 0.145 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.145 2.520 1.375 ;
        RECT  2.390 0.720 2.470 1.375 ;
        RECT  2.110 1.145 2.390 1.375 ;
        RECT  1.990 0.895 2.110 1.375 ;
        RECT  1.720 1.145 1.990 1.375 ;
        RECT  1.600 0.895 1.720 1.375 ;
        RECT  1.290 1.145 1.600 1.375 ;
        RECT  1.210 1.000 1.290 1.375 ;
        RECT  0.125 1.145 1.210 1.375 ;
        RECT  0.055 0.865 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.205 0.185 2.275 0.465 ;
        RECT  2.205 0.695 2.275 1.065 ;
        RECT  2.065 0.355 2.205 0.465 ;
        RECT  2.065 0.695 2.205 0.815 ;
        RECT  1.495 0.355 1.715 0.465 ;
        RECT  1.495 0.695 1.715 0.815 ;
        RECT  1.425 0.185 1.495 0.465 ;
        RECT  1.425 0.695 1.495 1.065 ;
        RECT  2.075 0.545 2.410 0.615 ;
        RECT  1.335 0.545 1.710 0.615 ;
        RECT  1.265 0.345 1.335 0.930 ;
        RECT  1.145 0.345 1.265 0.415 ;
        RECT  0.725 0.860 1.265 0.930 ;
        RECT  1.075 0.215 1.145 0.415 ;
        RECT  0.220 0.215 1.075 0.285 ;
        RECT  0.615 0.860 0.725 1.075 ;
    END
END OR3D6BWP40

MACRO OR3D8BWP40
    CLASS CORE ;
    FOREIGN OR3D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.480000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 0.700 3.260 1.025 ;
        RECT  3.185 0.185 3.255 0.465 ;
        RECT  2.855 0.345 3.185 0.465 ;
        RECT  2.855 0.700 3.180 0.820 ;
        RECT  2.835 0.185 2.855 0.465 ;
        RECT  2.835 0.700 2.855 1.045 ;
        RECT  2.785 0.185 2.835 1.045 ;
        RECT  2.780 0.345 2.785 1.045 ;
        RECT  2.625 0.345 2.780 0.820 ;
        RECT  2.455 0.345 2.625 0.465 ;
        RECT  2.460 0.700 2.625 0.820 ;
        RECT  2.380 0.700 2.460 1.025 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.055 0.345 2.385 0.465 ;
        RECT  2.060 0.700 2.380 0.820 ;
        RECT  1.980 0.700 2.060 1.025 ;
        RECT  1.985 0.185 2.055 0.465 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 0.495 0.540 0.625 ;
        RECT  0.175 0.495 0.255 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.495 1.135 0.765 ;
        RECT  0.780 0.495 1.005 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.560 0.495 1.645 0.765 ;
        RECT  1.335 0.495 1.560 0.615 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 -0.115 3.500 0.115 ;
        RECT  3.370 -0.115 3.450 0.465 ;
        RECT  3.080 -0.115 3.370 0.115 ;
        RECT  2.960 -0.115 3.080 0.265 ;
        RECT  2.680 -0.115 2.960 0.115 ;
        RECT  2.560 -0.115 2.680 0.265 ;
        RECT  2.280 -0.115 2.560 0.115 ;
        RECT  2.160 -0.115 2.280 0.265 ;
        RECT  1.855 -0.115 2.160 0.115 ;
        RECT  1.775 -0.115 1.855 0.275 ;
        RECT  1.460 -0.115 1.775 0.115 ;
        RECT  1.380 -0.115 1.460 0.275 ;
        RECT  1.080 -0.115 1.380 0.115 ;
        RECT  1.000 -0.115 1.080 0.275 ;
        RECT  0.700 -0.115 1.000 0.115 ;
        RECT  0.620 -0.115 0.700 0.275 ;
        RECT  0.320 -0.115 0.620 0.115 ;
        RECT  0.240 -0.115 0.320 0.275 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.145 3.500 1.375 ;
        RECT  3.370 0.720 3.450 1.375 ;
        RECT  3.080 1.145 3.370 1.375 ;
        RECT  2.960 0.890 3.080 1.375 ;
        RECT  2.680 1.145 2.960 1.375 ;
        RECT  2.560 0.890 2.680 1.375 ;
        RECT  2.280 1.145 2.560 1.375 ;
        RECT  2.160 0.890 2.280 1.375 ;
        RECT  1.855 1.145 2.160 1.375 ;
        RECT  1.775 0.860 1.855 1.375 ;
        RECT  1.460 1.145 1.775 1.375 ;
        RECT  1.380 0.985 1.460 1.375 ;
        RECT  0.000 1.145 1.380 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.180 0.700 3.260 1.025 ;
        RECT  3.185 0.185 3.255 0.465 ;
        RECT  2.905 0.345 3.185 0.465 ;
        RECT  2.905 0.700 3.180 0.820 ;
        RECT  2.455 0.345 2.555 0.465 ;
        RECT  2.460 0.700 2.555 0.820 ;
        RECT  2.380 0.700 2.460 1.025 ;
        RECT  2.385 0.185 2.455 0.465 ;
        RECT  2.055 0.345 2.385 0.465 ;
        RECT  2.060 0.700 2.380 0.820 ;
        RECT  1.980 0.700 2.060 1.025 ;
        RECT  1.985 0.185 2.055 0.465 ;
        RECT  1.880 0.545 2.485 0.615 ;
        RECT  1.810 0.345 1.880 0.615 ;
        RECT  1.645 0.345 1.810 0.415 ;
        RECT  1.550 0.845 1.670 1.055 ;
        RECT  1.575 0.185 1.645 0.415 ;
        RECT  1.265 0.345 1.575 0.415 ;
        RECT  1.265 0.845 1.550 0.915 ;
        RECT  1.195 0.185 1.265 0.415 ;
        RECT  1.195 0.845 1.265 1.075 ;
        RECT  0.885 0.345 1.195 0.415 ;
        RECT  0.790 0.845 1.195 0.915 ;
        RECT  0.220 0.985 1.100 1.055 ;
        RECT  0.815 0.185 0.885 0.415 ;
        RECT  0.700 0.345 0.815 0.415 ;
        RECT  0.620 0.345 0.700 0.915 ;
        RECT  0.505 0.345 0.620 0.415 ;
        RECT  0.125 0.845 0.620 0.915 ;
        RECT  0.435 0.185 0.505 0.415 ;
        RECT  0.130 0.345 0.435 0.415 ;
        RECT  0.050 0.285 0.130 0.415 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END OR3D8BWP40

MACRO OR4D0BWP40
    CLASS CORE ;
    FOREIGN OR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.058000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.185 1.225 1.060 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.670 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.870 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.115 1.260 0.115 ;
        RECT  0.880 -0.115 1.000 0.250 ;
        RECT  0.565 -0.115 0.880 0.115 ;
        RECT  0.445 -0.115 0.565 0.140 ;
        RECT  0.130 -0.115 0.445 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.145 1.260 1.375 ;
        RECT  0.880 1.010 1.000 1.375 ;
        RECT  0.000 1.145 0.880 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.335 1.055 0.915 ;
        RECT  0.780 0.335 0.985 0.405 ;
        RECT  0.125 0.845 0.985 0.915 ;
        RECT  0.710 0.210 0.780 0.405 ;
        RECT  0.220 0.210 0.710 0.280 ;
        RECT  0.055 0.845 0.125 1.055 ;
    END
END OR4D0BWP40

MACRO OR4D1BWP40
    CLASS CORE ;
    FOREIGN OR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.260 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.116000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.185 1.225 1.060 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.385 0.670 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.025000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.870 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 -0.115 1.260 0.115 ;
        RECT  0.880 -0.115 1.000 0.250 ;
        RECT  0.565 -0.115 0.880 0.115 ;
        RECT  0.445 -0.115 0.565 0.140 ;
        RECT  0.130 -0.115 0.445 0.115 ;
        RECT  0.050 -0.115 0.130 0.315 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.145 1.260 1.375 ;
        RECT  0.880 1.010 1.000 1.375 ;
        RECT  0.000 1.145 0.880 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.335 1.055 0.915 ;
        RECT  0.780 0.335 0.985 0.405 ;
        RECT  0.135 0.845 0.985 0.915 ;
        RECT  0.710 0.210 0.780 0.405 ;
        RECT  0.220 0.210 0.710 0.280 ;
        RECT  0.050 0.845 0.135 1.010 ;
    END
END OR4D1BWP40

MACRO OR4D2BWP40
    CLASS CORE ;
    FOREIGN OR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.495 1.365 0.625 ;
        RECT  1.090 0.195 1.160 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.805 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.645 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.850 0.785 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.115 1.400 0.115 ;
        RECT  1.270 -0.115 1.345 0.425 ;
        RECT  0.980 -0.115 1.270 0.115 ;
        RECT  0.860 -0.115 0.980 0.275 ;
        RECT  0.550 -0.115 0.860 0.115 ;
        RECT  0.430 -0.115 0.550 0.275 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 1.145 1.400 1.375 ;
        RECT  1.275 0.715 1.345 1.375 ;
        RECT  0.970 1.145 1.275 1.375 ;
        RECT  0.850 1.050 0.970 1.375 ;
        RECT  0.000 1.145 0.850 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.345 1.020 0.980 ;
        RECT  0.750 0.345 0.950 0.415 ;
        RECT  0.035 0.910 0.950 0.980 ;
        RECT  0.670 0.185 0.750 0.415 ;
        RECT  0.320 0.345 0.670 0.415 ;
        RECT  0.225 0.185 0.320 0.415 ;
    END
END OR4D2BWP40

MACRO OR4D3BWP40
    CLASS CORE ;
    FOREIGN OR4D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.212000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.195 1.505 0.455 ;
        RECT  1.435 0.705 1.505 1.045 ;
        RECT  1.415 0.195 1.435 1.045 ;
        RECT  1.225 0.355 1.415 0.805 ;
        RECT  1.110 0.355 1.225 0.455 ;
        RECT  1.110 0.705 1.225 0.805 ;
        RECT  1.040 0.195 1.110 0.455 ;
        RECT  1.040 0.705 1.110 1.045 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.495 0.385 0.805 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.495 0.665 0.625 ;
        RECT  0.455 0.495 0.525 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.825 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.115 1.540 0.115 ;
        RECT  1.200 -0.115 1.320 0.275 ;
        RECT  0.930 -0.115 1.200 0.115 ;
        RECT  0.810 -0.115 0.930 0.275 ;
        RECT  0.530 -0.115 0.810 0.115 ;
        RECT  0.410 -0.115 0.530 0.275 ;
        RECT  0.130 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.130 0.415 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.540 1.375 ;
        RECT  1.200 0.905 1.320 1.375 ;
        RECT  0.930 1.145 1.200 1.375 ;
        RECT  0.810 1.050 0.930 1.375 ;
        RECT  0.000 1.145 0.810 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.110 0.355 1.155 0.455 ;
        RECT  1.110 0.705 1.155 0.805 ;
        RECT  1.040 0.195 1.110 0.455 ;
        RECT  1.040 0.705 1.110 1.045 ;
        RECT  0.970 0.545 1.075 0.615 ;
        RECT  0.900 0.345 0.970 0.960 ;
        RECT  0.700 0.345 0.900 0.415 ;
        RECT  0.035 0.890 0.900 0.960 ;
        RECT  0.620 0.185 0.700 0.415 ;
        RECT  0.320 0.345 0.620 0.415 ;
        RECT  0.225 0.185 0.320 0.415 ;
    END
END OR4D3BWP40

MACRO OR4D4BWP40
    CLASS CORE ;
    FOREIGN OR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.249600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.185 2.395 0.465 ;
        RECT  2.325 0.745 2.395 1.025 ;
        RECT  2.275 0.355 2.325 0.465 ;
        RECT  2.275 0.745 2.325 0.815 ;
        RECT  2.065 0.355 2.275 0.815 ;
        RECT  2.015 0.355 2.065 0.465 ;
        RECT  2.005 0.745 2.065 0.815 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.745 2.005 1.025 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.985 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.495 1.235 0.765 ;
        RECT  0.665 0.695 1.130 0.765 ;
        RECT  0.580 0.495 0.665 0.765 ;
        RECT  0.545 0.495 0.580 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.335 0.355 1.410 0.765 ;
        RECT  0.420 0.355 1.335 0.425 ;
        RECT  0.315 0.355 0.420 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.520 1.650 0.915 ;
        RECT  0.245 0.845 1.565 0.915 ;
        RECT  0.165 0.495 0.245 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 -0.115 2.660 0.115 ;
        RECT  2.530 -0.115 2.610 0.475 ;
        RECT  2.230 -0.115 2.530 0.115 ;
        RECT  2.110 -0.115 2.230 0.275 ;
        RECT  1.780 -0.115 2.110 0.115 ;
        RECT  1.700 -0.115 1.780 0.300 ;
        RECT  1.360 -0.115 1.700 0.115 ;
        RECT  1.240 -0.115 1.360 0.140 ;
        RECT  0.940 -0.115 1.240 0.115 ;
        RECT  0.820 -0.115 0.940 0.145 ;
        RECT  0.530 -0.115 0.820 0.115 ;
        RECT  0.410 -0.115 0.530 0.145 ;
        RECT  0.125 -0.115 0.410 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.660 1.375 ;
        RECT  2.530 0.700 2.610 1.375 ;
        RECT  2.230 1.145 2.530 1.375 ;
        RECT  2.110 0.890 2.230 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.125 1.800 1.375 ;
        RECT  0.125 1.145 1.680 1.375 ;
        RECT  0.055 0.980 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.345 0.185 2.395 0.465 ;
        RECT  2.345 0.745 2.395 1.025 ;
        RECT  1.945 0.185 1.995 0.465 ;
        RECT  1.935 0.745 1.995 1.025 ;
        RECT  1.855 0.545 1.985 0.635 ;
        RECT  1.785 0.370 1.855 1.055 ;
        RECT  1.600 0.370 1.785 0.440 ;
        RECT  0.820 0.985 1.785 1.055 ;
        RECT  1.530 0.215 1.600 0.440 ;
        RECT  0.220 0.215 1.530 0.285 ;
    END
END OR4D4BWP40

MACRO OR4D6BWP40
    CLASS CORE ;
    FOREIGN OR4D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.366600 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.185 2.780 0.470 ;
        RECT  2.700 0.745 2.780 1.025 ;
        RECT  2.415 0.355 2.700 0.470 ;
        RECT  2.415 0.745 2.700 0.815 ;
        RECT  2.405 0.355 2.415 0.815 ;
        RECT  2.400 0.185 2.405 0.815 ;
        RECT  2.325 0.185 2.400 1.025 ;
        RECT  2.205 0.355 2.325 0.815 ;
        RECT  2.015 0.355 2.205 0.465 ;
        RECT  2.005 0.745 2.205 0.815 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.745 2.005 1.025 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.735 0.495 0.985 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.495 1.225 0.765 ;
        RECT  0.665 0.695 1.120 0.765 ;
        RECT  0.595 0.495 0.665 0.765 ;
        RECT  0.570 0.495 0.595 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.355 1.430 0.765 ;
        RECT  0.440 0.355 1.295 0.425 ;
        RECT  0.315 0.355 0.440 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.565 0.520 1.650 0.915 ;
        RECT  0.245 0.845 1.565 0.915 ;
        RECT  0.145 0.495 0.245 0.915 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 -0.115 3.080 0.115 ;
        RECT  2.915 -0.115 2.995 0.475 ;
        RECT  2.610 -0.115 2.915 0.115 ;
        RECT  2.490 -0.115 2.610 0.275 ;
        RECT  2.230 -0.115 2.490 0.115 ;
        RECT  2.110 -0.115 2.230 0.275 ;
        RECT  1.780 -0.115 2.110 0.115 ;
        RECT  1.700 -0.115 1.780 0.300 ;
        RECT  1.360 -0.115 1.700 0.115 ;
        RECT  1.240 -0.115 1.360 0.140 ;
        RECT  0.940 -0.115 1.240 0.115 ;
        RECT  0.820 -0.115 0.940 0.145 ;
        RECT  0.550 -0.115 0.820 0.115 ;
        RECT  0.430 -0.115 0.550 0.145 ;
        RECT  0.125 -0.115 0.430 0.115 ;
        RECT  0.055 -0.115 0.125 0.420 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 1.145 3.080 1.375 ;
        RECT  2.915 0.700 2.995 1.375 ;
        RECT  2.610 1.145 2.915 1.375 ;
        RECT  2.490 0.885 2.610 1.375 ;
        RECT  2.230 1.145 2.490 1.375 ;
        RECT  2.110 0.885 2.230 1.375 ;
        RECT  1.800 1.145 2.110 1.375 ;
        RECT  1.680 1.125 1.800 1.375 ;
        RECT  0.125 1.145 1.680 1.375 ;
        RECT  0.055 1.000 0.125 1.375 ;
        RECT  0.000 1.145 0.055 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.700 0.185 2.780 0.470 ;
        RECT  2.700 0.745 2.780 1.025 ;
        RECT  2.485 0.355 2.700 0.470 ;
        RECT  2.485 0.745 2.700 0.815 ;
        RECT  2.015 0.355 2.135 0.465 ;
        RECT  2.005 0.745 2.135 0.815 ;
        RECT  1.945 0.185 2.015 0.465 ;
        RECT  1.935 0.745 2.005 1.025 ;
        RECT  1.855 0.545 2.130 0.615 ;
        RECT  1.785 0.370 1.855 1.055 ;
        RECT  1.600 0.370 1.785 0.440 ;
        RECT  0.815 0.985 1.785 1.055 ;
        RECT  1.530 0.215 1.600 0.440 ;
        RECT  0.240 0.215 1.530 0.285 ;
    END
END OR4D6BWP40

MACRO OR4D8BWP40
    CLASS CORE ;
    FOREIGN OR4D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.496000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.660 0.695 3.740 0.995 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.355 0.345 3.665 0.465 ;
        RECT  3.360 0.695 3.660 0.815 ;
        RECT  3.280 0.695 3.360 0.995 ;
        RECT  3.285 0.185 3.355 0.465 ;
        RECT  3.255 0.345 3.285 0.465 ;
        RECT  3.255 0.695 3.280 0.815 ;
        RECT  3.045 0.345 3.255 0.815 ;
        RECT  2.975 0.345 3.045 0.465 ;
        RECT  2.975 0.695 3.045 0.815 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.900 0.695 2.975 0.995 ;
        RECT  2.595 0.345 2.905 0.465 ;
        RECT  2.600 0.695 2.900 0.815 ;
        RECT  2.520 0.695 2.600 0.995 ;
        RECT  2.525 0.185 2.595 0.465 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.495 0.525 0.765 ;
        RECT  0.175 0.495 0.440 0.625 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 0.495 1.135 0.625 ;
        RECT  0.735 0.495 0.820 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.495 1.785 0.765 ;
        RECT  1.365 0.495 1.705 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.096000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.205 0.765 ;
        RECT  1.855 0.495 2.125 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.975 -0.115 4.060 0.115 ;
        RECT  3.895 -0.115 3.975 0.465 ;
        RECT  3.570 -0.115 3.895 0.115 ;
        RECT  3.450 -0.115 3.570 0.275 ;
        RECT  3.190 -0.115 3.450 0.115 ;
        RECT  3.070 -0.115 3.190 0.275 ;
        RECT  2.810 -0.115 3.070 0.115 ;
        RECT  2.690 -0.115 2.810 0.275 ;
        RECT  2.410 -0.115 2.690 0.115 ;
        RECT  2.330 -0.115 2.410 0.275 ;
        RECT  2.030 -0.115 2.330 0.115 ;
        RECT  1.950 -0.115 2.030 0.275 ;
        RECT  1.650 -0.115 1.950 0.115 ;
        RECT  1.570 -0.115 1.650 0.275 ;
        RECT  1.270 -0.115 1.570 0.115 ;
        RECT  1.190 -0.115 1.270 0.275 ;
        RECT  0.890 -0.115 1.190 0.115 ;
        RECT  0.810 -0.115 0.890 0.275 ;
        RECT  0.510 -0.115 0.810 0.115 ;
        RECT  0.430 -0.115 0.510 0.275 ;
        RECT  0.130 -0.115 0.430 0.115 ;
        RECT  0.050 -0.115 0.130 0.400 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.985 1.145 4.060 1.375 ;
        RECT  3.875 0.720 3.985 1.375 ;
        RECT  3.570 1.145 3.875 1.375 ;
        RECT  3.450 0.885 3.570 1.375 ;
        RECT  3.190 1.145 3.450 1.375 ;
        RECT  3.070 0.885 3.190 1.375 ;
        RECT  2.810 1.145 3.070 1.375 ;
        RECT  2.690 0.885 2.810 1.375 ;
        RECT  2.410 1.145 2.690 1.375 ;
        RECT  2.330 0.805 2.410 1.375 ;
        RECT  2.030 1.145 2.330 1.375 ;
        RECT  1.950 0.985 2.030 1.375 ;
        RECT  0.000 1.145 1.950 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.660 0.695 3.740 0.995 ;
        RECT  3.665 0.185 3.735 0.465 ;
        RECT  3.355 0.345 3.665 0.465 ;
        RECT  3.360 0.695 3.660 0.815 ;
        RECT  3.325 0.695 3.360 0.995 ;
        RECT  3.325 0.185 3.355 0.465 ;
        RECT  2.905 0.185 2.975 0.465 ;
        RECT  2.900 0.695 2.975 0.995 ;
        RECT  2.595 0.345 2.905 0.465 ;
        RECT  2.600 0.695 2.900 0.815 ;
        RECT  2.520 0.695 2.600 0.995 ;
        RECT  2.525 0.185 2.595 0.465 ;
        RECT  2.400 0.545 2.965 0.615 ;
        RECT  2.320 0.345 2.400 0.615 ;
        RECT  2.240 0.345 2.320 0.415 ;
        RECT  2.120 0.205 2.240 0.415 ;
        RECT  2.120 0.845 2.240 1.055 ;
        RECT  1.860 0.345 2.120 0.415 ;
        RECT  1.840 0.845 2.120 0.915 ;
        RECT  1.740 0.205 1.860 0.415 ;
        RECT  1.760 0.845 1.840 1.055 ;
        RECT  1.360 0.985 1.760 1.055 ;
        RECT  1.480 0.345 1.740 0.415 ;
        RECT  1.270 0.845 1.670 0.915 ;
        RECT  1.360 0.205 1.480 0.415 ;
        RECT  1.100 0.345 1.360 0.415 ;
        RECT  1.195 0.685 1.270 0.915 ;
        RECT  0.790 0.845 1.195 0.915 ;
        RECT  0.980 0.205 1.100 0.415 ;
        RECT  0.225 0.985 1.100 1.055 ;
        RECT  0.720 0.345 0.980 0.415 ;
        RECT  0.665 0.205 0.720 0.415 ;
        RECT  0.600 0.205 0.665 0.915 ;
        RECT  0.595 0.345 0.600 0.915 ;
        RECT  0.340 0.345 0.595 0.415 ;
        RECT  0.145 0.845 0.595 0.915 ;
        RECT  0.220 0.205 0.340 0.415 ;
        RECT  0.035 0.845 0.145 1.075 ;
    END
END OR4D8BWP40

MACRO SDFCNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.300 4.865 1.050 ;
        RECT  4.775 0.300 4.795 0.445 ;
        RECT  4.775 0.910 4.795 1.050 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.420 0.525 4.510 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.660 -0.115 4.900 0.115 ;
        RECT  4.580 -0.115 4.660 0.235 ;
        RECT  4.050 -0.115 4.580 0.115 ;
        RECT  3.980 -0.115 4.050 0.435 ;
        RECT  3.100 -0.115 3.980 0.115 ;
        RECT  3.005 -0.115 3.100 0.330 ;
        RECT  2.680 -0.115 3.005 0.115 ;
        RECT  2.610 -0.115 2.680 0.270 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.145 4.900 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.230 1.145 4.560 1.375 ;
        RECT  4.160 1.005 4.230 1.375 ;
        RECT  4.050 1.145 4.160 1.375 ;
        RECT  3.980 1.005 4.050 1.375 ;
        RECT  3.225 1.145 3.980 1.375 ;
        RECT  3.105 0.920 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.305 4.705 0.920 ;
        RECT  4.200 0.305 4.635 0.375 ;
        RECT  4.480 0.850 4.635 0.920 ;
        RECT  4.330 0.495 4.525 0.765 ;
        RECT  4.410 0.850 4.480 1.075 ;
        RECT  4.335 1.005 4.410 1.075 ;
        RECT  3.665 0.845 4.325 0.915 ;
        RECT  4.130 0.305 4.200 0.735 ;
        RECT  3.885 0.665 4.130 0.735 ;
        RECT  3.755 0.695 3.800 0.765 ;
        RECT  3.685 0.195 3.755 0.765 ;
        RECT  3.305 0.195 3.685 0.265 ;
        RECT  3.595 0.845 3.665 1.025 ;
        RECT  3.565 0.345 3.595 1.025 ;
        RECT  3.520 0.345 3.565 0.915 ;
        RECT  3.180 0.410 3.250 0.840 ;
        RECT  2.865 0.410 3.180 0.490 ;
        RECT  2.395 0.770 3.180 0.840 ;
        RECT  2.720 0.570 3.100 0.640 ;
        RECT  2.790 0.340 2.865 0.490 ;
        RECT  2.650 0.340 2.720 0.640 ;
        RECT  2.190 0.920 2.705 0.990 ;
        RECT  2.490 0.340 2.650 0.410 ;
        RECT  2.465 0.490 2.580 0.690 ;
        RECT  2.420 0.195 2.490 0.410 ;
        RECT  2.090 0.195 2.420 0.265 ;
        RECT  2.295 0.635 2.395 0.840 ;
        RECT  2.195 0.340 2.295 0.555 ;
        RECT  2.190 0.485 2.195 0.555 ;
        RECT  2.120 0.485 2.190 0.990 ;
        RECT  2.020 0.195 2.090 0.405 ;
        RECT  2.000 0.195 2.020 0.960 ;
        RECT  1.950 0.335 2.000 0.960 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.805 0.875 1.860 0.945 ;
        RECT  1.735 0.875 1.805 1.055 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  0.715 0.985 1.735 1.055 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.660 0.725 1.705 0.795 ;
        RECT  1.580 0.725 1.660 0.890 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.375 0.525 4.445 0.595 ;
        RECT  2.500 0.525 2.570 0.595 ;
    END
END SDFCNQD0BWP40

MACRO SDFCNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.075 ;
        RECT  4.775 0.185 4.795 0.465 ;
        RECT  4.775 0.735 4.795 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.440 0.525 4.500 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 -0.115 4.900 0.115 ;
        RECT  4.550 -0.115 4.680 0.255 ;
        RECT  4.050 -0.115 4.550 0.115 ;
        RECT  3.980 -0.115 4.050 0.435 ;
        RECT  3.100 -0.115 3.980 0.115 ;
        RECT  2.980 -0.115 3.100 0.290 ;
        RECT  2.680 -0.115 2.980 0.115 ;
        RECT  2.610 -0.115 2.680 0.255 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.145 4.900 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.230 1.145 4.560 1.375 ;
        RECT  4.160 1.005 4.230 1.375 ;
        RECT  4.050 1.145 4.160 1.375 ;
        RECT  3.980 1.005 4.050 1.375 ;
        RECT  3.225 1.145 3.980 1.375 ;
        RECT  3.105 0.940 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.335 4.705 0.920 ;
        RECT  4.200 0.335 4.635 0.405 ;
        RECT  4.480 0.850 4.635 0.920 ;
        RECT  4.330 0.495 4.525 0.765 ;
        RECT  4.410 0.850 4.480 1.075 ;
        RECT  4.335 1.005 4.410 1.075 ;
        RECT  3.595 0.845 4.325 0.915 ;
        RECT  4.130 0.335 4.200 0.735 ;
        RECT  3.885 0.665 4.130 0.735 ;
        RECT  3.755 0.695 3.800 0.765 ;
        RECT  3.685 0.195 3.755 0.765 ;
        RECT  3.340 0.195 3.685 0.265 ;
        RECT  3.520 0.345 3.595 0.915 ;
        RECT  3.200 0.370 3.270 0.850 ;
        RECT  2.875 0.370 3.200 0.440 ;
        RECT  2.395 0.780 3.200 0.850 ;
        RECT  2.725 0.540 3.110 0.625 ;
        RECT  2.795 0.310 2.875 0.440 ;
        RECT  2.655 0.335 2.725 0.625 ;
        RECT  2.190 0.920 2.705 0.990 ;
        RECT  2.495 0.335 2.655 0.405 ;
        RECT  2.465 0.480 2.585 0.710 ;
        RECT  2.425 0.195 2.495 0.405 ;
        RECT  2.100 0.195 2.425 0.265 ;
        RECT  2.290 0.635 2.395 0.850 ;
        RECT  2.200 0.345 2.300 0.560 ;
        RECT  2.190 0.490 2.200 0.560 ;
        RECT  2.120 0.490 2.190 0.990 ;
        RECT  2.020 0.195 2.100 0.405 ;
        RECT  2.000 0.195 2.020 0.960 ;
        RECT  1.950 0.335 2.000 0.960 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.380 0.525 4.450 0.595 ;
        RECT  2.490 0.525 2.560 0.595 ;
    END
END SDFCNQD1BWP40

MACRO SDFCNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.144300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.420 0.525 4.515 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 -0.115 5.180 0.115 ;
        RECT  5.030 -0.115 5.105 0.480 ;
        RECT  4.680 -0.115 5.030 0.115 ;
        RECT  4.550 -0.115 4.680 0.255 ;
        RECT  4.050 -0.115 4.550 0.115 ;
        RECT  3.980 -0.115 4.050 0.435 ;
        RECT  3.120 -0.115 3.980 0.115 ;
        RECT  3.000 -0.115 3.120 0.235 ;
        RECT  2.680 -0.115 3.000 0.115 ;
        RECT  2.610 -0.115 2.680 0.290 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 1.145 5.180 1.375 ;
        RECT  5.030 0.655 5.105 1.375 ;
        RECT  4.680 1.145 5.030 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.230 1.145 4.560 1.375 ;
        RECT  4.160 1.005 4.230 1.375 ;
        RECT  4.050 1.145 4.160 1.375 ;
        RECT  3.980 1.005 4.050 1.375 ;
        RECT  3.225 1.145 3.980 1.375 ;
        RECT  3.105 0.920 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.335 4.705 0.920 ;
        RECT  4.200 0.335 4.635 0.405 ;
        RECT  4.480 0.850 4.635 0.920 ;
        RECT  4.330 0.495 4.525 0.765 ;
        RECT  4.410 0.850 4.480 1.075 ;
        RECT  4.335 1.005 4.410 1.075 ;
        RECT  3.595 0.845 4.325 0.915 ;
        RECT  4.130 0.335 4.200 0.735 ;
        RECT  3.885 0.665 4.130 0.735 ;
        RECT  3.755 0.695 3.800 0.765 ;
        RECT  3.685 0.195 3.755 0.765 ;
        RECT  3.310 0.195 3.685 0.265 ;
        RECT  3.520 0.345 3.595 0.915 ;
        RECT  3.275 0.335 3.345 0.840 ;
        RECT  2.800 0.335 3.275 0.405 ;
        RECT  2.350 0.770 3.275 0.840 ;
        RECT  2.730 0.545 3.150 0.615 ;
        RECT  2.660 0.360 2.730 0.615 ;
        RECT  2.190 0.920 2.725 0.990 ;
        RECT  2.530 0.360 2.660 0.430 ;
        RECT  2.430 0.510 2.590 0.690 ;
        RECT  2.460 0.195 2.530 0.430 ;
        RECT  2.090 0.195 2.460 0.265 ;
        RECT  2.270 0.615 2.350 0.840 ;
        RECT  2.195 0.335 2.295 0.545 ;
        RECT  2.190 0.475 2.195 0.545 ;
        RECT  2.120 0.475 2.190 0.990 ;
        RECT  2.020 0.195 2.090 0.405 ;
        RECT  2.000 0.195 2.020 0.960 ;
        RECT  1.950 0.335 2.000 0.960 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.385 0.525 4.455 0.595 ;
        RECT  2.480 0.525 2.550 0.595 ;
    END
END SDFCNQD2BWP40

MACRO SDFCNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.264900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.745 5.860 1.000 ;
        RECT  5.775 0.205 5.850 0.485 ;
        RECT  5.765 0.205 5.775 1.000 ;
        RECT  5.750 0.355 5.765 1.000 ;
        RECT  5.565 0.355 5.750 0.830 ;
        RECT  5.460 0.355 5.565 0.485 ;
        RECT  5.460 0.710 5.565 0.830 ;
        RECT  5.380 0.205 5.460 0.485 ;
        RECT  5.380 0.710 5.460 1.000 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.050600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.395 0.525 4.875 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.090 -0.115 6.160 0.115 ;
        RECT  6.020 -0.115 6.090 0.480 ;
        RECT  5.645 -0.115 6.020 0.115 ;
        RECT  5.570 -0.115 5.645 0.275 ;
        RECT  5.290 -0.115 5.570 0.115 ;
        RECT  5.155 -0.115 5.290 0.140 ;
        RECT  4.890 -0.115 5.155 0.115 ;
        RECT  4.755 -0.115 4.890 0.140 ;
        RECT  4.070 -0.115 4.755 0.115 ;
        RECT  4.000 -0.115 4.070 0.435 ;
        RECT  3.100 -0.115 4.000 0.115 ;
        RECT  2.980 -0.115 3.100 0.235 ;
        RECT  2.680 -0.115 2.980 0.115 ;
        RECT  2.610 -0.115 2.680 0.255 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.090 1.145 6.160 1.375 ;
        RECT  6.020 0.710 6.090 1.375 ;
        RECT  5.640 1.145 6.020 1.375 ;
        RECT  5.570 0.960 5.640 1.375 ;
        RECT  5.260 1.145 5.570 1.375 ;
        RECT  5.185 1.000 5.260 1.375 ;
        RECT  4.670 1.145 5.185 1.375 ;
        RECT  4.550 1.025 4.670 1.375 ;
        RECT  4.260 1.145 4.550 1.375 ;
        RECT  4.170 0.995 4.260 1.375 ;
        RECT  4.070 1.145 4.170 1.375 ;
        RECT  4.000 0.920 4.070 1.375 ;
        RECT  3.225 1.145 4.000 1.375 ;
        RECT  3.105 0.925 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.845 0.745 5.860 1.000 ;
        RECT  5.845 0.205 5.850 0.485 ;
        RECT  5.460 0.355 5.495 0.485 ;
        RECT  5.460 0.710 5.495 0.830 ;
        RECT  5.380 0.205 5.460 0.485 ;
        RECT  5.380 0.710 5.460 1.000 ;
        RECT  5.235 0.210 5.310 0.925 ;
        RECT  4.360 0.210 5.235 0.280 ;
        RECT  4.270 0.855 5.235 0.925 ;
        RECT  4.150 0.370 5.070 0.440 ;
        RECT  4.660 0.520 4.920 0.675 ;
        RECT  3.595 0.570 4.475 0.640 ;
        RECT  4.200 0.720 4.270 0.925 ;
        RECT  3.895 0.720 4.200 0.790 ;
        RECT  3.390 0.995 3.820 1.065 ;
        RECT  3.595 0.845 3.670 0.915 ;
        RECT  3.520 0.345 3.595 0.915 ;
        RECT  3.390 0.195 3.470 0.265 ;
        RECT  3.320 0.195 3.390 1.065 ;
        RECT  3.130 0.335 3.200 0.840 ;
        RECT  2.765 0.335 3.130 0.405 ;
        RECT  2.355 0.770 3.130 0.840 ;
        RECT  2.695 0.545 3.050 0.615 ;
        RECT  2.190 0.920 2.705 0.990 ;
        RECT  2.625 0.325 2.695 0.615 ;
        RECT  2.530 0.325 2.625 0.395 ;
        RECT  2.430 0.485 2.550 0.700 ;
        RECT  2.460 0.195 2.530 0.395 ;
        RECT  2.090 0.195 2.460 0.265 ;
        RECT  2.285 0.625 2.355 0.840 ;
        RECT  2.195 0.335 2.300 0.545 ;
        RECT  2.190 0.475 2.195 0.545 ;
        RECT  2.120 0.475 2.190 0.990 ;
        RECT  2.020 0.195 2.090 0.405 ;
        RECT  2.000 0.195 2.020 0.960 ;
        RECT  1.950 0.335 2.000 0.960 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.745 0.525 4.815 0.595 ;
        RECT  2.455 0.525 2.525 0.595 ;
    END
END SDFCNQD4BWP40

MACRO SDFCNQND0BWP40
    CLASS CORE ;
    FOREIGN SDFCNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.050 ;
        RECT  4.775 0.185 4.795 0.330 ;
        RECT  4.775 0.905 4.795 1.050 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.245 0.525 4.245 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.655 -0.115 4.900 0.115 ;
        RECT  4.585 -0.115 4.655 0.290 ;
        RECT  4.080 -0.115 4.585 0.115 ;
        RECT  3.945 -0.115 4.080 0.225 ;
        RECT  3.125 -0.115 3.945 0.115 ;
        RECT  3.005 -0.115 3.125 0.235 ;
        RECT  2.680 -0.115 3.005 0.115 ;
        RECT  2.610 -0.115 2.680 0.410 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.145 4.900 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.240 1.145 4.560 1.375 ;
        RECT  4.170 1.025 4.240 1.375 ;
        RECT  4.040 1.145 4.170 1.375 ;
        RECT  3.970 1.025 4.040 1.375 ;
        RECT  3.225 1.145 3.970 1.375 ;
        RECT  3.105 0.920 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.705 0.520 4.710 0.660 ;
        RECT  4.635 0.520 4.705 0.955 ;
        RECT  4.320 0.885 4.635 0.955 ;
        RECT  4.390 0.325 4.460 0.805 ;
        RECT  3.965 0.325 4.390 0.395 ;
        RECT  4.250 0.705 4.320 0.955 ;
        RECT  4.045 0.480 4.265 0.635 ;
        RECT  3.825 0.705 4.250 0.775 ;
        RECT  3.650 0.855 4.180 0.925 ;
        RECT  3.895 0.325 3.965 0.600 ;
        RECT  3.755 0.325 3.825 0.775 ;
        RECT  3.375 0.995 3.775 1.065 ;
        RECT  3.535 0.785 3.650 0.925 ;
        RECT  3.465 0.345 3.535 0.925 ;
        RECT  3.375 0.195 3.480 0.265 ;
        RECT  3.305 0.195 3.375 1.065 ;
        RECT  3.155 0.315 3.225 0.840 ;
        RECT  2.790 0.315 3.155 0.385 ;
        RECT  2.595 0.770 3.155 0.840 ;
        RECT  2.955 0.490 3.070 0.630 ;
        RECT  2.540 0.490 2.955 0.560 ;
        RECT  2.205 0.920 2.735 0.990 ;
        RECT  2.515 0.630 2.595 0.840 ;
        RECT  2.470 0.195 2.540 0.560 ;
        RECT  2.065 0.195 2.470 0.265 ;
        RECT  2.275 0.495 2.400 0.745 ;
        RECT  2.205 0.345 2.305 0.415 ;
        RECT  2.135 0.345 2.205 0.990 ;
        RECT  2.020 0.195 2.065 0.435 ;
        RECT  1.975 0.195 2.020 0.960 ;
        RECT  1.950 0.335 1.975 0.960 ;
        RECT  0.640 0.195 1.895 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.345 1.775 0.795 ;
        RECT  1.590 0.345 1.705 0.415 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.125 0.525 4.195 0.595 ;
        RECT  2.305 0.525 2.375 0.595 ;
    END
END SDFCNQND0BWP40

MACRO SDFCNQND1BWP40
    CLASS CORE ;
    FOREIGN SDFCNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.075 ;
        RECT  4.775 0.185 4.795 0.465 ;
        RECT  4.775 0.735 4.795 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.225 0.525 4.255 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.655 -0.115 4.900 0.115 ;
        RECT  4.585 -0.115 4.655 0.390 ;
        RECT  4.050 -0.115 4.585 0.115 ;
        RECT  3.980 -0.115 4.050 0.285 ;
        RECT  3.125 -0.115 3.980 0.115 ;
        RECT  3.005 -0.115 3.125 0.235 ;
        RECT  2.680 -0.115 3.005 0.115 ;
        RECT  2.610 -0.115 2.680 0.405 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.145 4.900 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.240 1.145 4.560 1.375 ;
        RECT  4.170 1.025 4.240 1.375 ;
        RECT  4.040 1.145 4.170 1.375 ;
        RECT  3.970 1.025 4.040 1.375 ;
        RECT  3.225 1.145 3.970 1.375 ;
        RECT  3.105 0.930 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.705 0.520 4.710 0.660 ;
        RECT  4.635 0.520 4.705 0.955 ;
        RECT  4.320 0.885 4.635 0.955 ;
        RECT  4.390 0.355 4.460 0.805 ;
        RECT  3.990 0.355 4.390 0.425 ;
        RECT  4.250 0.705 4.320 0.955 ;
        RECT  4.070 0.510 4.310 0.635 ;
        RECT  3.825 0.705 4.250 0.775 ;
        RECT  3.650 0.855 4.180 0.925 ;
        RECT  3.920 0.355 3.990 0.615 ;
        RECT  3.755 0.325 3.825 0.775 ;
        RECT  3.375 0.995 3.775 1.065 ;
        RECT  3.535 0.785 3.650 0.925 ;
        RECT  3.465 0.345 3.535 0.925 ;
        RECT  3.375 0.195 3.480 0.265 ;
        RECT  3.305 0.195 3.375 1.065 ;
        RECT  3.150 0.315 3.220 0.840 ;
        RECT  2.790 0.315 3.150 0.385 ;
        RECT  2.590 0.770 3.150 0.840 ;
        RECT  2.955 0.485 3.070 0.630 ;
        RECT  2.540 0.485 2.955 0.555 ;
        RECT  2.205 0.920 2.730 0.990 ;
        RECT  2.515 0.625 2.590 0.840 ;
        RECT  2.470 0.195 2.540 0.555 ;
        RECT  2.065 0.195 2.470 0.265 ;
        RECT  2.275 0.485 2.390 0.760 ;
        RECT  2.205 0.335 2.315 0.405 ;
        RECT  2.135 0.335 2.205 0.990 ;
        RECT  2.020 0.195 2.065 0.435 ;
        RECT  1.975 0.195 2.020 0.960 ;
        RECT  1.950 0.335 1.975 0.960 ;
        RECT  0.640 0.195 1.895 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.135 0.525 4.205 0.595 ;
        RECT  2.300 0.525 2.370 0.595 ;
    END
END SDFCNQND1BWP40

MACRO SDFCNQND2BWP40
    CLASS CORE ;
    FOREIGN SDFCNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.036000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.240 0.525 4.270 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 -0.115 5.180 0.115 ;
        RECT  5.035 -0.115 5.105 0.475 ;
        RECT  4.655 -0.115 5.035 0.115 ;
        RECT  4.585 -0.115 4.655 0.390 ;
        RECT  4.050 -0.115 4.585 0.115 ;
        RECT  3.980 -0.115 4.050 0.285 ;
        RECT  3.125 -0.115 3.980 0.115 ;
        RECT  3.005 -0.115 3.125 0.235 ;
        RECT  2.680 -0.115 3.005 0.115 ;
        RECT  2.610 -0.115 2.680 0.405 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.105 1.145 5.180 1.375 ;
        RECT  5.035 0.675 5.105 1.375 ;
        RECT  4.680 1.145 5.035 1.375 ;
        RECT  4.560 1.025 4.680 1.375 ;
        RECT  4.240 1.145 4.560 1.375 ;
        RECT  4.170 1.025 4.240 1.375 ;
        RECT  4.040 1.145 4.170 1.375 ;
        RECT  3.970 1.025 4.040 1.375 ;
        RECT  3.225 1.145 3.970 1.375 ;
        RECT  3.105 0.925 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.705 0.520 4.710 0.660 ;
        RECT  4.635 0.520 4.705 0.955 ;
        RECT  4.320 0.885 4.635 0.955 ;
        RECT  4.390 0.355 4.460 0.805 ;
        RECT  3.990 0.355 4.390 0.425 ;
        RECT  4.250 0.705 4.320 0.955 ;
        RECT  4.070 0.500 4.305 0.635 ;
        RECT  3.825 0.705 4.250 0.775 ;
        RECT  3.650 0.855 4.180 0.925 ;
        RECT  3.910 0.355 3.990 0.605 ;
        RECT  3.755 0.325 3.825 0.775 ;
        RECT  3.375 0.995 3.775 1.065 ;
        RECT  3.535 0.785 3.650 0.925 ;
        RECT  3.465 0.345 3.535 0.925 ;
        RECT  3.375 0.195 3.480 0.265 ;
        RECT  3.305 0.195 3.375 1.065 ;
        RECT  3.155 0.315 3.225 0.840 ;
        RECT  2.790 0.315 3.155 0.385 ;
        RECT  2.595 0.770 3.155 0.840 ;
        RECT  2.930 0.485 3.055 0.615 ;
        RECT  2.540 0.485 2.930 0.555 ;
        RECT  2.215 0.920 2.705 0.990 ;
        RECT  2.515 0.625 2.595 0.840 ;
        RECT  2.470 0.195 2.540 0.555 ;
        RECT  2.065 0.195 2.470 0.265 ;
        RECT  2.285 0.485 2.390 0.820 ;
        RECT  2.215 0.335 2.330 0.405 ;
        RECT  2.135 0.335 2.215 0.990 ;
        RECT  2.020 0.195 2.065 0.435 ;
        RECT  1.975 0.195 2.020 0.960 ;
        RECT  1.950 0.335 1.975 0.960 ;
        RECT  0.640 0.195 1.895 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.150 0.525 4.220 0.595 ;
        RECT  2.305 0.525 2.375 0.595 ;
    END
END SDFCNQND2BWP40

MACRO SDFCNQND4BWP40
    CLASS CORE ;
    FOREIGN SDFCNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.370 0.745 5.480 1.000 ;
        RECT  5.385 0.205 5.470 0.485 ;
        RECT  5.355 0.355 5.385 0.485 ;
        RECT  5.355 0.745 5.370 0.830 ;
        RECT  5.145 0.355 5.355 0.830 ;
        RECT  5.090 0.355 5.145 0.470 ;
        RECT  5.090 0.710 5.145 0.830 ;
        RECT  5.005 0.205 5.090 0.470 ;
        RECT  5.005 0.710 5.090 1.000 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.245 0.525 4.785 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.115 5.740 0.115 ;
        RECT  5.590 -0.115 5.660 0.475 ;
        RECT  5.265 -0.115 5.590 0.115 ;
        RECT  5.195 -0.115 5.265 0.275 ;
        RECT  4.900 -0.115 5.195 0.115 ;
        RECT  4.780 -0.115 4.900 0.145 ;
        RECT  3.980 -0.115 4.780 0.115 ;
        RECT  3.910 -0.115 3.980 0.285 ;
        RECT  3.125 -0.115 3.910 0.115 ;
        RECT  3.005 -0.115 3.125 0.235 ;
        RECT  2.680 -0.115 3.005 0.115 ;
        RECT  2.610 -0.115 2.680 0.420 ;
        RECT  1.500 -0.115 2.610 0.115 ;
        RECT  1.380 -0.115 1.500 0.125 ;
        RECT  1.190 -0.115 1.380 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.145 5.740 1.375 ;
        RECT  5.590 0.705 5.660 1.375 ;
        RECT  5.265 1.145 5.590 1.375 ;
        RECT  5.195 0.915 5.265 1.375 ;
        RECT  4.885 1.145 5.195 1.375 ;
        RECT  4.815 0.835 4.885 1.375 ;
        RECT  4.505 1.145 4.815 1.375 ;
        RECT  4.415 1.095 4.505 1.375 ;
        RECT  4.100 1.145 4.415 1.375 ;
        RECT  3.970 1.035 4.100 1.375 ;
        RECT  3.225 1.145 3.970 1.375 ;
        RECT  3.105 1.040 3.225 1.375 ;
        RECT  2.515 1.145 3.105 1.375 ;
        RECT  2.405 1.065 2.515 1.375 ;
        RECT  1.460 1.145 2.405 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.745 5.480 1.000 ;
        RECT  5.425 0.205 5.470 0.485 ;
        RECT  5.005 0.205 5.075 0.470 ;
        RECT  5.005 0.710 5.075 1.000 ;
        RECT  4.925 0.545 5.045 0.615 ;
        RECT  4.855 0.220 4.925 0.615 ;
        RECT  4.210 0.220 4.855 0.295 ;
        RECT  4.625 0.495 4.780 0.765 ;
        RECT  4.545 0.925 4.710 1.000 ;
        RECT  4.475 0.375 4.545 1.000 ;
        RECT  4.400 0.375 4.475 0.445 ;
        RECT  4.020 0.545 4.475 0.615 ;
        RECT  4.300 0.855 4.375 1.005 ;
        RECT  3.930 0.855 4.300 0.925 ;
        RECT  3.860 0.705 4.295 0.775 ;
        RECT  4.140 0.220 4.210 0.425 ;
        RECT  3.860 0.355 4.140 0.425 ;
        RECT  3.860 0.845 3.930 0.925 ;
        RECT  3.790 0.355 3.860 0.775 ;
        RECT  3.540 0.845 3.860 0.915 ;
        RECT  3.670 0.355 3.790 0.425 ;
        RECT  3.655 0.995 3.780 1.075 ;
        RECT  3.375 0.995 3.655 1.065 ;
        RECT  3.470 0.335 3.540 0.915 ;
        RECT  3.375 0.195 3.435 0.265 ;
        RECT  3.305 0.195 3.375 1.065 ;
        RECT  3.145 0.315 3.215 0.840 ;
        RECT  2.790 0.315 3.145 0.385 ;
        RECT  2.600 0.770 3.145 0.840 ;
        RECT  2.945 0.495 3.060 0.625 ;
        RECT  2.530 0.495 2.945 0.565 ;
        RECT  2.205 0.920 2.705 0.990 ;
        RECT  2.525 0.635 2.600 0.840 ;
        RECT  2.460 0.195 2.530 0.565 ;
        RECT  2.065 0.195 2.460 0.265 ;
        RECT  2.285 0.495 2.390 0.750 ;
        RECT  2.205 0.345 2.305 0.415 ;
        RECT  2.135 0.345 2.205 0.990 ;
        RECT  2.020 0.195 2.065 0.435 ;
        RECT  1.975 0.195 2.020 0.960 ;
        RECT  1.950 0.335 1.975 0.960 ;
        RECT  0.640 0.195 1.895 0.265 ;
        RECT  1.680 0.875 1.860 0.945 ;
        RECT  1.705 0.350 1.775 0.795 ;
        RECT  1.590 0.350 1.705 0.435 ;
        RECT  1.560 0.725 1.705 0.795 ;
        RECT  1.610 0.875 1.680 1.055 ;
        RECT  0.715 0.985 1.610 1.055 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.820 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.665 0.525 4.735 0.595 ;
        RECT  2.305 0.525 2.375 0.595 ;
    END
END SDFCNQND4BWP40

MACRO SDFCSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.215 5.565 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.390 -0.115 5.600 0.115 ;
        RECT  5.255 -0.115 5.390 0.350 ;
        RECT  4.360 -0.115 5.255 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.200 -0.115 3.455 0.115 ;
        RECT  1.080 -0.115 1.200 0.125 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.380 1.145 5.600 1.375 ;
        RECT  5.260 0.950 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  4.955 0.930 5.075 1.000 ;
        RECT  4.785 0.510 5.005 0.630 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.875 0.710 4.955 1.000 ;
        RECT  3.920 0.930 4.875 1.000 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.790 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.365 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.710 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  1.720 0.575 1.800 0.645 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.350 1.720 0.790 ;
        RECT  1.590 0.350 1.650 0.420 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFCSNQD0BWP40

MACRO SDFCSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.032200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.370 -0.115 5.600 0.115 ;
        RECT  5.275 -0.115 5.370 0.310 ;
        RECT  4.360 -0.115 5.275 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.200 -0.115 3.455 0.115 ;
        RECT  1.080 -0.115 1.200 0.125 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.380 1.145 5.600 1.375 ;
        RECT  5.260 0.865 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  3.920 0.930 5.075 1.000 ;
        RECT  4.785 0.460 5.005 0.580 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.710 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  1.720 0.575 1.800 0.645 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.350 1.720 0.790 ;
        RECT  1.590 0.350 1.650 0.420 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFCSNQD1BWP40

MACRO SDFCSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.032200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 -0.115 5.880 0.115 ;
        RECT  5.740 -0.115 5.810 0.485 ;
        RECT  5.390 -0.115 5.740 0.115 ;
        RECT  5.255 -0.115 5.390 0.310 ;
        RECT  4.360 -0.115 5.255 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.200 -0.115 3.455 0.115 ;
        RECT  1.080 -0.115 1.200 0.125 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 1.145 5.880 1.375 ;
        RECT  5.740 0.690 5.810 1.375 ;
        RECT  5.380 1.145 5.740 1.375 ;
        RECT  5.260 0.955 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  3.920 0.930 5.075 1.000 ;
        RECT  4.785 0.460 5.005 0.580 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.715 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  1.720 0.575 1.800 0.645 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.350 1.720 0.790 ;
        RECT  1.590 0.350 1.650 0.420 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFCSNQD2BWP40

MACRO SDFCSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.450 5.870 0.765 ;
        RECT  5.765 0.525 5.775 0.635 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.405 0.195 6.500 0.485 ;
        RECT  6.405 0.710 6.500 0.995 ;
        RECT  6.335 0.355 6.405 0.485 ;
        RECT  6.335 0.710 6.405 0.830 ;
        RECT  6.125 0.355 6.335 0.830 ;
        RECT  6.100 0.355 6.125 0.485 ;
        RECT  6.100 0.710 6.125 0.830 ;
        RECT  6.025 0.215 6.100 0.485 ;
        RECT  6.025 0.710 6.100 0.995 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.044600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.315 0.355 4.445 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 -0.115 6.720 0.115 ;
        RECT  6.595 -0.115 6.665 0.440 ;
        RECT  6.290 -0.115 6.595 0.115 ;
        RECT  6.205 -0.115 6.290 0.265 ;
        RECT  5.920 -0.115 6.205 0.115 ;
        RECT  5.830 -0.115 5.920 0.310 ;
        RECT  5.170 -0.115 5.830 0.115 ;
        RECT  5.050 -0.115 5.170 0.140 ;
        RECT  4.370 -0.115 5.050 0.115 ;
        RECT  4.235 -0.115 4.370 0.130 ;
        RECT  3.525 -0.115 4.235 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.200 -0.115 3.455 0.115 ;
        RECT  1.080 -0.115 1.200 0.125 ;
        RECT  0.340 -0.115 1.080 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.145 6.720 1.375 ;
        RECT  6.595 0.680 6.665 1.375 ;
        RECT  6.310 1.145 6.595 1.375 ;
        RECT  6.190 0.960 6.310 1.375 ;
        RECT  5.910 1.145 6.190 1.375 ;
        RECT  5.835 0.955 5.910 1.375 ;
        RECT  5.000 1.145 5.835 1.375 ;
        RECT  4.880 1.070 5.000 1.375 ;
        RECT  4.370 1.145 4.880 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.405 0.195 6.500 0.485 ;
        RECT  6.405 0.710 6.500 0.995 ;
        RECT  6.025 0.215 6.055 0.485 ;
        RECT  6.025 0.710 6.055 0.995 ;
        RECT  5.625 0.210 5.695 1.000 ;
        RECT  5.045 0.930 5.625 1.000 ;
        RECT  5.515 0.620 5.555 0.740 ;
        RECT  5.445 0.210 5.515 0.860 ;
        RECT  4.765 0.210 5.445 0.280 ;
        RECT  5.330 0.790 5.445 0.860 ;
        RECT  4.845 0.350 5.350 0.420 ;
        RECT  4.965 0.605 5.045 1.000 ;
        RECT  3.920 0.930 4.965 1.000 ;
        RECT  4.695 0.210 4.765 0.860 ;
        RECT  4.690 0.335 4.695 0.860 ;
        RECT  4.675 0.335 4.690 0.445 ;
        RECT  4.205 0.790 4.690 0.860 ;
        RECT  4.585 0.580 4.620 0.700 ;
        RECT  4.515 0.200 4.585 0.700 ;
        RECT  3.980 0.200 4.515 0.270 ;
        RECT  4.135 0.445 4.205 0.860 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.935 0.195 3.980 0.270 ;
        RECT  3.685 0.195 3.935 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.715 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  0.640 0.195 1.920 0.265 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  1.720 0.575 1.800 0.645 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.350 1.720 0.790 ;
        RECT  1.590 0.350 1.650 0.420 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFCSNQD4BWP40

MACRO SDFKCNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFKCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.495 1.035 0.565 ;
        RECT  0.870 0.215 0.955 0.565 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.355 1.505 0.640 ;
        RECT  1.310 0.510 1.385 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.195 4.725 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.011800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 -0.115 4.760 0.115 ;
        RECT  4.445 -0.115 4.515 0.305 ;
        RECT  4.145 -0.115 4.445 0.115 ;
        RECT  4.075 -0.115 4.145 0.315 ;
        RECT  3.385 -0.115 4.075 0.115 ;
        RECT  3.315 -0.115 3.385 0.420 ;
        RECT  3.010 -0.115 3.315 0.115 ;
        RECT  2.890 -0.115 3.010 0.210 ;
        RECT  2.030 -0.115 2.890 0.115 ;
        RECT  1.910 -0.115 2.030 0.125 ;
        RECT  1.490 -0.115 1.910 0.115 ;
        RECT  1.370 -0.115 1.490 0.265 ;
        RECT  1.095 -0.115 1.370 0.115 ;
        RECT  1.025 -0.115 1.095 0.415 ;
        RECT  0.125 -0.115 1.025 0.115 ;
        RECT  0.055 -0.115 0.125 0.305 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 1.145 4.760 1.375 ;
        RECT  4.445 0.955 4.515 1.375 ;
        RECT  4.150 1.145 4.445 1.375 ;
        RECT  4.080 0.950 4.150 1.375 ;
        RECT  3.385 1.145 4.080 1.375 ;
        RECT  3.315 0.785 3.385 1.375 ;
        RECT  3.005 1.145 3.315 1.375 ;
        RECT  2.895 0.890 3.005 1.375 ;
        RECT  2.050 1.145 2.895 1.375 ;
        RECT  1.930 1.135 2.050 1.375 ;
        RECT  1.500 1.145 1.930 1.375 ;
        RECT  1.380 1.110 1.500 1.375 ;
        RECT  1.140 1.145 1.380 1.375 ;
        RECT  1.020 1.050 1.140 1.375 ;
        RECT  0.340 1.145 1.020 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.395 4.515 0.820 ;
        RECT  4.335 0.395 4.445 0.465 ;
        RECT  4.335 0.750 4.445 0.820 ;
        RECT  4.010 0.545 4.340 0.615 ;
        RECT  4.265 0.195 4.335 0.465 ;
        RECT  4.265 0.750 4.335 1.070 ;
        RECT  3.970 0.395 4.265 0.465 ;
        RECT  3.940 0.545 4.010 1.045 ;
        RECT  3.880 0.545 3.940 0.615 ;
        RECT  3.660 0.975 3.940 1.045 ;
        RECT  3.800 0.220 3.880 0.615 ;
        RECT  3.800 0.770 3.870 0.890 ;
        RECT  3.660 0.220 3.800 0.290 ;
        RECT  3.690 0.770 3.800 0.840 ;
        RECT  3.620 0.440 3.690 0.840 ;
        RECT  3.120 0.300 3.190 0.980 ;
        RECT  2.905 0.745 3.120 0.815 ;
        RECT  2.980 0.280 3.050 0.640 ;
        RECT  2.605 0.280 2.980 0.350 ;
        RECT  2.835 0.695 2.905 0.815 ;
        RECT  2.745 0.420 2.820 0.490 ;
        RECT  2.745 0.885 2.815 0.955 ;
        RECT  2.675 0.420 2.745 0.955 ;
        RECT  2.535 0.205 2.605 0.925 ;
        RECT  1.655 0.205 2.445 0.275 ;
        RECT  2.345 0.865 2.415 1.065 ;
        RECT  1.580 0.995 2.345 1.065 ;
        RECT  2.235 0.355 2.305 0.795 ;
        RECT  2.135 0.355 2.235 0.425 ;
        RECT  2.135 0.725 2.235 0.795 ;
        RECT  2.065 0.545 2.155 0.615 ;
        RECT  1.995 0.355 2.065 0.830 ;
        RECT  1.740 0.355 1.995 0.425 ;
        RECT  1.750 0.750 1.995 0.830 ;
        RECT  1.585 0.205 1.655 0.330 ;
        RECT  1.575 0.510 1.645 0.920 ;
        RECT  0.695 0.850 1.575 0.920 ;
        RECT  1.240 0.710 1.330 0.780 ;
        RECT  1.240 0.190 1.275 0.310 ;
        RECT  1.170 0.190 1.240 0.780 ;
        RECT  0.855 0.710 1.170 0.780 ;
        RECT  0.775 0.635 0.855 0.780 ;
        RECT  0.625 0.200 0.695 0.920 ;
        RECT  0.505 0.205 0.545 0.915 ;
        RECT  0.475 0.205 0.505 1.065 ;
        RECT  0.380 0.205 0.475 0.275 ;
        RECT  0.435 0.845 0.475 1.065 ;
        RECT  0.125 0.845 0.435 0.915 ;
        RECT  0.055 0.845 0.125 1.005 ;
    END
END SDFKCNQD0BWP40

MACRO SDFKCNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFKCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.495 1.060 0.565 ;
        RECT  0.870 0.215 0.955 0.565 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.355 1.505 0.625 ;
        RECT  1.305 0.545 1.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.635 0.185 4.725 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 -0.115 4.760 0.115 ;
        RECT  4.445 -0.115 4.515 0.305 ;
        RECT  4.145 -0.115 4.445 0.115 ;
        RECT  4.075 -0.115 4.145 0.315 ;
        RECT  3.385 -0.115 4.075 0.115 ;
        RECT  3.315 -0.115 3.385 0.445 ;
        RECT  3.040 -0.115 3.315 0.115 ;
        RECT  2.920 -0.115 3.040 0.210 ;
        RECT  2.060 -0.115 2.920 0.115 ;
        RECT  1.940 -0.115 2.060 0.130 ;
        RECT  1.490 -0.115 1.940 0.115 ;
        RECT  1.375 -0.115 1.490 0.265 ;
        RECT  1.095 -0.115 1.375 0.115 ;
        RECT  1.025 -0.115 1.095 0.415 ;
        RECT  0.125 -0.115 1.025 0.115 ;
        RECT  0.055 -0.115 0.125 0.400 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 1.145 4.760 1.375 ;
        RECT  4.445 0.835 4.515 1.375 ;
        RECT  4.150 1.145 4.445 1.375 ;
        RECT  4.080 0.950 4.150 1.375 ;
        RECT  3.385 1.145 4.080 1.375 ;
        RECT  3.315 0.700 3.385 1.375 ;
        RECT  3.015 1.145 3.315 1.375 ;
        RECT  2.945 0.865 3.015 1.375 ;
        RECT  2.040 1.145 2.945 1.375 ;
        RECT  1.920 1.135 2.040 1.375 ;
        RECT  1.500 1.145 1.920 1.375 ;
        RECT  1.380 1.110 1.500 1.375 ;
        RECT  1.115 1.145 1.380 1.375 ;
        RECT  1.045 1.020 1.115 1.375 ;
        RECT  0.315 1.145 1.045 1.375 ;
        RECT  0.245 0.870 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.395 4.515 0.755 ;
        RECT  4.335 0.395 4.445 0.465 ;
        RECT  4.335 0.685 4.445 0.755 ;
        RECT  4.010 0.545 4.340 0.615 ;
        RECT  4.265 0.195 4.335 0.465 ;
        RECT  4.265 0.685 4.335 1.070 ;
        RECT  3.970 0.395 4.265 0.465 ;
        RECT  3.940 0.545 4.010 1.045 ;
        RECT  3.880 0.545 3.940 0.615 ;
        RECT  3.660 0.975 3.940 1.045 ;
        RECT  3.800 0.220 3.880 0.615 ;
        RECT  3.800 0.770 3.870 0.890 ;
        RECT  3.660 0.220 3.800 0.290 ;
        RECT  3.690 0.770 3.800 0.840 ;
        RECT  3.620 0.440 3.690 0.840 ;
        RECT  3.150 0.300 3.220 0.980 ;
        RECT  3.135 0.300 3.150 0.415 ;
        RECT  3.135 0.720 3.150 0.980 ;
        RECT  2.945 0.720 3.135 0.790 ;
        RECT  3.065 0.470 3.080 0.590 ;
        RECT  2.995 0.280 3.065 0.590 ;
        RECT  2.605 0.280 2.995 0.350 ;
        RECT  2.875 0.670 2.945 0.790 ;
        RECT  2.785 0.420 2.835 0.490 ;
        RECT  2.785 0.885 2.830 0.955 ;
        RECT  2.715 0.420 2.785 0.955 ;
        RECT  2.535 0.280 2.605 0.965 ;
        RECT  1.655 0.205 2.435 0.275 ;
        RECT  2.345 0.865 2.415 1.065 ;
        RECT  2.285 0.355 2.355 0.795 ;
        RECT  1.580 0.995 2.345 1.065 ;
        RECT  2.135 0.355 2.285 0.425 ;
        RECT  2.135 0.725 2.285 0.795 ;
        RECT  2.065 0.545 2.155 0.615 ;
        RECT  1.995 0.355 2.065 0.850 ;
        RECT  1.740 0.355 1.995 0.425 ;
        RECT  1.765 0.780 1.995 0.850 ;
        RECT  1.585 0.205 1.655 0.410 ;
        RECT  1.575 0.510 1.645 0.920 ;
        RECT  0.695 0.850 1.575 0.920 ;
        RECT  1.235 0.710 1.330 0.780 ;
        RECT  1.235 0.190 1.275 0.310 ;
        RECT  1.165 0.190 1.235 0.780 ;
        RECT  0.845 0.710 1.165 0.780 ;
        RECT  0.775 0.635 0.845 0.780 ;
        RECT  0.625 0.200 0.695 1.075 ;
        RECT  0.505 0.205 0.545 0.790 ;
        RECT  0.475 0.205 0.505 0.990 ;
        RECT  0.380 0.205 0.475 0.275 ;
        RECT  0.435 0.720 0.475 0.990 ;
        RECT  0.125 0.720 0.435 0.790 ;
        RECT  0.055 0.720 0.125 1.075 ;
    END
END SDFKCNQD1BWP40

MACRO SDFKCNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFKCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.495 1.060 0.565 ;
        RECT  0.870 0.215 0.955 0.565 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.355 1.505 0.625 ;
        RECT  1.305 0.545 1.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.645 0.185 4.735 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 -0.115 5.040 0.115 ;
        RECT  4.885 -0.115 4.970 0.470 ;
        RECT  4.515 -0.115 4.885 0.115 ;
        RECT  4.445 -0.115 4.515 0.305 ;
        RECT  4.145 -0.115 4.445 0.115 ;
        RECT  4.075 -0.115 4.145 0.315 ;
        RECT  3.385 -0.115 4.075 0.115 ;
        RECT  3.315 -0.115 3.385 0.445 ;
        RECT  3.040 -0.115 3.315 0.115 ;
        RECT  2.920 -0.115 3.040 0.210 ;
        RECT  2.060 -0.115 2.920 0.115 ;
        RECT  1.940 -0.115 2.060 0.130 ;
        RECT  1.490 -0.115 1.940 0.115 ;
        RECT  1.375 -0.115 1.490 0.265 ;
        RECT  1.095 -0.115 1.375 0.115 ;
        RECT  1.025 -0.115 1.095 0.415 ;
        RECT  0.125 -0.115 1.025 0.115 ;
        RECT  0.055 -0.115 0.125 0.400 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.970 1.145 5.040 1.375 ;
        RECT  4.885 0.670 4.970 1.375 ;
        RECT  4.515 1.145 4.885 1.375 ;
        RECT  4.445 0.835 4.515 1.375 ;
        RECT  4.150 1.145 4.445 1.375 ;
        RECT  4.080 0.950 4.150 1.375 ;
        RECT  3.385 1.145 4.080 1.375 ;
        RECT  3.315 0.700 3.385 1.375 ;
        RECT  3.015 1.145 3.315 1.375 ;
        RECT  2.945 0.865 3.015 1.375 ;
        RECT  2.040 1.145 2.945 1.375 ;
        RECT  1.920 1.135 2.040 1.375 ;
        RECT  1.500 1.145 1.920 1.375 ;
        RECT  1.380 1.110 1.500 1.375 ;
        RECT  1.115 1.145 1.380 1.375 ;
        RECT  1.045 1.020 1.115 1.375 ;
        RECT  0.315 1.145 1.045 1.375 ;
        RECT  0.245 0.870 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.445 0.395 4.515 0.755 ;
        RECT  4.335 0.395 4.445 0.465 ;
        RECT  4.335 0.685 4.445 0.755 ;
        RECT  4.010 0.545 4.340 0.615 ;
        RECT  4.265 0.195 4.335 0.465 ;
        RECT  4.265 0.685 4.335 1.070 ;
        RECT  3.970 0.395 4.265 0.465 ;
        RECT  3.940 0.545 4.010 1.045 ;
        RECT  3.880 0.545 3.940 0.615 ;
        RECT  3.660 0.975 3.940 1.045 ;
        RECT  3.800 0.220 3.880 0.615 ;
        RECT  3.800 0.770 3.870 0.890 ;
        RECT  3.660 0.220 3.800 0.290 ;
        RECT  3.690 0.770 3.800 0.840 ;
        RECT  3.620 0.440 3.690 0.840 ;
        RECT  3.150 0.300 3.220 0.980 ;
        RECT  3.135 0.300 3.150 0.415 ;
        RECT  3.135 0.720 3.150 0.980 ;
        RECT  2.945 0.720 3.135 0.790 ;
        RECT  3.065 0.470 3.080 0.590 ;
        RECT  2.995 0.280 3.065 0.590 ;
        RECT  2.605 0.280 2.995 0.350 ;
        RECT  2.875 0.670 2.945 0.790 ;
        RECT  2.785 0.420 2.835 0.490 ;
        RECT  2.785 0.885 2.830 0.955 ;
        RECT  2.715 0.420 2.785 0.955 ;
        RECT  2.535 0.280 2.605 0.965 ;
        RECT  1.655 0.205 2.435 0.275 ;
        RECT  2.345 0.865 2.415 1.065 ;
        RECT  2.285 0.355 2.355 0.795 ;
        RECT  1.580 0.995 2.345 1.065 ;
        RECT  2.135 0.355 2.285 0.425 ;
        RECT  2.135 0.725 2.285 0.795 ;
        RECT  2.065 0.545 2.155 0.615 ;
        RECT  1.995 0.355 2.065 0.850 ;
        RECT  1.740 0.355 1.995 0.425 ;
        RECT  1.765 0.780 1.995 0.850 ;
        RECT  1.585 0.205 1.655 0.410 ;
        RECT  1.575 0.510 1.645 0.920 ;
        RECT  0.695 0.850 1.575 0.920 ;
        RECT  1.235 0.710 1.330 0.780 ;
        RECT  1.235 0.190 1.275 0.310 ;
        RECT  1.165 0.190 1.235 0.780 ;
        RECT  0.845 0.710 1.165 0.780 ;
        RECT  0.775 0.635 0.845 0.780 ;
        RECT  0.625 0.200 0.695 1.075 ;
        RECT  0.505 0.205 0.545 0.790 ;
        RECT  0.475 0.205 0.505 0.990 ;
        RECT  0.380 0.205 0.475 0.275 ;
        RECT  0.435 0.720 0.475 0.990 ;
        RECT  0.125 0.720 0.435 0.790 ;
        RECT  0.055 0.720 0.125 1.075 ;
    END
END SDFKCNQD2BWP40

MACRO SDFKCNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFKCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.495 1.060 0.565 ;
        RECT  0.870 0.215 0.955 0.565 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.355 1.505 0.625 ;
        RECT  1.305 0.545 1.385 0.625 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.265 0.205 5.355 0.465 ;
        RECT  5.265 0.685 5.355 1.075 ;
        RECT  5.215 0.380 5.265 0.465 ;
        RECT  5.215 0.685 5.265 0.770 ;
        RECT  5.005 0.380 5.215 0.770 ;
        RECT  4.995 0.380 5.005 0.465 ;
        RECT  4.995 0.685 5.005 0.770 ;
        RECT  4.905 0.205 4.995 0.465 ;
        RECT  4.905 0.685 4.995 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.245 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.495 1.925 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 0.355 0.405 0.640 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 -0.115 5.600 0.115 ;
        RECT  5.475 -0.115 5.545 0.445 ;
        RECT  5.165 -0.115 5.475 0.115 ;
        RECT  5.095 -0.115 5.165 0.255 ;
        RECT  4.785 -0.115 5.095 0.115 ;
        RECT  4.715 -0.115 4.785 0.445 ;
        RECT  4.405 -0.115 4.715 0.115 ;
        RECT  4.335 -0.115 4.405 0.305 ;
        RECT  3.585 -0.115 4.335 0.115 ;
        RECT  3.515 -0.115 3.585 0.380 ;
        RECT  3.040 -0.115 3.515 0.115 ;
        RECT  2.920 -0.115 3.040 0.210 ;
        RECT  2.060 -0.115 2.920 0.115 ;
        RECT  1.940 -0.115 2.060 0.130 ;
        RECT  1.490 -0.115 1.940 0.115 ;
        RECT  1.375 -0.115 1.490 0.265 ;
        RECT  1.095 -0.115 1.375 0.115 ;
        RECT  1.025 -0.115 1.095 0.415 ;
        RECT  0.125 -0.115 1.025 0.115 ;
        RECT  0.055 -0.115 0.125 0.400 ;
        RECT  0.000 -0.115 0.055 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 1.145 5.600 1.375 ;
        RECT  5.475 0.715 5.545 1.375 ;
        RECT  5.165 1.145 5.475 1.375 ;
        RECT  5.095 0.885 5.165 1.375 ;
        RECT  4.785 1.145 5.095 1.375 ;
        RECT  4.715 0.715 4.785 1.375 ;
        RECT  4.410 1.145 4.715 1.375 ;
        RECT  4.340 0.950 4.410 1.375 ;
        RECT  3.585 1.145 4.340 1.375 ;
        RECT  3.515 0.740 3.585 1.375 ;
        RECT  3.015 1.145 3.515 1.375 ;
        RECT  2.945 0.865 3.015 1.375 ;
        RECT  2.040 1.145 2.945 1.375 ;
        RECT  1.920 1.135 2.040 1.375 ;
        RECT  1.500 1.145 1.920 1.375 ;
        RECT  1.380 1.110 1.500 1.375 ;
        RECT  1.115 1.145 1.380 1.375 ;
        RECT  1.045 1.020 1.115 1.375 ;
        RECT  0.315 1.145 1.045 1.375 ;
        RECT  0.245 0.870 0.315 1.375 ;
        RECT  0.000 1.145 0.245 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.205 5.355 0.465 ;
        RECT  5.285 0.685 5.355 1.075 ;
        RECT  4.905 0.205 4.935 0.465 ;
        RECT  4.905 0.685 4.935 1.075 ;
        RECT  4.595 0.395 4.645 0.785 ;
        RECT  4.575 0.185 4.595 1.070 ;
        RECT  4.525 0.185 4.575 0.465 ;
        RECT  4.525 0.715 4.575 1.070 ;
        RECT  4.220 0.395 4.525 0.465 ;
        RECT  4.270 0.545 4.505 0.615 ;
        RECT  4.200 0.545 4.270 1.050 ;
        RECT  4.150 0.545 4.200 0.615 ;
        RECT  3.930 0.980 4.200 1.050 ;
        RECT  4.070 0.240 4.150 0.615 ;
        RECT  4.060 0.780 4.130 0.900 ;
        RECT  3.930 0.240 4.070 0.310 ;
        RECT  3.960 0.780 4.060 0.850 ;
        RECT  3.890 0.440 3.960 0.850 ;
        RECT  3.715 0.315 3.785 0.520 ;
        RECT  3.715 0.600 3.785 0.955 ;
        RECT  3.385 0.450 3.715 0.520 ;
        RECT  3.385 0.600 3.715 0.670 ;
        RECT  3.315 0.315 3.385 0.520 ;
        RECT  3.315 0.600 3.385 0.955 ;
        RECT  3.150 0.300 3.220 0.980 ;
        RECT  3.135 0.300 3.150 0.415 ;
        RECT  3.135 0.720 3.150 0.980 ;
        RECT  2.945 0.720 3.135 0.790 ;
        RECT  3.065 0.470 3.080 0.590 ;
        RECT  2.995 0.280 3.065 0.590 ;
        RECT  2.605 0.280 2.995 0.350 ;
        RECT  2.875 0.670 2.945 0.790 ;
        RECT  2.785 0.420 2.835 0.490 ;
        RECT  2.785 0.885 2.830 0.955 ;
        RECT  2.715 0.420 2.785 0.955 ;
        RECT  2.535 0.280 2.605 0.965 ;
        RECT  1.655 0.205 2.435 0.275 ;
        RECT  2.345 0.865 2.415 1.065 ;
        RECT  2.285 0.355 2.355 0.795 ;
        RECT  1.580 0.995 2.345 1.065 ;
        RECT  2.135 0.355 2.285 0.425 ;
        RECT  2.135 0.725 2.285 0.795 ;
        RECT  2.065 0.545 2.155 0.615 ;
        RECT  1.995 0.355 2.065 0.850 ;
        RECT  1.740 0.355 1.995 0.425 ;
        RECT  1.765 0.780 1.995 0.850 ;
        RECT  1.585 0.205 1.655 0.410 ;
        RECT  1.575 0.510 1.645 0.920 ;
        RECT  0.695 0.850 1.575 0.920 ;
        RECT  1.235 0.710 1.330 0.780 ;
        RECT  1.235 0.190 1.275 0.310 ;
        RECT  1.165 0.190 1.235 0.780 ;
        RECT  0.845 0.710 1.165 0.780 ;
        RECT  0.775 0.635 0.845 0.780 ;
        RECT  0.625 0.200 0.695 1.075 ;
        RECT  0.505 0.205 0.545 0.790 ;
        RECT  0.475 0.205 0.505 0.990 ;
        RECT  0.380 0.205 0.475 0.275 ;
        RECT  0.435 0.720 0.475 0.990 ;
        RECT  0.125 0.720 0.435 0.790 ;
        RECT  0.055 0.720 0.125 1.075 ;
    END
END SDFKCNQD4BWP40

MACRO SDFKCSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFKCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.765 0.230 0.835 ;
        RECT  0.035 0.495 0.125 0.835 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.500 1.635 0.570 ;
        RECT  1.425 0.215 1.505 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.355 2.065 0.640 ;
        RECT  1.880 0.520 1.930 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.195 0.195 5.285 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.765 0.595 0.835 ;
        RECT  0.455 0.765 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.485 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.011800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.875 ;
        RECT  0.435 0.475 0.875 0.545 ;
        RECT  0.735 0.805 0.875 0.875 ;
        RECT  0.355 0.410 0.435 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.075 -0.115 5.320 0.115 ;
        RECT  5.005 -0.115 5.075 0.305 ;
        RECT  4.705 -0.115 5.005 0.115 ;
        RECT  4.635 -0.115 4.705 0.315 ;
        RECT  3.945 -0.115 4.635 0.115 ;
        RECT  3.875 -0.115 3.945 0.420 ;
        RECT  3.570 -0.115 3.875 0.115 ;
        RECT  3.450 -0.115 3.570 0.210 ;
        RECT  2.590 -0.115 3.450 0.115 ;
        RECT  2.470 -0.115 2.590 0.135 ;
        RECT  2.050 -0.115 2.470 0.115 ;
        RECT  1.930 -0.115 2.050 0.270 ;
        RECT  1.655 -0.115 1.930 0.115 ;
        RECT  1.585 -0.115 1.655 0.420 ;
        RECT  0.315 -0.115 1.585 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.075 1.145 5.320 1.375 ;
        RECT  5.005 0.955 5.075 1.375 ;
        RECT  4.710 1.145 5.005 1.375 ;
        RECT  4.640 0.950 4.710 1.375 ;
        RECT  3.945 1.145 4.640 1.375 ;
        RECT  3.875 0.785 3.945 1.375 ;
        RECT  3.565 1.145 3.875 1.375 ;
        RECT  3.455 0.890 3.565 1.375 ;
        RECT  2.610 1.145 3.455 1.375 ;
        RECT  2.490 1.130 2.610 1.375 ;
        RECT  2.035 1.145 2.490 1.375 ;
        RECT  1.965 1.025 2.035 1.375 ;
        RECT  1.675 1.145 1.965 1.375 ;
        RECT  1.605 1.025 1.675 1.375 ;
        RECT  0.930 1.145 1.605 1.375 ;
        RECT  0.810 1.110 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.005 0.395 5.075 0.820 ;
        RECT  4.895 0.395 5.005 0.465 ;
        RECT  4.895 0.750 5.005 0.820 ;
        RECT  4.570 0.545 4.900 0.615 ;
        RECT  4.825 0.195 4.895 0.465 ;
        RECT  4.825 0.750 4.895 1.070 ;
        RECT  4.530 0.395 4.825 0.465 ;
        RECT  4.500 0.545 4.570 1.045 ;
        RECT  4.440 0.545 4.500 0.615 ;
        RECT  4.220 0.975 4.500 1.045 ;
        RECT  4.360 0.220 4.440 0.615 ;
        RECT  4.360 0.770 4.430 0.890 ;
        RECT  4.220 0.220 4.360 0.290 ;
        RECT  4.250 0.770 4.360 0.840 ;
        RECT  4.180 0.440 4.250 0.840 ;
        RECT  3.680 0.300 3.750 0.980 ;
        RECT  3.465 0.745 3.680 0.815 ;
        RECT  3.540 0.280 3.610 0.640 ;
        RECT  3.165 0.280 3.540 0.350 ;
        RECT  3.395 0.695 3.465 0.815 ;
        RECT  3.305 0.420 3.380 0.490 ;
        RECT  3.305 0.885 3.375 0.955 ;
        RECT  3.235 0.420 3.305 0.955 ;
        RECT  3.095 0.205 3.165 0.925 ;
        RECT  2.215 0.205 2.980 0.275 ;
        RECT  2.905 0.865 2.975 1.060 ;
        RECT  2.140 0.990 2.905 1.060 ;
        RECT  2.795 0.345 2.865 0.790 ;
        RECT  2.705 0.345 2.795 0.465 ;
        RECT  2.700 0.710 2.795 0.790 ;
        RECT  2.625 0.545 2.695 0.615 ;
        RECT  2.555 0.355 2.625 0.825 ;
        RECT  2.300 0.355 2.555 0.425 ;
        RECT  2.325 0.755 2.555 0.825 ;
        RECT  2.145 0.205 2.215 0.365 ;
        RECT  2.135 0.510 2.205 0.920 ;
        RECT  1.300 0.850 2.135 0.920 ;
        RECT  1.810 0.710 1.890 0.780 ;
        RECT  1.810 0.190 1.835 0.310 ;
        RECT  1.740 0.190 1.810 0.780 ;
        RECT  1.415 0.710 1.740 0.780 ;
        RECT  1.345 0.640 1.415 0.780 ;
        RECT  1.265 0.850 1.300 0.960 ;
        RECT  1.195 0.195 1.265 0.960 ;
        RECT  1.030 0.235 1.105 1.030 ;
        RECT  1.005 0.235 1.030 0.405 ;
        RECT  0.610 0.960 1.030 1.030 ;
        RECT  0.610 0.335 1.005 0.405 ;
        RECT  0.410 0.195 0.920 0.265 ;
        RECT  0.385 0.625 0.805 0.695 ;
        RECT  0.315 0.625 0.385 0.975 ;
        RECT  0.275 0.625 0.315 0.695 ;
        RECT  0.125 0.905 0.315 0.975 ;
        RECT  0.195 0.355 0.275 0.695 ;
        RECT  0.125 0.355 0.195 0.425 ;
        RECT  0.055 0.195 0.125 0.425 ;
        RECT  0.055 0.905 0.125 1.075 ;
    END
END SDFKCSNQD0BWP40

MACRO SDFKCSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFKCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.765 0.230 0.835 ;
        RECT  0.035 0.495 0.125 0.835 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.500 1.635 0.570 ;
        RECT  1.425 0.215 1.505 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.028400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.355 2.065 0.640 ;
        RECT  1.880 0.520 1.930 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.195 0.195 5.285 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.765 0.595 0.835 ;
        RECT  0.455 0.765 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.485 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.014800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.875 ;
        RECT  0.435 0.475 0.875 0.545 ;
        RECT  0.735 0.805 0.875 0.875 ;
        RECT  0.355 0.410 0.435 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.075 -0.115 5.320 0.115 ;
        RECT  5.005 -0.115 5.075 0.305 ;
        RECT  4.705 -0.115 5.005 0.115 ;
        RECT  4.635 -0.115 4.705 0.310 ;
        RECT  3.945 -0.115 4.635 0.115 ;
        RECT  3.875 -0.115 3.945 0.445 ;
        RECT  3.600 -0.115 3.875 0.115 ;
        RECT  3.480 -0.115 3.600 0.210 ;
        RECT  2.620 -0.115 3.480 0.115 ;
        RECT  2.500 -0.115 2.620 0.130 ;
        RECT  2.050 -0.115 2.500 0.115 ;
        RECT  1.935 -0.115 2.050 0.265 ;
        RECT  1.655 -0.115 1.935 0.115 ;
        RECT  1.585 -0.115 1.655 0.420 ;
        RECT  0.315 -0.115 1.585 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.075 1.145 5.320 1.375 ;
        RECT  5.005 0.835 5.075 1.375 ;
        RECT  4.710 1.145 5.005 1.375 ;
        RECT  4.640 0.950 4.710 1.375 ;
        RECT  3.945 1.145 4.640 1.375 ;
        RECT  3.875 0.700 3.945 1.375 ;
        RECT  3.575 1.145 3.875 1.375 ;
        RECT  3.505 0.865 3.575 1.375 ;
        RECT  2.600 1.145 3.505 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.035 1.145 2.480 1.375 ;
        RECT  1.965 1.025 2.035 1.375 ;
        RECT  1.675 1.145 1.965 1.375 ;
        RECT  1.605 1.025 1.675 1.375 ;
        RECT  0.930 1.145 1.605 1.375 ;
        RECT  0.810 1.110 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.005 0.395 5.075 0.755 ;
        RECT  4.895 0.395 5.005 0.465 ;
        RECT  4.895 0.685 5.005 0.755 ;
        RECT  4.570 0.545 4.900 0.615 ;
        RECT  4.825 0.210 4.895 0.465 ;
        RECT  4.825 0.685 4.895 1.070 ;
        RECT  4.510 0.395 4.825 0.465 ;
        RECT  4.500 0.545 4.570 1.045 ;
        RECT  4.425 0.545 4.500 0.615 ;
        RECT  4.220 0.975 4.500 1.045 ;
        RECT  4.360 0.770 4.430 0.890 ;
        RECT  4.345 0.240 4.425 0.615 ;
        RECT  4.250 0.770 4.360 0.840 ;
        RECT  4.220 0.240 4.345 0.310 ;
        RECT  4.180 0.440 4.250 0.840 ;
        RECT  3.710 0.300 3.780 0.980 ;
        RECT  3.695 0.300 3.710 0.415 ;
        RECT  3.695 0.720 3.710 0.980 ;
        RECT  3.505 0.720 3.695 0.790 ;
        RECT  3.625 0.470 3.640 0.590 ;
        RECT  3.555 0.280 3.625 0.590 ;
        RECT  3.165 0.280 3.555 0.350 ;
        RECT  3.435 0.670 3.505 0.790 ;
        RECT  3.345 0.420 3.395 0.490 ;
        RECT  3.345 0.885 3.390 0.955 ;
        RECT  3.275 0.420 3.345 0.955 ;
        RECT  3.095 0.280 3.165 0.965 ;
        RECT  2.215 0.205 2.995 0.275 ;
        RECT  2.905 0.865 2.975 1.060 ;
        RECT  2.845 0.355 2.915 0.795 ;
        RECT  2.140 0.990 2.905 1.060 ;
        RECT  2.695 0.355 2.845 0.425 ;
        RECT  2.695 0.725 2.845 0.795 ;
        RECT  2.625 0.545 2.715 0.615 ;
        RECT  2.555 0.355 2.625 0.850 ;
        RECT  2.300 0.355 2.555 0.425 ;
        RECT  2.325 0.780 2.555 0.850 ;
        RECT  2.145 0.205 2.215 0.410 ;
        RECT  2.135 0.510 2.205 0.920 ;
        RECT  1.265 0.850 2.135 0.920 ;
        RECT  1.810 0.710 1.890 0.780 ;
        RECT  1.810 0.190 1.835 0.310 ;
        RECT  1.740 0.190 1.810 0.780 ;
        RECT  1.425 0.710 1.740 0.780 ;
        RECT  1.345 0.640 1.425 0.780 ;
        RECT  1.195 0.195 1.265 0.920 ;
        RECT  1.030 0.235 1.105 1.030 ;
        RECT  1.005 0.235 1.030 0.405 ;
        RECT  0.610 0.960 1.030 1.030 ;
        RECT  0.610 0.335 1.005 0.405 ;
        RECT  0.410 0.195 0.920 0.265 ;
        RECT  0.385 0.625 0.805 0.695 ;
        RECT  0.315 0.625 0.385 0.975 ;
        RECT  0.275 0.625 0.315 0.695 ;
        RECT  0.125 0.905 0.315 0.975 ;
        RECT  0.195 0.355 0.275 0.695 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.905 0.125 1.075 ;
    END
END SDFKCSNQD1BWP40

MACRO SDFKCSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFKCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.765 0.230 0.835 ;
        RECT  0.035 0.495 0.125 0.835 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.500 1.635 0.570 ;
        RECT  1.425 0.215 1.505 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.028400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.355 2.065 0.640 ;
        RECT  1.880 0.520 1.930 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.205 0.185 5.295 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.765 0.595 0.835 ;
        RECT  0.455 0.765 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.485 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.014800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.875 ;
        RECT  0.435 0.475 0.875 0.545 ;
        RECT  0.735 0.805 0.875 0.875 ;
        RECT  0.355 0.410 0.435 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.530 -0.115 5.600 0.115 ;
        RECT  5.445 -0.115 5.530 0.470 ;
        RECT  5.075 -0.115 5.445 0.115 ;
        RECT  5.005 -0.115 5.075 0.305 ;
        RECT  4.705 -0.115 5.005 0.115 ;
        RECT  4.635 -0.115 4.705 0.310 ;
        RECT  3.945 -0.115 4.635 0.115 ;
        RECT  3.875 -0.115 3.945 0.445 ;
        RECT  3.600 -0.115 3.875 0.115 ;
        RECT  3.480 -0.115 3.600 0.210 ;
        RECT  2.620 -0.115 3.480 0.115 ;
        RECT  2.500 -0.115 2.620 0.130 ;
        RECT  2.050 -0.115 2.500 0.115 ;
        RECT  1.935 -0.115 2.050 0.265 ;
        RECT  1.655 -0.115 1.935 0.115 ;
        RECT  1.585 -0.115 1.655 0.420 ;
        RECT  0.315 -0.115 1.585 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.145 5.600 1.375 ;
        RECT  5.445 0.670 5.530 1.375 ;
        RECT  5.075 1.145 5.445 1.375 ;
        RECT  5.005 0.835 5.075 1.375 ;
        RECT  4.710 1.145 5.005 1.375 ;
        RECT  4.640 0.950 4.710 1.375 ;
        RECT  3.945 1.145 4.640 1.375 ;
        RECT  3.875 0.700 3.945 1.375 ;
        RECT  3.575 1.145 3.875 1.375 ;
        RECT  3.505 0.865 3.575 1.375 ;
        RECT  2.600 1.145 3.505 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.035 1.145 2.480 1.375 ;
        RECT  1.965 1.025 2.035 1.375 ;
        RECT  1.675 1.145 1.965 1.375 ;
        RECT  1.605 1.025 1.675 1.375 ;
        RECT  0.930 1.145 1.605 1.375 ;
        RECT  0.810 1.110 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.005 0.395 5.075 0.755 ;
        RECT  4.895 0.395 5.005 0.465 ;
        RECT  4.895 0.685 5.005 0.755 ;
        RECT  4.570 0.545 4.900 0.615 ;
        RECT  4.825 0.210 4.895 0.465 ;
        RECT  4.825 0.685 4.895 1.070 ;
        RECT  4.510 0.395 4.825 0.465 ;
        RECT  4.500 0.545 4.570 1.045 ;
        RECT  4.425 0.545 4.500 0.615 ;
        RECT  4.220 0.975 4.500 1.045 ;
        RECT  4.360 0.770 4.430 0.890 ;
        RECT  4.345 0.240 4.425 0.615 ;
        RECT  4.250 0.770 4.360 0.840 ;
        RECT  4.220 0.240 4.345 0.310 ;
        RECT  4.180 0.440 4.250 0.840 ;
        RECT  3.710 0.300 3.780 0.980 ;
        RECT  3.695 0.300 3.710 0.415 ;
        RECT  3.695 0.720 3.710 0.980 ;
        RECT  3.505 0.720 3.695 0.790 ;
        RECT  3.625 0.470 3.640 0.590 ;
        RECT  3.555 0.280 3.625 0.590 ;
        RECT  3.165 0.280 3.555 0.350 ;
        RECT  3.435 0.670 3.505 0.790 ;
        RECT  3.345 0.420 3.395 0.490 ;
        RECT  3.345 0.885 3.390 0.955 ;
        RECT  3.275 0.420 3.345 0.955 ;
        RECT  3.095 0.280 3.165 0.965 ;
        RECT  2.215 0.205 2.995 0.275 ;
        RECT  2.905 0.865 2.975 1.060 ;
        RECT  2.845 0.355 2.915 0.795 ;
        RECT  2.140 0.990 2.905 1.060 ;
        RECT  2.695 0.355 2.845 0.425 ;
        RECT  2.695 0.725 2.845 0.795 ;
        RECT  2.625 0.545 2.715 0.615 ;
        RECT  2.555 0.355 2.625 0.850 ;
        RECT  2.300 0.355 2.555 0.425 ;
        RECT  2.325 0.780 2.555 0.850 ;
        RECT  2.145 0.205 2.215 0.410 ;
        RECT  2.135 0.510 2.205 0.920 ;
        RECT  1.265 0.850 2.135 0.920 ;
        RECT  1.810 0.710 1.890 0.780 ;
        RECT  1.810 0.190 1.835 0.310 ;
        RECT  1.740 0.190 1.810 0.780 ;
        RECT  1.425 0.710 1.740 0.780 ;
        RECT  1.345 0.640 1.425 0.780 ;
        RECT  1.195 0.195 1.265 0.920 ;
        RECT  1.030 0.235 1.105 1.030 ;
        RECT  1.005 0.235 1.030 0.405 ;
        RECT  0.610 0.960 1.030 1.030 ;
        RECT  0.610 0.335 1.005 0.405 ;
        RECT  0.410 0.195 0.920 0.265 ;
        RECT  0.385 0.625 0.805 0.695 ;
        RECT  0.315 0.625 0.385 0.975 ;
        RECT  0.275 0.625 0.315 0.695 ;
        RECT  0.125 0.905 0.315 0.975 ;
        RECT  0.195 0.355 0.275 0.695 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.905 0.125 1.075 ;
    END
END SDFKCSNQD2BWP40

MACRO SDFKCSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFKCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.125 0.765 0.230 0.835 ;
        RECT  0.035 0.495 0.125 0.835 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.500 1.635 0.570 ;
        RECT  1.425 0.215 1.505 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.028400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.355 2.065 0.640 ;
        RECT  1.880 0.520 1.930 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.825 0.205 5.915 0.465 ;
        RECT  5.825 0.685 5.915 1.075 ;
        RECT  5.775 0.380 5.825 0.465 ;
        RECT  5.775 0.685 5.825 0.770 ;
        RECT  5.565 0.380 5.775 0.770 ;
        RECT  5.555 0.380 5.565 0.465 ;
        RECT  5.555 0.685 5.565 0.770 ;
        RECT  5.465 0.205 5.555 0.465 ;
        RECT  5.465 0.685 5.555 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 0.765 0.595 0.835 ;
        RECT  0.455 0.765 0.525 1.045 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.495 2.485 0.625 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.014800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.875 0.475 0.945 0.875 ;
        RECT  0.435 0.475 0.875 0.545 ;
        RECT  0.735 0.805 0.875 0.875 ;
        RECT  0.355 0.410 0.435 0.545 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 -0.115 6.160 0.115 ;
        RECT  6.035 -0.115 6.105 0.445 ;
        RECT  5.725 -0.115 6.035 0.115 ;
        RECT  5.655 -0.115 5.725 0.255 ;
        RECT  5.345 -0.115 5.655 0.115 ;
        RECT  5.275 -0.115 5.345 0.305 ;
        RECT  4.965 -0.115 5.275 0.115 ;
        RECT  4.895 -0.115 4.965 0.305 ;
        RECT  4.145 -0.115 4.895 0.115 ;
        RECT  4.075 -0.115 4.145 0.380 ;
        RECT  3.600 -0.115 4.075 0.115 ;
        RECT  3.480 -0.115 3.600 0.210 ;
        RECT  2.620 -0.115 3.480 0.115 ;
        RECT  2.500 -0.115 2.620 0.130 ;
        RECT  2.050 -0.115 2.500 0.115 ;
        RECT  1.930 -0.115 2.050 0.265 ;
        RECT  1.655 -0.115 1.930 0.115 ;
        RECT  1.585 -0.115 1.655 0.420 ;
        RECT  0.315 -0.115 1.585 0.115 ;
        RECT  0.245 -0.115 0.315 0.285 ;
        RECT  0.000 -0.115 0.245 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.105 1.145 6.160 1.375 ;
        RECT  6.035 0.715 6.105 1.375 ;
        RECT  5.725 1.145 6.035 1.375 ;
        RECT  5.655 0.885 5.725 1.375 ;
        RECT  5.345 1.145 5.655 1.375 ;
        RECT  5.275 0.715 5.345 1.375 ;
        RECT  4.970 1.145 5.275 1.375 ;
        RECT  4.900 0.950 4.970 1.375 ;
        RECT  4.145 1.145 4.900 1.375 ;
        RECT  4.075 0.740 4.145 1.375 ;
        RECT  3.575 1.145 4.075 1.375 ;
        RECT  3.505 0.865 3.575 1.375 ;
        RECT  2.600 1.145 3.505 1.375 ;
        RECT  2.480 1.135 2.600 1.375 ;
        RECT  2.035 1.145 2.480 1.375 ;
        RECT  1.965 1.025 2.035 1.375 ;
        RECT  1.675 1.145 1.965 1.375 ;
        RECT  1.605 1.025 1.675 1.375 ;
        RECT  0.930 1.145 1.605 1.375 ;
        RECT  0.810 1.110 0.930 1.375 ;
        RECT  0.340 1.145 0.810 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.845 0.205 5.915 0.465 ;
        RECT  5.845 0.685 5.915 1.075 ;
        RECT  5.465 0.205 5.495 0.465 ;
        RECT  5.465 0.685 5.495 1.075 ;
        RECT  5.155 0.395 5.205 0.785 ;
        RECT  5.135 0.185 5.155 1.070 ;
        RECT  5.085 0.185 5.135 0.465 ;
        RECT  5.085 0.715 5.135 1.070 ;
        RECT  4.780 0.395 5.085 0.465 ;
        RECT  4.830 0.545 5.065 0.615 ;
        RECT  4.760 0.545 4.830 1.050 ;
        RECT  4.710 0.545 4.760 0.615 ;
        RECT  4.490 0.980 4.760 1.050 ;
        RECT  4.630 0.240 4.710 0.615 ;
        RECT  4.620 0.780 4.690 0.900 ;
        RECT  4.490 0.240 4.630 0.310 ;
        RECT  4.520 0.780 4.620 0.850 ;
        RECT  4.450 0.440 4.520 0.850 ;
        RECT  4.275 0.315 4.345 0.520 ;
        RECT  4.275 0.600 4.345 0.955 ;
        RECT  3.945 0.450 4.275 0.520 ;
        RECT  3.945 0.600 4.275 0.670 ;
        RECT  3.875 0.315 3.945 0.520 ;
        RECT  3.875 0.600 3.945 0.955 ;
        RECT  3.710 0.300 3.780 0.980 ;
        RECT  3.695 0.300 3.710 0.415 ;
        RECT  3.695 0.720 3.710 0.980 ;
        RECT  3.505 0.720 3.695 0.790 ;
        RECT  3.625 0.470 3.640 0.590 ;
        RECT  3.555 0.280 3.625 0.590 ;
        RECT  3.165 0.280 3.555 0.350 ;
        RECT  3.435 0.670 3.505 0.790 ;
        RECT  3.345 0.420 3.395 0.490 ;
        RECT  3.345 0.885 3.390 0.955 ;
        RECT  3.275 0.420 3.345 0.955 ;
        RECT  3.095 0.280 3.165 0.965 ;
        RECT  2.215 0.205 2.995 0.275 ;
        RECT  2.905 0.865 2.975 1.060 ;
        RECT  2.845 0.355 2.915 0.795 ;
        RECT  2.140 0.990 2.905 1.060 ;
        RECT  2.695 0.355 2.845 0.425 ;
        RECT  2.695 0.725 2.845 0.795 ;
        RECT  2.625 0.545 2.715 0.615 ;
        RECT  2.555 0.355 2.625 0.850 ;
        RECT  2.300 0.355 2.555 0.425 ;
        RECT  2.325 0.780 2.555 0.850 ;
        RECT  2.145 0.205 2.215 0.410 ;
        RECT  2.135 0.510 2.205 0.920 ;
        RECT  1.265 0.850 2.135 0.920 ;
        RECT  1.810 0.710 1.890 0.780 ;
        RECT  1.810 0.190 1.835 0.310 ;
        RECT  1.740 0.190 1.810 0.780 ;
        RECT  1.425 0.710 1.740 0.780 ;
        RECT  1.345 0.640 1.425 0.780 ;
        RECT  1.195 0.195 1.265 0.920 ;
        RECT  1.030 0.235 1.105 1.030 ;
        RECT  1.005 0.235 1.030 0.405 ;
        RECT  0.610 0.960 1.030 1.030 ;
        RECT  0.610 0.335 1.005 0.405 ;
        RECT  0.410 0.195 0.920 0.265 ;
        RECT  0.385 0.625 0.805 0.695 ;
        RECT  0.315 0.625 0.385 0.975 ;
        RECT  0.275 0.625 0.315 0.695 ;
        RECT  0.125 0.905 0.315 0.975 ;
        RECT  0.195 0.355 0.275 0.695 ;
        RECT  0.145 0.355 0.195 0.425 ;
        RECT  0.055 0.185 0.145 0.425 ;
        RECT  0.055 0.905 0.125 1.075 ;
    END
END SDFKCSNQD4BWP40

MACRO SDFKSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFKSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.495 1.440 0.625 ;
        RECT  1.225 0.495 1.320 0.565 ;
        RECT  1.155 0.215 1.225 0.565 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.810 0.640 ;
        RECT  1.690 0.505 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.055 0.195 5.145 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.755 0.680 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.285 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 -0.115 5.180 0.115 ;
        RECT  4.865 -0.115 4.935 0.315 ;
        RECT  4.565 -0.115 4.865 0.115 ;
        RECT  4.495 -0.115 4.565 0.315 ;
        RECT  3.795 -0.115 4.495 0.115 ;
        RECT  3.725 -0.115 3.795 0.435 ;
        RECT  3.420 -0.115 3.725 0.115 ;
        RECT  3.300 -0.115 3.420 0.210 ;
        RECT  2.410 -0.115 3.300 0.115 ;
        RECT  2.290 -0.115 2.410 0.125 ;
        RECT  1.860 -0.115 2.290 0.115 ;
        RECT  1.740 -0.115 1.860 0.270 ;
        RECT  1.465 -0.115 1.740 0.115 ;
        RECT  1.395 -0.115 1.465 0.420 ;
        RECT  0.685 -0.115 1.395 0.115 ;
        RECT  0.615 -0.115 0.685 0.285 ;
        RECT  0.340 -0.115 0.615 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 1.145 5.180 1.375 ;
        RECT  4.865 0.945 4.935 1.375 ;
        RECT  4.565 1.145 4.865 1.375 ;
        RECT  4.495 0.950 4.565 1.375 ;
        RECT  3.795 1.145 4.495 1.375 ;
        RECT  3.725 0.785 3.795 1.375 ;
        RECT  3.415 1.145 3.725 1.375 ;
        RECT  3.305 0.890 3.415 1.375 ;
        RECT  2.430 1.145 3.305 1.375 ;
        RECT  2.310 1.140 2.430 1.375 ;
        RECT  1.870 1.145 2.310 1.375 ;
        RECT  1.750 1.110 1.870 1.375 ;
        RECT  1.530 1.145 1.750 1.375 ;
        RECT  1.410 1.020 1.530 1.375 ;
        RECT  0.340 1.145 1.410 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.395 4.935 0.820 ;
        RECT  4.755 0.395 4.865 0.465 ;
        RECT  4.755 0.750 4.865 0.820 ;
        RECT  4.425 0.545 4.760 0.615 ;
        RECT  4.685 0.195 4.755 0.465 ;
        RECT  4.685 0.750 4.755 1.070 ;
        RECT  4.370 0.395 4.685 0.465 ;
        RECT  4.355 0.545 4.425 1.045 ;
        RECT  4.290 0.545 4.355 0.615 ;
        RECT  4.070 0.975 4.355 1.045 ;
        RECT  4.220 0.225 4.290 0.615 ;
        RECT  4.215 0.775 4.285 0.885 ;
        RECT  4.070 0.225 4.220 0.295 ;
        RECT  4.095 0.775 4.215 0.845 ;
        RECT  4.025 0.440 4.095 0.845 ;
        RECT  3.530 0.300 3.600 0.980 ;
        RECT  3.315 0.745 3.530 0.815 ;
        RECT  3.390 0.280 3.460 0.640 ;
        RECT  2.995 0.280 3.390 0.350 ;
        RECT  3.245 0.695 3.315 0.815 ;
        RECT  3.155 0.420 3.230 0.490 ;
        RECT  3.155 0.885 3.225 0.955 ;
        RECT  3.085 0.420 3.155 0.955 ;
        RECT  2.925 0.205 2.995 0.925 ;
        RECT  2.785 0.355 2.855 0.780 ;
        RECT  2.025 0.205 2.830 0.275 ;
        RECT  2.735 0.860 2.805 1.055 ;
        RECT  2.515 0.355 2.785 0.425 ;
        RECT  2.625 0.710 2.785 0.780 ;
        RECT  2.120 0.985 2.735 1.055 ;
        RECT  2.555 0.710 2.625 0.905 ;
        RECT  2.435 0.545 2.525 0.615 ;
        RECT  2.365 0.355 2.435 0.905 ;
        RECT  2.115 0.355 2.365 0.425 ;
        RECT  2.130 0.835 2.365 0.905 ;
        RECT  2.050 0.985 2.120 1.070 ;
        RECT  1.950 1.000 2.050 1.070 ;
        RECT  1.955 0.205 2.025 0.345 ;
        RECT  1.880 0.510 1.950 0.930 ;
        RECT  1.065 0.860 1.880 0.930 ;
        RECT  1.620 0.720 1.690 0.790 ;
        RECT  1.620 0.195 1.645 0.315 ;
        RECT  1.550 0.195 1.620 0.790 ;
        RECT  1.215 0.720 1.550 0.790 ;
        RECT  1.145 0.640 1.215 0.790 ;
        RECT  0.995 0.185 1.065 1.055 ;
        RECT  0.875 0.355 0.910 1.055 ;
        RECT  0.840 0.185 0.875 1.055 ;
        RECT  0.805 0.185 0.840 0.425 ;
        RECT  0.805 0.945 0.840 1.055 ;
        RECT  0.505 0.355 0.805 0.425 ;
        RECT  0.505 0.935 0.720 1.005 ;
        RECT  0.435 0.195 0.505 0.425 ;
        RECT  0.435 0.935 0.505 1.070 ;
        RECT  0.340 0.505 0.385 0.670 ;
        RECT  0.270 0.345 0.340 0.915 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.125 0.845 0.270 0.915 ;
        RECT  0.055 0.195 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.015 ;
    END
END SDFKSNQD0BWP40

MACRO SDFKSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFKSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.495 1.440 0.625 ;
        RECT  1.225 0.495 1.320 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.810 0.640 ;
        RECT  1.690 0.505 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.055 0.185 5.145 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.755 0.680 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.285 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 -0.115 5.180 0.115 ;
        RECT  4.865 -0.115 4.935 0.305 ;
        RECT  4.565 -0.115 4.865 0.115 ;
        RECT  4.495 -0.115 4.565 0.330 ;
        RECT  3.795 -0.115 4.495 0.115 ;
        RECT  3.725 -0.115 3.795 0.435 ;
        RECT  3.420 -0.115 3.725 0.115 ;
        RECT  3.300 -0.115 3.420 0.210 ;
        RECT  2.410 -0.115 3.300 0.115 ;
        RECT  2.290 -0.115 2.410 0.130 ;
        RECT  1.860 -0.115 2.290 0.115 ;
        RECT  1.740 -0.115 1.860 0.265 ;
        RECT  1.465 -0.115 1.740 0.115 ;
        RECT  1.365 -0.115 1.465 0.420 ;
        RECT  0.710 -0.115 1.365 0.115 ;
        RECT  0.570 -0.115 0.710 0.150 ;
        RECT  0.340 -0.115 0.570 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 1.145 5.180 1.375 ;
        RECT  4.865 0.835 4.935 1.375 ;
        RECT  4.570 1.145 4.865 1.375 ;
        RECT  4.500 0.950 4.570 1.375 ;
        RECT  3.795 1.145 4.500 1.375 ;
        RECT  3.725 0.690 3.795 1.375 ;
        RECT  3.395 1.145 3.725 1.375 ;
        RECT  3.325 0.865 3.395 1.375 ;
        RECT  2.450 1.145 3.325 1.375 ;
        RECT  2.330 1.115 2.450 1.375 ;
        RECT  1.870 1.145 2.330 1.375 ;
        RECT  1.750 1.110 1.870 1.375 ;
        RECT  1.520 1.145 1.750 1.375 ;
        RECT  1.400 1.010 1.520 1.375 ;
        RECT  0.340 1.145 1.400 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.405 4.935 0.755 ;
        RECT  4.755 0.405 4.865 0.475 ;
        RECT  4.755 0.685 4.865 0.755 ;
        RECT  4.685 0.210 4.755 0.475 ;
        RECT  4.685 0.685 4.755 1.070 ;
        RECT  4.430 0.545 4.735 0.615 ;
        RECT  4.370 0.405 4.685 0.475 ;
        RECT  4.360 0.545 4.430 1.045 ;
        RECT  4.290 0.545 4.360 0.615 ;
        RECT  4.070 0.975 4.360 1.045 ;
        RECT  4.210 0.240 4.290 0.615 ;
        RECT  4.210 0.770 4.280 0.890 ;
        RECT  4.070 0.240 4.210 0.310 ;
        RECT  4.100 0.770 4.210 0.840 ;
        RECT  4.030 0.440 4.100 0.840 ;
        RECT  3.530 0.300 3.600 0.980 ;
        RECT  3.515 0.300 3.530 0.415 ;
        RECT  3.515 0.720 3.530 0.980 ;
        RECT  3.325 0.720 3.515 0.790 ;
        RECT  3.445 0.470 3.460 0.590 ;
        RECT  3.375 0.280 3.445 0.590 ;
        RECT  2.995 0.280 3.375 0.350 ;
        RECT  3.255 0.670 3.325 0.790 ;
        RECT  3.165 0.420 3.220 0.490 ;
        RECT  3.165 0.885 3.210 0.955 ;
        RECT  3.095 0.420 3.165 0.955 ;
        RECT  2.925 0.280 2.995 0.980 ;
        RECT  2.025 0.205 2.835 0.275 ;
        RECT  2.780 0.865 2.835 0.935 ;
        RECT  2.710 0.865 2.780 1.045 ;
        RECT  2.160 0.975 2.710 1.045 ;
        RECT  2.625 0.355 2.695 0.765 ;
        RECT  2.515 0.355 2.625 0.425 ;
        RECT  2.555 0.695 2.625 0.890 ;
        RECT  2.435 0.545 2.540 0.620 ;
        RECT  2.365 0.355 2.435 0.905 ;
        RECT  2.110 0.355 2.365 0.425 ;
        RECT  2.130 0.835 2.365 0.905 ;
        RECT  2.090 0.975 2.160 1.070 ;
        RECT  1.950 1.000 2.090 1.070 ;
        RECT  1.955 0.205 2.025 0.410 ;
        RECT  1.890 0.510 1.960 0.930 ;
        RECT  1.065 0.860 1.890 0.930 ;
        RECT  1.605 0.720 1.690 0.790 ;
        RECT  1.605 0.190 1.645 0.310 ;
        RECT  1.535 0.190 1.605 0.790 ;
        RECT  1.225 0.720 1.535 0.790 ;
        RECT  1.135 0.640 1.225 0.790 ;
        RECT  0.995 0.210 1.065 1.060 ;
        RECT  0.875 0.280 0.910 0.840 ;
        RECT  0.840 0.280 0.875 1.060 ;
        RECT  0.505 0.280 0.840 0.350 ;
        RECT  0.805 0.770 0.840 1.060 ;
        RECT  0.615 0.770 0.685 1.025 ;
        RECT  0.505 0.860 0.615 0.930 ;
        RECT  0.435 0.185 0.505 0.350 ;
        RECT  0.435 0.770 0.505 1.025 ;
        RECT  0.340 0.505 0.385 0.670 ;
        RECT  0.270 0.345 0.340 0.915 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.125 0.845 0.270 0.915 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFKSNQD1BWP40

MACRO SDFKSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFKSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.460 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.495 1.440 0.625 ;
        RECT  1.225 0.495 1.320 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.810 0.640 ;
        RECT  1.690 0.505 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.065 0.185 5.155 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.755 0.680 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.285 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.390 -0.115 5.460 0.115 ;
        RECT  5.305 -0.115 5.390 0.470 ;
        RECT  4.935 -0.115 5.305 0.115 ;
        RECT  4.865 -0.115 4.935 0.305 ;
        RECT  4.565 -0.115 4.865 0.115 ;
        RECT  4.495 -0.115 4.565 0.330 ;
        RECT  3.795 -0.115 4.495 0.115 ;
        RECT  3.725 -0.115 3.795 0.435 ;
        RECT  3.420 -0.115 3.725 0.115 ;
        RECT  3.300 -0.115 3.420 0.210 ;
        RECT  2.410 -0.115 3.300 0.115 ;
        RECT  2.290 -0.115 2.410 0.130 ;
        RECT  1.860 -0.115 2.290 0.115 ;
        RECT  1.740 -0.115 1.860 0.265 ;
        RECT  1.465 -0.115 1.740 0.115 ;
        RECT  1.365 -0.115 1.465 0.420 ;
        RECT  0.710 -0.115 1.365 0.115 ;
        RECT  0.570 -0.115 0.710 0.150 ;
        RECT  0.340 -0.115 0.570 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.390 1.145 5.460 1.375 ;
        RECT  5.305 0.670 5.390 1.375 ;
        RECT  4.935 1.145 5.305 1.375 ;
        RECT  4.865 0.835 4.935 1.375 ;
        RECT  4.570 1.145 4.865 1.375 ;
        RECT  4.500 0.950 4.570 1.375 ;
        RECT  3.795 1.145 4.500 1.375 ;
        RECT  3.725 0.690 3.795 1.375 ;
        RECT  3.395 1.145 3.725 1.375 ;
        RECT  3.325 0.865 3.395 1.375 ;
        RECT  2.450 1.145 3.325 1.375 ;
        RECT  2.330 1.115 2.450 1.375 ;
        RECT  1.870 1.145 2.330 1.375 ;
        RECT  1.750 1.110 1.870 1.375 ;
        RECT  1.520 1.145 1.750 1.375 ;
        RECT  1.400 1.010 1.520 1.375 ;
        RECT  0.340 1.145 1.400 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.865 0.405 4.935 0.755 ;
        RECT  4.755 0.405 4.865 0.475 ;
        RECT  4.755 0.685 4.865 0.755 ;
        RECT  4.685 0.210 4.755 0.475 ;
        RECT  4.685 0.685 4.755 1.070 ;
        RECT  4.430 0.545 4.735 0.615 ;
        RECT  4.370 0.405 4.685 0.475 ;
        RECT  4.360 0.545 4.430 1.045 ;
        RECT  4.290 0.545 4.360 0.615 ;
        RECT  4.070 0.975 4.360 1.045 ;
        RECT  4.210 0.240 4.290 0.615 ;
        RECT  4.210 0.770 4.280 0.890 ;
        RECT  4.070 0.240 4.210 0.310 ;
        RECT  4.100 0.770 4.210 0.840 ;
        RECT  4.030 0.440 4.100 0.840 ;
        RECT  3.530 0.300 3.600 0.980 ;
        RECT  3.515 0.300 3.530 0.415 ;
        RECT  3.515 0.720 3.530 0.980 ;
        RECT  3.325 0.720 3.515 0.790 ;
        RECT  3.445 0.470 3.460 0.590 ;
        RECT  3.375 0.280 3.445 0.590 ;
        RECT  2.995 0.280 3.375 0.350 ;
        RECT  3.255 0.670 3.325 0.790 ;
        RECT  3.165 0.420 3.220 0.490 ;
        RECT  3.165 0.885 3.210 0.955 ;
        RECT  3.095 0.420 3.165 0.955 ;
        RECT  2.925 0.280 2.995 0.980 ;
        RECT  2.025 0.205 2.835 0.275 ;
        RECT  2.780 0.865 2.835 0.935 ;
        RECT  2.710 0.865 2.780 1.045 ;
        RECT  2.160 0.975 2.710 1.045 ;
        RECT  2.625 0.355 2.695 0.765 ;
        RECT  2.515 0.355 2.625 0.425 ;
        RECT  2.555 0.695 2.625 0.890 ;
        RECT  2.435 0.545 2.540 0.620 ;
        RECT  2.365 0.355 2.435 0.905 ;
        RECT  2.110 0.355 2.365 0.425 ;
        RECT  2.130 0.835 2.365 0.905 ;
        RECT  2.090 0.975 2.160 1.070 ;
        RECT  1.950 1.000 2.090 1.070 ;
        RECT  1.955 0.205 2.025 0.410 ;
        RECT  1.890 0.510 1.960 0.930 ;
        RECT  1.065 0.860 1.890 0.930 ;
        RECT  1.605 0.720 1.690 0.790 ;
        RECT  1.605 0.190 1.645 0.310 ;
        RECT  1.535 0.190 1.605 0.790 ;
        RECT  1.225 0.720 1.535 0.790 ;
        RECT  1.135 0.640 1.225 0.790 ;
        RECT  0.995 0.210 1.065 1.060 ;
        RECT  0.875 0.280 0.910 0.840 ;
        RECT  0.840 0.280 0.875 1.060 ;
        RECT  0.505 0.280 0.840 0.350 ;
        RECT  0.805 0.770 0.840 1.060 ;
        RECT  0.615 0.770 0.685 1.025 ;
        RECT  0.505 0.860 0.615 0.930 ;
        RECT  0.435 0.185 0.505 0.350 ;
        RECT  0.435 0.770 0.505 1.025 ;
        RECT  0.340 0.505 0.385 0.670 ;
        RECT  0.270 0.345 0.340 0.915 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.125 0.845 0.270 0.915 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFKSNQD2BWP40

MACRO SDFKSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFKSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.190 0.765 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.495 1.440 0.625 ;
        RECT  1.225 0.495 1.320 0.570 ;
        RECT  1.155 0.215 1.225 0.570 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.715 0.355 1.810 0.640 ;
        RECT  1.690 0.505 1.715 0.640 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.685 0.205 5.775 0.465 ;
        RECT  5.685 0.685 5.775 1.075 ;
        RECT  5.635 0.380 5.685 0.465 ;
        RECT  5.635 0.685 5.685 0.770 ;
        RECT  5.425 0.380 5.635 0.770 ;
        RECT  5.415 0.380 5.425 0.465 ;
        RECT  5.415 0.685 5.425 0.770 ;
        RECT  5.325 0.205 5.415 0.465 ;
        RECT  5.325 0.685 5.415 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.495 0.755 0.680 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 0.495 2.285 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.965 -0.115 6.020 0.115 ;
        RECT  5.895 -0.115 5.965 0.445 ;
        RECT  5.585 -0.115 5.895 0.115 ;
        RECT  5.515 -0.115 5.585 0.255 ;
        RECT  5.205 -0.115 5.515 0.115 ;
        RECT  5.135 -0.115 5.205 0.305 ;
        RECT  4.825 -0.115 5.135 0.115 ;
        RECT  4.755 -0.115 4.825 0.305 ;
        RECT  4.005 -0.115 4.755 0.115 ;
        RECT  3.935 -0.115 4.005 0.380 ;
        RECT  3.420 -0.115 3.935 0.115 ;
        RECT  3.300 -0.115 3.420 0.210 ;
        RECT  2.410 -0.115 3.300 0.115 ;
        RECT  2.290 -0.115 2.410 0.130 ;
        RECT  1.860 -0.115 2.290 0.115 ;
        RECT  1.740 -0.115 1.860 0.265 ;
        RECT  1.465 -0.115 1.740 0.115 ;
        RECT  1.365 -0.115 1.465 0.420 ;
        RECT  0.710 -0.115 1.365 0.115 ;
        RECT  0.570 -0.115 0.710 0.150 ;
        RECT  0.340 -0.115 0.570 0.115 ;
        RECT  0.220 -0.115 0.340 0.275 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.965 1.145 6.020 1.375 ;
        RECT  5.895 0.715 5.965 1.375 ;
        RECT  5.585 1.145 5.895 1.375 ;
        RECT  5.515 0.885 5.585 1.375 ;
        RECT  5.205 1.145 5.515 1.375 ;
        RECT  5.135 0.715 5.205 1.375 ;
        RECT  4.830 1.145 5.135 1.375 ;
        RECT  4.760 0.950 4.830 1.375 ;
        RECT  4.005 1.145 4.760 1.375 ;
        RECT  3.935 0.740 4.005 1.375 ;
        RECT  3.395 1.145 3.935 1.375 ;
        RECT  3.325 0.865 3.395 1.375 ;
        RECT  2.450 1.145 3.325 1.375 ;
        RECT  2.330 1.115 2.450 1.375 ;
        RECT  1.870 1.145 2.330 1.375 ;
        RECT  1.750 1.110 1.870 1.375 ;
        RECT  1.520 1.145 1.750 1.375 ;
        RECT  1.400 1.010 1.520 1.375 ;
        RECT  0.340 1.145 1.400 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.705 0.205 5.775 0.465 ;
        RECT  5.705 0.685 5.775 1.075 ;
        RECT  5.325 0.205 5.355 0.465 ;
        RECT  5.325 0.685 5.355 1.075 ;
        RECT  5.015 0.395 5.065 0.785 ;
        RECT  4.995 0.185 5.015 1.070 ;
        RECT  4.945 0.185 4.995 0.465 ;
        RECT  4.945 0.715 4.995 1.070 ;
        RECT  4.640 0.395 4.945 0.465 ;
        RECT  4.690 0.545 4.925 0.615 ;
        RECT  4.620 0.545 4.690 1.050 ;
        RECT  4.570 0.545 4.620 0.615 ;
        RECT  4.350 0.980 4.620 1.050 ;
        RECT  4.490 0.240 4.570 0.615 ;
        RECT  4.480 0.780 4.550 0.900 ;
        RECT  4.350 0.240 4.490 0.310 ;
        RECT  4.380 0.780 4.480 0.850 ;
        RECT  4.310 0.440 4.380 0.850 ;
        RECT  4.135 0.315 4.205 0.520 ;
        RECT  4.135 0.600 4.205 0.955 ;
        RECT  3.805 0.450 4.135 0.520 ;
        RECT  3.805 0.600 4.135 0.670 ;
        RECT  3.735 0.315 3.805 0.520 ;
        RECT  3.735 0.600 3.805 0.955 ;
        RECT  3.530 0.300 3.600 0.980 ;
        RECT  3.515 0.300 3.530 0.415 ;
        RECT  3.515 0.720 3.530 0.980 ;
        RECT  3.325 0.720 3.515 0.790 ;
        RECT  3.445 0.470 3.460 0.590 ;
        RECT  3.375 0.280 3.445 0.590 ;
        RECT  2.995 0.280 3.375 0.350 ;
        RECT  3.255 0.670 3.325 0.790 ;
        RECT  3.165 0.420 3.220 0.490 ;
        RECT  3.165 0.885 3.210 0.955 ;
        RECT  3.095 0.420 3.165 0.955 ;
        RECT  2.925 0.280 2.995 0.980 ;
        RECT  2.025 0.205 2.835 0.275 ;
        RECT  2.780 0.865 2.835 0.935 ;
        RECT  2.710 0.865 2.780 1.045 ;
        RECT  2.160 0.975 2.710 1.045 ;
        RECT  2.625 0.355 2.695 0.765 ;
        RECT  2.515 0.355 2.625 0.425 ;
        RECT  2.555 0.695 2.625 0.890 ;
        RECT  2.435 0.545 2.540 0.620 ;
        RECT  2.365 0.355 2.435 0.905 ;
        RECT  2.110 0.355 2.365 0.425 ;
        RECT  2.130 0.835 2.365 0.905 ;
        RECT  2.090 0.975 2.160 1.070 ;
        RECT  1.950 1.000 2.090 1.070 ;
        RECT  1.955 0.205 2.025 0.410 ;
        RECT  1.890 0.510 1.960 0.930 ;
        RECT  1.065 0.860 1.890 0.930 ;
        RECT  1.605 0.720 1.690 0.790 ;
        RECT  1.605 0.190 1.645 0.310 ;
        RECT  1.535 0.190 1.605 0.790 ;
        RECT  1.225 0.720 1.535 0.790 ;
        RECT  1.135 0.640 1.225 0.790 ;
        RECT  0.995 0.210 1.065 1.060 ;
        RECT  0.875 0.280 0.910 0.840 ;
        RECT  0.840 0.280 0.875 1.060 ;
        RECT  0.505 0.280 0.840 0.350 ;
        RECT  0.805 0.770 0.840 1.060 ;
        RECT  0.615 0.770 0.685 1.025 ;
        RECT  0.505 0.860 0.615 0.930 ;
        RECT  0.435 0.185 0.505 0.350 ;
        RECT  0.435 0.770 0.505 1.025 ;
        RECT  0.340 0.505 0.385 0.670 ;
        RECT  0.270 0.345 0.340 0.915 ;
        RECT  0.125 0.345 0.270 0.415 ;
        RECT  0.125 0.845 0.270 0.915 ;
        RECT  0.055 0.185 0.125 0.415 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFKSNQD4BWP40

MACRO SDFMQD0BWP40
    CLASS CORE ;
    FOREIGN SDFMQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.275 0.475 2.360 0.810 ;
        RECT  2.220 0.475 2.275 0.635 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.062000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.045 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.305 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.355 1.995 0.595 ;
        RECT  1.570 0.505 1.800 0.595 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.530 0.495 2.765 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.315 -0.115 5.600 0.115 ;
        RECT  5.245 -0.115 5.315 0.315 ;
        RECT  4.945 -0.115 5.245 0.115 ;
        RECT  4.875 -0.115 4.945 0.315 ;
        RECT  4.225 -0.115 4.875 0.115 ;
        RECT  4.080 -0.115 4.225 0.125 ;
        RECT  3.530 -0.115 4.080 0.115 ;
        RECT  3.410 -0.115 3.530 0.125 ;
        RECT  2.750 -0.115 3.410 0.115 ;
        RECT  2.625 -0.115 2.750 0.140 ;
        RECT  2.420 -0.115 2.625 0.115 ;
        RECT  2.300 -0.115 2.420 0.125 ;
        RECT  0.945 -0.115 2.300 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.315 1.145 5.600 1.375 ;
        RECT  5.245 0.935 5.315 1.375 ;
        RECT  4.940 1.145 5.245 1.375 ;
        RECT  4.810 1.130 4.940 1.375 ;
        RECT  4.150 1.145 4.810 1.375 ;
        RECT  4.030 0.970 4.150 1.375 ;
        RECT  3.565 1.145 4.030 1.375 ;
        RECT  3.445 0.870 3.565 1.375 ;
        RECT  2.420 1.145 3.445 1.375 ;
        RECT  2.300 1.130 2.420 1.375 ;
        RECT  0.950 1.145 2.300 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 1.010 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.395 5.355 0.810 ;
        RECT  5.135 0.395 5.285 0.465 ;
        RECT  5.135 0.740 5.285 0.810 ;
        RECT  4.985 0.545 5.185 0.615 ;
        RECT  5.065 0.185 5.135 0.465 ;
        RECT  5.065 0.740 5.135 1.025 ;
        RECT  4.835 0.395 5.065 0.465 ;
        RECT  4.915 0.545 4.985 0.930 ;
        RECT  4.515 0.860 4.915 0.930 ;
        RECT  4.765 0.395 4.835 0.600 ;
        RECT  4.615 0.195 4.695 0.780 ;
        RECT  4.450 0.195 4.615 0.265 ;
        RECT  4.435 0.350 4.515 0.930 ;
        RECT  4.340 0.185 4.450 0.265 ;
        RECT  4.320 0.185 4.340 0.890 ;
        RECT  4.270 0.195 4.320 0.890 ;
        RECT  3.170 0.195 4.270 0.265 ;
        RECT  3.835 0.785 4.270 0.890 ;
        RECT  3.800 0.520 4.190 0.640 ;
        RECT  3.660 0.335 3.730 0.880 ;
        RECT  3.395 0.570 3.660 0.690 ;
        RECT  3.315 0.345 3.345 0.480 ;
        RECT  3.315 0.800 3.335 0.925 ;
        RECT  3.245 0.345 3.315 0.925 ;
        RECT  3.070 0.995 3.260 1.065 ;
        RECT  3.085 0.350 3.155 0.760 ;
        RECT  3.030 0.690 3.085 0.760 ;
        RECT  3.000 0.845 3.070 1.065 ;
        RECT  2.940 0.845 3.000 0.915 ;
        RECT  2.940 0.210 2.985 0.505 ;
        RECT  2.870 0.210 2.940 0.915 ;
        RECT  2.720 0.985 2.880 1.075 ;
        RECT  2.565 0.210 2.870 0.280 ;
        RECT  2.445 0.845 2.870 0.915 ;
        RECT  0.455 0.985 2.720 1.055 ;
        RECT  2.450 0.210 2.565 0.390 ;
        RECT  2.150 0.335 2.235 0.405 ;
        RECT  2.150 0.715 2.200 0.915 ;
        RECT  2.080 0.335 2.150 0.915 ;
        RECT  2.075 0.675 2.080 0.915 ;
        RECT  1.500 0.675 2.075 0.745 ;
        RECT  1.730 0.205 2.010 0.275 ;
        RECT  1.905 0.815 2.005 0.915 ;
        RECT  1.030 0.840 1.905 0.915 ;
        RECT  1.660 0.205 1.730 0.415 ;
        RECT  1.055 0.345 1.660 0.415 ;
        RECT  0.455 0.205 1.580 0.275 ;
        RECT  1.375 0.495 1.500 0.745 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  3.925 0.525 3.995 0.595 ;
        RECT  3.085 0.525 3.155 0.595 ;
        LAYER M2 ;
        RECT  3.030 0.525 4.045 0.595 ;
    END
END SDFMQD0BWP40

MACRO SDFMQD1BWP40
    CLASS CORE ;
    FOREIGN SDFMQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.030000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.265 0.475 2.350 0.810 ;
        RECT  2.210 0.475 2.265 0.635 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.124000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.305 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.355 1.985 0.595 ;
        RECT  1.570 0.505 1.800 0.595 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 0.495 2.765 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.315 -0.115 5.600 0.115 ;
        RECT  5.245 -0.115 5.315 0.315 ;
        RECT  4.945 -0.115 5.245 0.115 ;
        RECT  4.875 -0.115 4.945 0.315 ;
        RECT  4.115 -0.115 4.875 0.115 ;
        RECT  4.040 -0.115 4.115 0.265 ;
        RECT  3.525 -0.115 4.040 0.115 ;
        RECT  3.405 -0.115 3.525 0.125 ;
        RECT  2.740 -0.115 3.405 0.115 ;
        RECT  2.615 -0.115 2.740 0.140 ;
        RECT  2.410 -0.115 2.615 0.115 ;
        RECT  2.290 -0.115 2.410 0.125 ;
        RECT  0.945 -0.115 2.290 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.315 1.145 5.600 1.375 ;
        RECT  5.245 0.895 5.315 1.375 ;
        RECT  4.940 1.145 5.245 1.375 ;
        RECT  4.810 1.130 4.940 1.375 ;
        RECT  4.140 1.145 4.810 1.375 ;
        RECT  4.020 0.870 4.140 1.375 ;
        RECT  3.535 1.145 4.020 1.375 ;
        RECT  3.450 0.750 3.535 1.375 ;
        RECT  2.410 1.145 3.450 1.375 ;
        RECT  2.290 1.130 2.410 1.375 ;
        RECT  0.950 1.145 2.290 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 1.020 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.325 0.395 5.395 0.810 ;
        RECT  5.135 0.395 5.325 0.465 ;
        RECT  5.135 0.740 5.325 0.810 ;
        RECT  4.985 0.545 5.210 0.615 ;
        RECT  5.065 0.185 5.135 0.465 ;
        RECT  5.065 0.740 5.135 1.025 ;
        RECT  4.835 0.395 5.065 0.465 ;
        RECT  4.915 0.545 4.985 0.960 ;
        RECT  4.520 0.890 4.915 0.960 ;
        RECT  4.765 0.395 4.835 0.600 ;
        RECT  4.625 0.195 4.695 0.795 ;
        RECT  4.370 0.195 4.625 0.265 ;
        RECT  4.450 0.335 4.520 0.960 ;
        RECT  4.300 0.195 4.370 0.790 ;
        RECT  3.905 0.355 4.300 0.425 ;
        RECT  3.905 0.720 4.300 0.790 ;
        RECT  3.790 0.520 4.180 0.640 ;
        RECT  3.835 0.195 3.905 0.425 ;
        RECT  3.835 0.720 3.905 0.965 ;
        RECT  3.150 0.195 3.835 0.265 ;
        RECT  3.720 0.745 3.725 0.865 ;
        RECT  3.650 0.335 3.720 0.865 ;
        RECT  3.640 0.530 3.650 0.865 ;
        RECT  3.380 0.530 3.640 0.650 ;
        RECT  3.310 0.350 3.335 0.470 ;
        RECT  3.240 0.350 3.310 0.925 ;
        RECT  3.125 0.995 3.230 1.065 ;
        RECT  3.075 0.350 3.145 0.760 ;
        RECT  3.055 0.845 3.125 1.065 ;
        RECT  3.000 0.690 3.075 0.760 ;
        RECT  2.930 0.845 3.055 0.915 ;
        RECT  2.930 0.210 2.975 0.505 ;
        RECT  2.860 0.210 2.930 0.915 ;
        RECT  2.710 0.985 2.870 1.075 ;
        RECT  2.555 0.210 2.860 0.280 ;
        RECT  2.435 0.845 2.860 0.915 ;
        RECT  0.455 0.985 2.710 1.055 ;
        RECT  2.440 0.210 2.555 0.390 ;
        RECT  2.140 0.335 2.225 0.405 ;
        RECT  2.140 0.715 2.190 0.915 ;
        RECT  2.070 0.335 2.140 0.915 ;
        RECT  2.065 0.675 2.070 0.915 ;
        RECT  1.500 0.675 2.065 0.745 ;
        RECT  1.730 0.205 2.000 0.275 ;
        RECT  1.895 0.815 1.995 0.915 ;
        RECT  1.030 0.840 1.895 0.915 ;
        RECT  1.660 0.205 1.730 0.415 ;
        RECT  1.055 0.345 1.660 0.415 ;
        RECT  0.455 0.205 1.580 0.275 ;
        RECT  1.375 0.495 1.500 0.745 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  3.900 0.525 3.970 0.595 ;
        RECT  3.075 0.525 3.145 0.595 ;
        LAYER M2 ;
        RECT  3.025 0.525 4.020 0.595 ;
    END
END SDFMQD1BWP40

MACRO SDFMQD2BWP40
    CLASS CORE ;
    FOREIGN SDFMQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.030000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.475 2.345 0.810 ;
        RECT  2.200 0.475 2.255 0.635 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.144000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.495 0.195 5.570 1.065 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.305 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.355 1.975 0.595 ;
        RECT  1.570 0.505 1.800 0.595 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 0.495 2.765 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.815 -0.115 5.880 0.115 ;
        RECT  5.735 -0.115 5.815 0.465 ;
        RECT  5.315 -0.115 5.735 0.115 ;
        RECT  5.245 -0.115 5.315 0.315 ;
        RECT  4.945 -0.115 5.245 0.115 ;
        RECT  4.875 -0.115 4.945 0.280 ;
        RECT  4.105 -0.115 4.875 0.115 ;
        RECT  4.030 -0.115 4.105 0.265 ;
        RECT  3.520 -0.115 4.030 0.115 ;
        RECT  3.400 -0.115 3.520 0.125 ;
        RECT  2.730 -0.115 3.400 0.115 ;
        RECT  2.605 -0.115 2.730 0.140 ;
        RECT  2.400 -0.115 2.605 0.115 ;
        RECT  2.280 -0.115 2.400 0.125 ;
        RECT  0.945 -0.115 2.280 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.805 1.145 5.880 1.375 ;
        RECT  5.730 0.655 5.805 1.375 ;
        RECT  5.315 1.145 5.730 1.375 ;
        RECT  5.245 0.895 5.315 1.375 ;
        RECT  4.940 1.145 5.245 1.375 ;
        RECT  4.810 1.130 4.940 1.375 ;
        RECT  4.130 1.145 4.810 1.375 ;
        RECT  4.010 0.870 4.130 1.375 ;
        RECT  3.525 1.145 4.010 1.375 ;
        RECT  3.435 0.745 3.525 1.375 ;
        RECT  2.400 1.145 3.435 1.375 ;
        RECT  2.280 1.130 2.400 1.375 ;
        RECT  0.950 1.145 2.280 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 1.030 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.325 0.395 5.395 0.810 ;
        RECT  5.135 0.395 5.325 0.465 ;
        RECT  5.135 0.740 5.325 0.810 ;
        RECT  4.985 0.545 5.210 0.615 ;
        RECT  5.065 0.185 5.135 0.465 ;
        RECT  5.065 0.740 5.135 1.025 ;
        RECT  4.825 0.395 5.065 0.465 ;
        RECT  4.915 0.545 4.985 0.930 ;
        RECT  4.525 0.860 4.915 0.930 ;
        RECT  4.755 0.395 4.825 0.600 ;
        RECT  4.605 0.195 4.685 0.780 ;
        RECT  4.360 0.195 4.605 0.265 ;
        RECT  4.455 0.340 4.525 0.930 ;
        RECT  4.290 0.195 4.360 0.790 ;
        RECT  3.895 0.355 4.290 0.425 ;
        RECT  3.900 0.720 4.290 0.790 ;
        RECT  3.780 0.520 4.180 0.640 ;
        RECT  3.825 0.720 3.900 0.955 ;
        RECT  3.825 0.195 3.895 0.425 ;
        RECT  3.150 0.195 3.825 0.265 ;
        RECT  3.640 0.345 3.710 0.855 ;
        RECT  3.365 0.515 3.640 0.635 ;
        RECT  3.295 0.370 3.355 0.445 ;
        RECT  3.225 0.370 3.295 0.925 ;
        RECT  3.135 0.995 3.220 1.065 ;
        RECT  3.065 0.350 3.135 0.760 ;
        RECT  3.065 0.845 3.135 1.065 ;
        RECT  2.990 0.690 3.065 0.760 ;
        RECT  2.920 0.845 3.065 0.915 ;
        RECT  2.920 0.210 2.965 0.505 ;
        RECT  2.850 0.210 2.920 0.915 ;
        RECT  2.700 0.985 2.860 1.075 ;
        RECT  2.545 0.210 2.850 0.280 ;
        RECT  2.425 0.845 2.850 0.915 ;
        RECT  0.455 0.985 2.700 1.055 ;
        RECT  2.430 0.210 2.545 0.390 ;
        RECT  2.130 0.335 2.215 0.405 ;
        RECT  2.130 0.715 2.180 0.915 ;
        RECT  2.060 0.335 2.130 0.915 ;
        RECT  2.055 0.675 2.060 0.915 ;
        RECT  1.500 0.675 2.055 0.745 ;
        RECT  1.730 0.205 1.990 0.275 ;
        RECT  1.885 0.815 1.985 0.915 ;
        RECT  1.030 0.840 1.885 0.915 ;
        RECT  1.660 0.205 1.730 0.405 ;
        RECT  1.290 0.335 1.660 0.405 ;
        RECT  1.085 0.195 1.580 0.265 ;
        RECT  1.375 0.485 1.500 0.745 ;
        RECT  1.230 0.335 1.290 0.415 ;
        RECT  1.055 0.345 1.230 0.415 ;
        RECT  1.015 0.195 1.085 0.275 ;
        RECT  0.455 0.205 1.015 0.275 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  3.880 0.525 3.950 0.595 ;
        RECT  3.065 0.525 3.135 0.595 ;
        LAYER M2 ;
        RECT  3.015 0.525 4.000 0.595 ;
    END
END SDFMQD2BWP40

MACRO SDFMQD4BWP40
    CLASS CORE ;
    FOREIGN SDFMQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.030000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.475 2.345 0.810 ;
        RECT  2.200 0.475 2.255 0.635 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.745 6.025 0.995 ;
        RECT  5.915 0.195 6.020 0.465 ;
        RECT  5.705 0.355 5.915 0.880 ;
        RECT  5.615 0.355 5.705 0.480 ;
        RECT  5.615 0.710 5.705 0.880 ;
        RECT  5.545 0.195 5.615 0.480 ;
        RECT  5.545 0.710 5.615 0.990 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.085 0.495 1.305 0.765 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.018600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.355 1.975 0.595 ;
        RECT  1.570 0.505 1.800 0.595 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 0.495 2.765 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.210 -0.115 6.300 0.115 ;
        RECT  6.130 -0.115 6.210 0.460 ;
        RECT  5.810 -0.115 6.130 0.115 ;
        RECT  5.730 -0.115 5.810 0.250 ;
        RECT  5.425 -0.115 5.730 0.115 ;
        RECT  5.355 -0.115 5.425 0.315 ;
        RECT  5.045 -0.115 5.355 0.115 ;
        RECT  4.975 -0.115 5.045 0.315 ;
        RECT  4.150 -0.115 4.975 0.115 ;
        RECT  4.030 -0.115 4.150 0.235 ;
        RECT  3.520 -0.115 4.030 0.115 ;
        RECT  3.400 -0.115 3.520 0.125 ;
        RECT  2.730 -0.115 3.400 0.115 ;
        RECT  2.605 -0.115 2.730 0.140 ;
        RECT  2.400 -0.115 2.605 0.115 ;
        RECT  2.280 -0.115 2.400 0.125 ;
        RECT  0.945 -0.115 2.280 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.210 1.145 6.300 1.375 ;
        RECT  6.130 0.705 6.210 1.375 ;
        RECT  5.810 1.145 6.130 1.375 ;
        RECT  5.730 0.995 5.810 1.375 ;
        RECT  5.425 1.145 5.730 1.375 ;
        RECT  5.355 0.895 5.425 1.375 ;
        RECT  5.040 1.145 5.355 1.375 ;
        RECT  4.910 1.130 5.040 1.375 ;
        RECT  4.195 1.145 4.910 1.375 ;
        RECT  4.075 0.870 4.195 1.375 ;
        RECT  3.525 1.145 4.075 1.375 ;
        RECT  3.435 0.755 3.525 1.375 ;
        RECT  2.400 1.145 3.435 1.375 ;
        RECT  2.280 1.130 2.400 1.375 ;
        RECT  0.950 1.145 2.280 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 1.025 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.985 0.745 6.025 0.995 ;
        RECT  5.985 0.195 6.020 0.465 ;
        RECT  5.615 0.355 5.635 0.480 ;
        RECT  5.615 0.710 5.635 0.880 ;
        RECT  5.545 0.195 5.615 0.480 ;
        RECT  5.545 0.710 5.615 0.990 ;
        RECT  5.380 0.395 5.450 0.810 ;
        RECT  5.235 0.395 5.380 0.465 ;
        RECT  5.235 0.740 5.380 0.810 ;
        RECT  5.085 0.545 5.300 0.615 ;
        RECT  5.165 0.185 5.235 0.465 ;
        RECT  5.165 0.740 5.235 1.025 ;
        RECT  4.925 0.395 5.165 0.465 ;
        RECT  5.015 0.545 5.085 0.930 ;
        RECT  4.610 0.860 5.015 0.930 ;
        RECT  4.855 0.395 4.925 0.600 ;
        RECT  4.705 0.195 4.785 0.780 ;
        RECT  4.460 0.195 4.705 0.265 ;
        RECT  4.540 0.345 4.610 0.930 ;
        RECT  4.390 0.195 4.460 0.790 ;
        RECT  3.900 0.360 4.390 0.430 ;
        RECT  3.915 0.720 4.390 0.790 ;
        RECT  3.780 0.510 4.270 0.640 ;
        RECT  3.840 0.720 3.915 0.950 ;
        RECT  3.825 0.195 3.900 0.430 ;
        RECT  3.150 0.195 3.825 0.265 ;
        RECT  3.640 0.335 3.710 0.855 ;
        RECT  3.375 0.530 3.640 0.650 ;
        RECT  3.300 0.360 3.355 0.445 ;
        RECT  3.230 0.360 3.300 0.925 ;
        RECT  3.080 0.995 3.220 1.065 ;
        RECT  3.065 0.350 3.135 0.760 ;
        RECT  3.010 0.845 3.080 1.065 ;
        RECT  2.990 0.690 3.065 0.760 ;
        RECT  2.920 0.845 3.010 0.915 ;
        RECT  2.920 0.210 2.965 0.505 ;
        RECT  2.850 0.210 2.920 0.915 ;
        RECT  2.700 0.985 2.860 1.075 ;
        RECT  2.545 0.210 2.850 0.280 ;
        RECT  2.425 0.845 2.850 0.915 ;
        RECT  0.455 0.985 2.700 1.055 ;
        RECT  2.430 0.210 2.545 0.390 ;
        RECT  2.130 0.335 2.215 0.405 ;
        RECT  2.130 0.770 2.180 0.915 ;
        RECT  2.060 0.335 2.130 0.915 ;
        RECT  2.055 0.675 2.060 0.915 ;
        RECT  1.500 0.675 2.055 0.745 ;
        RECT  1.730 0.205 1.990 0.275 ;
        RECT  1.885 0.815 1.985 0.915 ;
        RECT  1.030 0.840 1.885 0.915 ;
        RECT  1.660 0.205 1.730 0.415 ;
        RECT  1.055 0.345 1.660 0.415 ;
        RECT  0.455 0.205 1.580 0.275 ;
        RECT  1.375 0.495 1.500 0.745 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  3.910 0.525 3.980 0.595 ;
        RECT  3.065 0.525 3.135 0.595 ;
        LAYER M2 ;
        RECT  3.015 0.525 4.030 0.595 ;
    END
END SDFMQD4BWP40

MACRO SDFNCNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.320 4.865 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.495 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.665 -0.115 4.900 0.115 ;
        RECT  4.540 -0.115 4.665 0.255 ;
        RECT  4.080 -0.115 4.540 0.115 ;
        RECT  4.005 -0.115 4.080 0.425 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.670 1.145 4.900 1.375 ;
        RECT  4.550 1.025 4.670 1.375 ;
        RECT  4.270 1.145 4.550 1.375 ;
        RECT  4.185 0.995 4.270 1.375 ;
        RECT  4.105 1.145 4.185 1.375 ;
        RECT  3.985 0.870 4.105 1.375 ;
        RECT  3.315 1.145 3.985 1.375 ;
        RECT  3.205 0.815 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.325 4.705 0.915 ;
        RECT  4.165 0.325 4.635 0.395 ;
        RECT  4.470 0.845 4.635 0.915 ;
        RECT  4.375 0.495 4.530 0.765 ;
        RECT  4.360 0.845 4.470 1.035 ;
        RECT  4.280 0.845 4.360 0.915 ;
        RECT  4.210 0.695 4.280 0.915 ;
        RECT  3.685 0.540 4.275 0.610 ;
        RECT  3.910 0.695 4.210 0.765 ;
        RECT  3.710 0.995 3.860 1.075 ;
        RECT  3.675 0.815 3.745 0.885 ;
        RECT  3.465 0.995 3.710 1.065 ;
        RECT  3.675 0.310 3.685 0.610 ;
        RECT  3.605 0.310 3.675 0.885 ;
        RECT  3.465 0.195 3.530 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.375 0.525 4.445 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQD0BWP40

MACRO SDFNCNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.185 4.865 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.035200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.495 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.680 -0.115 4.900 0.115 ;
        RECT  4.555 -0.115 4.680 0.255 ;
        RECT  4.080 -0.115 4.555 0.115 ;
        RECT  4.005 -0.115 4.080 0.425 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.670 1.145 4.900 1.375 ;
        RECT  4.550 1.025 4.670 1.375 ;
        RECT  4.270 1.145 4.550 1.375 ;
        RECT  4.185 0.995 4.270 1.375 ;
        RECT  4.105 1.145 4.185 1.375 ;
        RECT  3.985 0.870 4.105 1.375 ;
        RECT  3.315 1.145 3.985 1.375 ;
        RECT  3.205 0.860 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.325 4.705 0.915 ;
        RECT  4.165 0.325 4.635 0.395 ;
        RECT  4.280 0.845 4.635 0.915 ;
        RECT  4.375 0.495 4.530 0.765 ;
        RECT  4.210 0.695 4.280 0.915 ;
        RECT  3.685 0.540 4.275 0.610 ;
        RECT  3.910 0.695 4.210 0.765 ;
        RECT  3.710 0.995 3.860 1.075 ;
        RECT  3.675 0.815 3.745 0.885 ;
        RECT  3.465 0.995 3.710 1.065 ;
        RECT  3.675 0.310 3.685 0.610 ;
        RECT  3.605 0.310 3.675 0.885 ;
        RECT  3.465 0.195 3.530 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.375 0.525 4.445 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQD1BWP40

MACRO SDFNCNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.795 0.185 4.865 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.040800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.495 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.090 -0.115 5.180 0.115 ;
        RECT  5.020 -0.115 5.090 0.485 ;
        RECT  4.680 -0.115 5.020 0.115 ;
        RECT  4.555 -0.115 4.680 0.255 ;
        RECT  4.080 -0.115 4.555 0.115 ;
        RECT  4.005 -0.115 4.080 0.425 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.090 1.145 5.180 1.375 ;
        RECT  5.020 0.675 5.090 1.375 ;
        RECT  4.670 1.145 5.020 1.375 ;
        RECT  4.550 1.025 4.670 1.375 ;
        RECT  4.270 1.145 4.550 1.375 ;
        RECT  4.185 0.995 4.270 1.375 ;
        RECT  4.105 1.145 4.185 1.375 ;
        RECT  3.985 0.870 4.105 1.375 ;
        RECT  3.315 1.145 3.985 1.375 ;
        RECT  3.205 0.860 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.635 0.325 4.705 0.915 ;
        RECT  4.165 0.325 4.635 0.395 ;
        RECT  4.280 0.845 4.635 0.915 ;
        RECT  4.375 0.495 4.530 0.765 ;
        RECT  4.210 0.695 4.280 0.915 ;
        RECT  3.685 0.540 4.275 0.610 ;
        RECT  3.910 0.695 4.210 0.765 ;
        RECT  3.710 0.995 3.860 1.075 ;
        RECT  3.675 0.815 3.745 0.885 ;
        RECT  3.465 0.995 3.710 1.065 ;
        RECT  3.675 0.310 3.685 0.610 ;
        RECT  3.605 0.310 3.675 0.885 ;
        RECT  3.465 0.195 3.530 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.375 0.525 4.445 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQD2BWP40

MACRO SDFNCNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.264900 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.745 5.860 1.000 ;
        RECT  5.775 0.205 5.850 0.485 ;
        RECT  5.765 0.205 5.775 1.000 ;
        RECT  5.750 0.355 5.765 1.000 ;
        RECT  5.565 0.355 5.750 0.830 ;
        RECT  5.460 0.355 5.565 0.465 ;
        RECT  5.460 0.710 5.565 0.830 ;
        RECT  5.380 0.195 5.460 0.465 ;
        RECT  5.380 0.710 5.460 1.000 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.050600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.845 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.090 -0.115 6.160 0.115 ;
        RECT  6.020 -0.115 6.090 0.480 ;
        RECT  5.645 -0.115 6.020 0.115 ;
        RECT  5.570 -0.115 5.645 0.275 ;
        RECT  5.280 -0.115 5.570 0.115 ;
        RECT  5.160 -0.115 5.280 0.155 ;
        RECT  4.890 -0.115 5.160 0.115 ;
        RECT  4.755 -0.115 4.890 0.155 ;
        RECT  4.080 -0.115 4.755 0.115 ;
        RECT  4.005 -0.115 4.080 0.425 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.090 1.145 6.160 1.375 ;
        RECT  6.020 0.695 6.090 1.375 ;
        RECT  5.640 1.145 6.020 1.375 ;
        RECT  5.570 0.960 5.640 1.375 ;
        RECT  5.260 1.145 5.570 1.375 ;
        RECT  5.185 1.000 5.260 1.375 ;
        RECT  4.670 1.145 5.185 1.375 ;
        RECT  4.550 1.025 4.670 1.375 ;
        RECT  4.270 1.145 4.550 1.375 ;
        RECT  4.180 0.995 4.270 1.375 ;
        RECT  4.105 1.145 4.180 1.375 ;
        RECT  3.985 0.895 4.105 1.375 ;
        RECT  3.315 1.145 3.985 1.375 ;
        RECT  3.205 1.040 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.845 0.745 5.860 1.000 ;
        RECT  5.845 0.205 5.850 0.485 ;
        RECT  5.460 0.355 5.495 0.465 ;
        RECT  5.460 0.710 5.495 0.830 ;
        RECT  5.380 0.195 5.460 0.465 ;
        RECT  5.380 0.710 5.460 1.000 ;
        RECT  5.310 0.545 5.460 0.615 ;
        RECT  5.235 0.225 5.310 0.925 ;
        RECT  4.360 0.225 5.235 0.295 ;
        RECT  4.280 0.855 5.235 0.925 ;
        RECT  4.260 0.375 5.070 0.445 ;
        RECT  4.845 0.625 5.035 0.765 ;
        RECT  4.670 0.525 4.845 0.765 ;
        RECT  3.685 0.570 4.475 0.640 ;
        RECT  4.210 0.720 4.280 0.925 ;
        RECT  4.190 0.295 4.260 0.445 ;
        RECT  3.910 0.720 4.210 0.790 ;
        RECT  3.710 0.995 3.860 1.075 ;
        RECT  3.675 0.815 3.745 0.885 ;
        RECT  3.465 0.995 3.710 1.065 ;
        RECT  3.675 0.310 3.685 0.640 ;
        RECT  3.605 0.310 3.675 0.885 ;
        RECT  3.465 0.195 3.530 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.725 0.525 4.795 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQD4BWP40

MACRO SDFNCNQND0BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.075 ;
        RECT  4.915 0.185 4.935 0.315 ;
        RECT  4.915 0.910 4.935 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.635 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.790 -0.115 5.040 0.115 ;
        RECT  4.670 -0.115 4.790 0.145 ;
        RECT  4.075 -0.115 4.670 0.115 ;
        RECT  4.005 -0.115 4.075 0.335 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.690 1.025 4.810 1.375 ;
        RECT  4.395 1.145 4.690 1.375 ;
        RECT  4.305 1.005 4.395 1.375 ;
        RECT  4.220 1.145 4.305 1.375 ;
        RECT  4.100 0.985 4.220 1.375 ;
        RECT  3.315 1.145 4.100 1.375 ;
        RECT  3.205 0.815 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.845 0.525 4.850 0.660 ;
        RECT  4.770 0.220 4.845 0.660 ;
        RECT  4.215 0.220 4.770 0.295 ;
        RECT  4.515 0.495 4.670 0.765 ;
        RECT  4.495 0.860 4.600 1.030 ;
        RECT  4.435 0.860 4.495 0.935 ;
        RECT  4.365 0.375 4.435 0.935 ;
        RECT  4.290 0.375 4.365 0.445 ;
        RECT  4.045 0.595 4.365 0.665 ;
        RECT  4.180 0.770 4.280 0.915 ;
        RECT  4.145 0.220 4.215 0.490 ;
        RECT  3.635 0.845 4.180 0.915 ;
        RECT  3.965 0.420 4.145 0.490 ;
        RECT  3.895 0.420 3.965 0.775 ;
        RECT  3.860 0.420 3.895 0.490 ;
        RECT  3.755 0.995 3.875 1.075 ;
        RECT  3.790 0.315 3.860 0.490 ;
        RECT  3.465 0.995 3.755 1.065 ;
        RECT  3.565 0.335 3.635 0.915 ;
        RECT  3.465 0.195 3.530 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.515 0.525 4.585 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQND0BWP40

MACRO SDFNCNQND1BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.075 ;
        RECT  4.915 0.185 4.935 0.465 ;
        RECT  4.915 0.735 4.935 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.038400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.635 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.790 -0.115 5.040 0.115 ;
        RECT  4.670 -0.115 4.790 0.145 ;
        RECT  4.075 -0.115 4.670 0.115 ;
        RECT  4.005 -0.115 4.075 0.335 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.810 1.145 5.040 1.375 ;
        RECT  4.690 0.880 4.810 1.375 ;
        RECT  4.395 1.145 4.690 1.375 ;
        RECT  4.305 1.005 4.395 1.375 ;
        RECT  4.220 1.145 4.305 1.375 ;
        RECT  4.100 0.985 4.220 1.375 ;
        RECT  3.315 1.145 4.100 1.375 ;
        RECT  3.205 0.860 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.845 0.525 4.850 0.660 ;
        RECT  4.770 0.220 4.845 0.660 ;
        RECT  4.215 0.220 4.770 0.295 ;
        RECT  4.515 0.495 4.670 0.765 ;
        RECT  4.435 0.860 4.600 0.935 ;
        RECT  4.365 0.375 4.435 0.935 ;
        RECT  4.290 0.375 4.365 0.445 ;
        RECT  4.045 0.595 4.365 0.665 ;
        RECT  4.180 0.770 4.280 0.915 ;
        RECT  4.145 0.220 4.215 0.490 ;
        RECT  3.635 0.845 4.180 0.915 ;
        RECT  3.965 0.420 4.145 0.490 ;
        RECT  3.895 0.420 3.965 0.775 ;
        RECT  3.860 0.420 3.895 0.490 ;
        RECT  3.755 0.995 3.875 1.075 ;
        RECT  3.790 0.315 3.860 0.490 ;
        RECT  3.475 0.995 3.755 1.065 ;
        RECT  3.565 0.335 3.635 0.915 ;
        RECT  3.475 0.195 3.520 0.265 ;
        RECT  3.385 0.195 3.475 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.515 0.525 4.585 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQND1BWP40

MACRO SDFNCNQND2BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.935 0.185 5.005 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.038400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.635 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.245 -0.115 5.320 0.115 ;
        RECT  5.175 -0.115 5.245 0.490 ;
        RECT  4.790 -0.115 5.175 0.115 ;
        RECT  4.670 -0.115 4.790 0.145 ;
        RECT  4.075 -0.115 4.670 0.115 ;
        RECT  4.005 -0.115 4.075 0.335 ;
        RECT  3.175 -0.115 4.005 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.245 1.145 5.320 1.375 ;
        RECT  5.175 0.670 5.245 1.375 ;
        RECT  4.810 1.145 5.175 1.375 ;
        RECT  4.690 0.880 4.810 1.375 ;
        RECT  4.395 1.145 4.690 1.375 ;
        RECT  4.305 1.005 4.395 1.375 ;
        RECT  4.220 1.145 4.305 1.375 ;
        RECT  4.100 0.985 4.220 1.375 ;
        RECT  3.315 1.145 4.100 1.375 ;
        RECT  3.205 0.860 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.845 0.520 4.850 0.660 ;
        RECT  4.770 0.220 4.845 0.660 ;
        RECT  4.215 0.220 4.770 0.295 ;
        RECT  4.515 0.495 4.670 0.765 ;
        RECT  4.435 0.860 4.600 0.935 ;
        RECT  4.365 0.375 4.435 0.935 ;
        RECT  4.290 0.375 4.365 0.445 ;
        RECT  4.045 0.595 4.365 0.665 ;
        RECT  4.180 0.770 4.280 0.915 ;
        RECT  4.145 0.220 4.215 0.490 ;
        RECT  3.635 0.845 4.180 0.915 ;
        RECT  3.965 0.420 4.145 0.490 ;
        RECT  3.895 0.420 3.965 0.775 ;
        RECT  3.860 0.420 3.895 0.490 ;
        RECT  3.755 0.995 3.875 1.075 ;
        RECT  3.790 0.315 3.860 0.490 ;
        RECT  3.465 0.995 3.755 1.065 ;
        RECT  3.565 0.335 3.635 0.915 ;
        RECT  3.465 0.195 3.525 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.515 0.525 4.585 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQND2BWP40

MACRO SDFNCNQND4BWP40
    CLASS CORE ;
    FOREIGN SDFNCNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.510 0.745 5.620 1.000 ;
        RECT  5.525 0.205 5.610 0.485 ;
        RECT  5.495 0.355 5.525 0.485 ;
        RECT  5.495 0.745 5.510 0.830 ;
        RECT  5.285 0.355 5.495 0.830 ;
        RECT  5.230 0.355 5.285 0.470 ;
        RECT  5.230 0.710 5.285 0.830 ;
        RECT  5.145 0.205 5.230 0.470 ;
        RECT  5.145 0.710 5.230 1.000 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.085 0.640 ;
        RECT  0.945 0.520 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.255 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.039200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.435 0.525 4.915 0.595 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.800 -0.115 5.880 0.115 ;
        RECT  5.730 -0.115 5.800 0.475 ;
        RECT  5.405 -0.115 5.730 0.115 ;
        RECT  5.335 -0.115 5.405 0.275 ;
        RECT  4.990 -0.115 5.335 0.115 ;
        RECT  4.870 -0.115 4.990 0.145 ;
        RECT  4.070 -0.115 4.870 0.115 ;
        RECT  4.000 -0.115 4.070 0.285 ;
        RECT  3.175 -0.115 4.000 0.115 ;
        RECT  3.055 -0.115 3.175 0.235 ;
        RECT  2.750 -0.115 3.055 0.115 ;
        RECT  2.620 -0.115 2.750 0.235 ;
        RECT  1.565 -0.115 2.620 0.115 ;
        RECT  1.440 -0.115 1.565 0.120 ;
        RECT  1.180 -0.115 1.440 0.115 ;
        RECT  1.060 -0.115 1.180 0.125 ;
        RECT  0.340 -0.115 1.060 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.800 1.145 5.880 1.375 ;
        RECT  5.730 0.705 5.800 1.375 ;
        RECT  5.405 1.145 5.730 1.375 ;
        RECT  5.335 0.915 5.405 1.375 ;
        RECT  5.010 1.145 5.335 1.375 ;
        RECT  4.930 0.835 5.010 1.375 ;
        RECT  4.595 1.145 4.930 1.375 ;
        RECT  4.505 1.095 4.595 1.375 ;
        RECT  4.190 1.145 4.505 1.375 ;
        RECT  4.060 1.035 4.190 1.375 ;
        RECT  3.315 1.145 4.060 1.375 ;
        RECT  3.205 0.860 3.315 1.375 ;
        RECT  2.620 1.145 3.205 1.375 ;
        RECT  2.500 1.070 2.620 1.375 ;
        RECT  1.460 1.145 2.500 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.565 0.745 5.620 1.000 ;
        RECT  5.565 0.205 5.610 0.485 ;
        RECT  5.145 0.205 5.215 0.470 ;
        RECT  5.145 0.710 5.215 1.000 ;
        RECT  5.055 0.545 5.185 0.615 ;
        RECT  4.985 0.220 5.055 0.615 ;
        RECT  4.300 0.220 4.985 0.295 ;
        RECT  4.715 0.495 4.870 0.765 ;
        RECT  4.635 0.925 4.800 1.000 ;
        RECT  4.565 0.375 4.635 1.000 ;
        RECT  4.490 0.375 4.565 0.445 ;
        RECT  4.110 0.545 4.565 0.615 ;
        RECT  4.390 0.855 4.465 1.005 ;
        RECT  4.020 0.855 4.390 0.925 ;
        RECT  3.950 0.705 4.385 0.775 ;
        RECT  4.230 0.220 4.300 0.425 ;
        RECT  3.950 0.355 4.230 0.425 ;
        RECT  3.950 0.845 4.020 0.925 ;
        RECT  3.880 0.355 3.950 0.775 ;
        RECT  3.630 0.845 3.950 0.915 ;
        RECT  3.760 0.355 3.880 0.425 ;
        RECT  3.745 0.995 3.870 1.075 ;
        RECT  3.465 0.995 3.745 1.065 ;
        RECT  3.560 0.335 3.630 0.915 ;
        RECT  3.465 0.195 3.525 0.265 ;
        RECT  3.385 0.195 3.465 1.065 ;
        RECT  3.040 0.335 3.110 0.860 ;
        RECT  2.860 0.335 3.040 0.405 ;
        RECT  2.475 0.790 3.040 0.860 ;
        RECT  2.760 0.510 2.900 0.580 ;
        RECT  2.315 0.930 2.810 1.000 ;
        RECT  2.690 0.335 2.760 0.580 ;
        RECT  2.540 0.335 2.690 0.405 ;
        RECT  2.545 0.475 2.620 0.710 ;
        RECT  2.405 0.475 2.545 0.610 ;
        RECT  2.470 0.195 2.540 0.405 ;
        RECT  2.385 0.680 2.475 0.860 ;
        RECT  2.130 0.195 2.470 0.265 ;
        RECT  2.315 0.360 2.335 0.480 ;
        RECT  2.245 0.360 2.315 1.000 ;
        RECT  2.105 0.520 2.175 0.920 ;
        RECT  2.060 0.195 2.130 0.405 ;
        RECT  1.470 0.850 2.105 0.920 ;
        RECT  2.035 0.335 2.060 0.405 ;
        RECT  1.965 0.335 2.035 0.780 ;
        RECT  1.945 0.690 1.965 0.780 ;
        RECT  0.640 0.195 1.940 0.265 ;
        RECT  0.715 0.990 1.880 1.060 ;
        RECT  1.695 0.350 1.765 0.780 ;
        RECT  1.590 0.350 1.695 0.420 ;
        RECT  1.560 0.710 1.695 0.780 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.920 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.850 1.400 0.920 ;
        RECT  0.865 0.335 0.945 0.445 ;
        RECT  0.865 0.835 0.940 0.905 ;
        RECT  0.795 0.335 0.865 0.905 ;
        RECT  0.645 0.810 0.715 1.060 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.795 0.525 4.865 0.595 ;
        RECT  2.485 0.525 2.555 0.595 ;
    END
END SDFNCNQND4BWP40

MACRO SDFNCSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFNCSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.215 5.565 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.390 -0.115 5.600 0.115 ;
        RECT  5.255 -0.115 5.390 0.350 ;
        RECT  4.360 -0.115 5.255 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.260 ;
        RECT  1.190 -0.115 3.455 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.380 1.145 5.600 1.375 ;
        RECT  5.260 0.940 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  4.945 0.930 5.075 1.000 ;
        RECT  4.785 0.510 5.005 0.630 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.865 0.705 4.945 1.000 ;
        RECT  3.920 0.930 4.865 1.000 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.790 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.365 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.715 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  0.640 0.195 1.900 0.265 ;
        RECT  1.720 0.530 1.855 0.600 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.345 1.720 0.790 ;
        RECT  1.590 0.345 1.650 0.415 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNCSNQD0BWP40

MACRO SDFNCSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFNCSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.205 5.565 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.033600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 -0.115 5.600 0.115 ;
        RECT  5.270 -0.115 5.365 0.310 ;
        RECT  4.360 -0.115 5.270 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.260 ;
        RECT  1.190 -0.115 3.455 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.380 1.145 5.600 1.375 ;
        RECT  5.260 0.870 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  3.920 0.930 5.075 1.000 ;
        RECT  4.785 0.460 5.005 0.580 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.715 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  1.800 0.195 1.880 0.420 ;
        RECT  1.720 0.515 1.855 0.585 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  0.640 0.195 1.800 0.265 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.345 1.720 0.790 ;
        RECT  1.590 0.345 1.650 0.415 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNCSNQD1BWP40

MACRO SDFNCSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFNCSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.450 5.320 0.765 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.033600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.235 0.490 4.465 0.675 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 -0.115 5.880 0.115 ;
        RECT  5.740 -0.115 5.810 0.485 ;
        RECT  5.390 -0.115 5.740 0.115 ;
        RECT  5.255 -0.115 5.390 0.310 ;
        RECT  4.360 -0.115 5.255 0.115 ;
        RECT  4.225 -0.115 4.360 0.250 ;
        RECT  3.525 -0.115 4.225 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.190 -0.115 3.455 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 1.145 5.880 1.375 ;
        RECT  5.740 0.690 5.810 1.375 ;
        RECT  5.380 1.145 5.740 1.375 ;
        RECT  5.260 0.865 5.380 1.375 ;
        RECT  4.975 1.145 5.260 1.375 ;
        RECT  4.845 1.095 4.975 1.375 ;
        RECT  4.370 1.145 4.845 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.075 0.285 5.145 1.000 ;
        RECT  3.920 0.930 5.075 1.000 ;
        RECT  4.785 0.460 5.005 0.580 ;
        RECT  4.460 0.195 4.975 0.265 ;
        RECT  4.710 0.335 4.785 0.860 ;
        RECT  4.675 0.335 4.710 0.445 ;
        RECT  4.450 0.790 4.710 0.860 ;
        RECT  4.605 0.520 4.630 0.700 ;
        RECT  4.535 0.340 4.605 0.700 ;
        RECT  4.030 0.340 4.535 0.410 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.960 0.195 4.030 0.410 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.685 0.195 3.960 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.720 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  1.800 0.195 1.880 0.420 ;
        RECT  1.720 0.515 1.855 0.585 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  0.640 0.195 1.800 0.265 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.345 1.720 0.790 ;
        RECT  1.590 0.345 1.650 0.415 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNCSNQD2BWP40

MACRO SDFNCSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFNCSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.026800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.775 0.450 5.870 0.765 ;
        RECT  5.765 0.525 5.775 0.635 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.405 0.195 6.500 0.485 ;
        RECT  6.405 0.710 6.500 0.995 ;
        RECT  6.335 0.355 6.405 0.485 ;
        RECT  6.335 0.710 6.405 0.830 ;
        RECT  6.125 0.355 6.335 0.830 ;
        RECT  6.100 0.355 6.125 0.485 ;
        RECT  6.100 0.710 6.125 0.830 ;
        RECT  6.025 0.215 6.100 0.485 ;
        RECT  6.025 0.710 6.100 0.980 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.495 1.085 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.044600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.315 0.355 4.445 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 -0.115 6.720 0.115 ;
        RECT  6.595 -0.115 6.665 0.440 ;
        RECT  6.290 -0.115 6.595 0.115 ;
        RECT  6.205 -0.115 6.290 0.265 ;
        RECT  5.920 -0.115 6.205 0.115 ;
        RECT  5.830 -0.115 5.920 0.310 ;
        RECT  5.170 -0.115 5.830 0.115 ;
        RECT  5.050 -0.115 5.170 0.140 ;
        RECT  4.370 -0.115 5.050 0.115 ;
        RECT  4.235 -0.115 4.370 0.130 ;
        RECT  3.525 -0.115 4.235 0.115 ;
        RECT  3.455 -0.115 3.525 0.400 ;
        RECT  1.190 -0.115 3.455 0.115 ;
        RECT  1.070 -0.115 1.190 0.125 ;
        RECT  0.340 -0.115 1.070 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.665 1.145 6.720 1.375 ;
        RECT  6.595 0.680 6.665 1.375 ;
        RECT  6.310 1.145 6.595 1.375 ;
        RECT  6.190 0.910 6.310 1.375 ;
        RECT  5.910 1.145 6.190 1.375 ;
        RECT  5.835 0.860 5.910 1.375 ;
        RECT  5.000 1.145 5.835 1.375 ;
        RECT  4.880 1.070 5.000 1.375 ;
        RECT  4.370 1.145 4.880 1.375 ;
        RECT  4.250 1.070 4.370 1.375 ;
        RECT  2.670 1.145 4.250 1.375 ;
        RECT  2.510 1.130 2.670 1.375 ;
        RECT  1.460 1.145 2.510 1.375 ;
        RECT  1.330 1.130 1.460 1.375 ;
        RECT  1.150 1.145 1.330 1.375 ;
        RECT  1.030 1.130 1.150 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.405 0.195 6.500 0.485 ;
        RECT  6.405 0.710 6.500 0.995 ;
        RECT  6.025 0.215 6.055 0.485 ;
        RECT  6.025 0.710 6.055 0.980 ;
        RECT  5.625 0.210 5.695 1.000 ;
        RECT  5.045 0.930 5.625 1.000 ;
        RECT  5.515 0.620 5.555 0.740 ;
        RECT  5.445 0.210 5.515 0.860 ;
        RECT  4.765 0.210 5.445 0.280 ;
        RECT  5.330 0.790 5.445 0.860 ;
        RECT  4.845 0.350 5.350 0.420 ;
        RECT  4.965 0.605 5.045 1.000 ;
        RECT  3.920 0.930 4.965 1.000 ;
        RECT  4.695 0.210 4.765 0.860 ;
        RECT  4.690 0.335 4.695 0.860 ;
        RECT  4.675 0.335 4.690 0.445 ;
        RECT  4.205 0.790 4.690 0.860 ;
        RECT  4.585 0.580 4.620 0.700 ;
        RECT  4.515 0.200 4.585 0.700 ;
        RECT  3.980 0.200 4.515 0.270 ;
        RECT  4.135 0.445 4.205 0.860 ;
        RECT  3.990 0.535 4.065 0.785 ;
        RECT  3.880 0.535 3.990 0.605 ;
        RECT  3.935 0.195 3.980 0.270 ;
        RECT  3.685 0.195 3.935 0.265 ;
        RECT  3.845 0.825 3.920 1.000 ;
        RECT  3.685 0.685 3.910 0.755 ;
        RECT  3.765 0.355 3.880 0.605 ;
        RECT  3.455 0.825 3.845 0.900 ;
        RECT  3.600 0.970 3.755 1.060 ;
        RECT  3.615 0.195 3.685 0.755 ;
        RECT  2.025 0.990 3.600 1.060 ;
        RECT  3.385 0.825 3.455 0.915 ;
        RECT  3.385 0.485 3.395 0.625 ;
        RECT  3.315 0.205 3.385 0.625 ;
        RECT  3.025 0.840 3.385 0.915 ;
        RECT  2.090 0.205 3.315 0.275 ;
        RECT  3.185 0.355 3.245 0.575 ;
        RECT  3.165 0.355 3.185 0.760 ;
        RECT  3.095 0.505 3.165 0.760 ;
        RECT  2.370 0.505 3.095 0.575 ;
        RECT  2.955 0.645 3.025 0.915 ;
        RECT  2.650 0.645 2.955 0.715 ;
        RECT  2.405 0.355 2.900 0.425 ;
        RECT  2.800 0.800 2.875 0.920 ;
        RECT  2.230 0.850 2.800 0.920 ;
        RECT  2.555 0.645 2.650 0.770 ;
        RECT  2.300 0.505 2.370 0.715 ;
        RECT  2.230 0.355 2.305 0.425 ;
        RECT  2.160 0.355 2.230 0.920 ;
        RECT  2.045 0.205 2.090 0.580 ;
        RECT  2.015 0.205 2.045 0.915 ;
        RECT  1.935 0.510 2.015 0.915 ;
        RECT  1.800 0.195 1.880 0.420 ;
        RECT  1.720 0.515 1.855 0.585 ;
        RECT  1.760 0.860 1.830 1.055 ;
        RECT  0.640 0.195 1.800 0.265 ;
        RECT  0.715 0.985 1.760 1.055 ;
        RECT  1.650 0.345 1.720 0.790 ;
        RECT  1.590 0.345 1.650 0.415 ;
        RECT  1.560 0.720 1.650 0.790 ;
        RECT  1.470 0.520 1.580 0.640 ;
        RECT  1.400 0.345 1.470 0.915 ;
        RECT  1.220 0.345 1.400 0.415 ;
        RECT  1.170 0.845 1.400 0.915 ;
        RECT  0.870 0.350 0.990 0.420 ;
        RECT  0.870 0.845 0.940 0.915 ;
        RECT  0.800 0.350 0.870 0.915 ;
        RECT  0.645 0.790 0.715 1.055 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.190 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNCSNQD4BWP40

MACRO SDFNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.045 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.625 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.060 -0.115 1.920 0.115 ;
        RECT  0.940 -0.115 1.060 0.125 ;
        RECT  0.340 -0.115 0.940 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.810 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.740 3.785 0.810 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.980 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  1.680 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQD0BWP40

MACRO SDFNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.625 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.045 -0.115 1.920 0.115 ;
        RECT  0.925 -0.115 1.045 0.125 ;
        RECT  0.340 -0.115 0.925 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.765 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.695 3.785 0.765 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  2.415 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  2.330 0.195 2.415 0.345 ;
        RECT  1.680 0.195 2.330 0.265 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQD1BWP40

MACRO SDFNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.050 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.625 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.275 -0.115 4.340 0.115 ;
        RECT  4.190 -0.115 4.275 0.450 ;
        RECT  3.815 -0.115 4.190 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.045 -0.115 1.920 0.115 ;
        RECT  0.925 -0.115 1.045 0.125 ;
        RECT  0.340 -0.115 0.925 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 1.145 4.340 1.375 ;
        RECT  4.190 0.710 4.270 1.375 ;
        RECT  3.815 1.145 4.190 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.765 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.695 3.785 0.765 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  2.420 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  2.330 0.195 2.420 0.345 ;
        RECT  1.680 0.195 2.330 0.265 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQD2BWP40

MACRO SDFNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.210 4.405 0.455 ;
        RECT  4.305 0.735 4.405 1.030 ;
        RECT  4.235 0.370 4.305 0.455 ;
        RECT  4.235 0.735 4.305 0.820 ;
        RECT  4.025 0.370 4.235 0.820 ;
        RECT  4.000 0.370 4.025 0.455 ;
        RECT  4.005 0.735 4.025 0.820 ;
        RECT  3.920 0.735 4.005 1.045 ;
        RECT  3.920 0.185 4.000 0.455 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.355 2.520 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.565 -0.115 4.620 0.115 ;
        RECT  4.495 -0.115 4.565 0.420 ;
        RECT  4.190 -0.115 4.495 0.115 ;
        RECT  4.115 -0.115 4.190 0.250 ;
        RECT  3.805 -0.115 4.115 0.115 ;
        RECT  3.735 -0.115 3.805 0.315 ;
        RECT  3.415 -0.115 3.735 0.115 ;
        RECT  3.345 -0.115 3.415 0.315 ;
        RECT  2.620 -0.115 3.345 0.115 ;
        RECT  2.500 -0.115 2.620 0.130 ;
        RECT  2.040 -0.115 2.500 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.040 -0.115 1.920 0.115 ;
        RECT  0.920 -0.115 1.040 0.125 ;
        RECT  0.340 -0.115 0.920 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.560 1.145 4.620 1.375 ;
        RECT  4.485 0.685 4.560 1.375 ;
        RECT  4.210 1.145 4.485 1.375 ;
        RECT  4.090 0.905 4.210 1.375 ;
        RECT  3.805 1.145 4.090 1.375 ;
        RECT  3.735 0.845 3.805 1.375 ;
        RECT  3.420 1.145 3.735 1.375 ;
        RECT  3.290 1.130 3.420 1.375 ;
        RECT  2.620 1.145 3.290 1.375 ;
        RECT  2.500 1.040 2.620 1.375 ;
        RECT  2.050 1.145 2.500 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.210 4.405 0.455 ;
        RECT  4.305 0.735 4.405 1.030 ;
        RECT  3.920 0.185 3.955 0.455 ;
        RECT  3.920 0.735 3.955 1.045 ;
        RECT  3.835 0.545 3.950 0.615 ;
        RECT  3.765 0.395 3.835 0.765 ;
        RECT  3.615 0.395 3.765 0.465 ;
        RECT  3.615 0.695 3.765 0.765 ;
        RECT  3.475 0.545 3.640 0.615 ;
        RECT  3.545 0.185 3.615 0.465 ;
        RECT  3.545 0.695 3.615 1.025 ;
        RECT  3.315 0.395 3.545 0.465 ;
        RECT  3.395 0.545 3.475 0.930 ;
        RECT  3.000 0.860 3.395 0.930 ;
        RECT  3.245 0.395 3.315 0.600 ;
        RECT  3.095 0.195 3.175 0.780 ;
        RECT  2.850 0.195 3.095 0.265 ;
        RECT  2.930 0.350 3.000 0.930 ;
        RECT  2.780 0.195 2.850 0.915 ;
        RECT  2.430 0.200 2.780 0.270 ;
        RECT  2.310 0.845 2.780 0.915 ;
        RECT  2.605 0.425 2.675 0.745 ;
        RECT  2.275 0.195 2.430 0.270 ;
        RECT  2.145 0.475 2.310 0.545 ;
        RECT  1.680 0.195 2.275 0.265 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.360 0.845 1.530 0.915 ;
        RECT  0.585 0.195 1.460 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.360 0.345 1.415 0.505 ;
        RECT  1.290 0.345 1.360 0.915 ;
        RECT  1.150 0.345 1.290 0.415 ;
        RECT  1.145 0.845 1.290 0.915 ;
        RECT  0.805 0.845 0.910 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.535 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.535 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.605 0.525 2.675 0.595 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.725 0.595 ;
    END
END SDFNQD4BWP40

MACRO SDFNQND0BWP40
    CLASS CORE ;
    FOREIGN SDFNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.045 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.615 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.045 -0.115 1.920 0.115 ;
        RECT  0.925 -0.115 1.045 0.125 ;
        RECT  0.340 -0.115 0.925 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.810 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.740 3.785 0.810 ;
        RECT  3.485 0.545 3.680 0.615 ;
        RECT  3.565 0.330 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.980 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  1.680 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQND0BWP40

MACRO SDFNQND1BWP40
    CLASS CORE ;
    FOREIGN SDFNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.625 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.060 -0.115 1.920 0.115 ;
        RECT  0.940 -0.115 1.060 0.125 ;
        RECT  0.340 -0.115 0.940 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.765 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.695 3.785 0.765 ;
        RECT  3.485 0.545 3.690 0.615 ;
        RECT  3.565 0.330 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  1.680 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQND1BWP40

MACRO SDFNQND2BWP40
    CLASS CORE ;
    FOREIGN SDFNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.040 1.065 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.625 2.635 0.765 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.275 -0.115 4.340 0.115 ;
        RECT  4.190 -0.115 4.275 0.450 ;
        RECT  3.815 -0.115 4.190 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.650 -0.115 3.375 0.115 ;
        RECT  2.530 -0.115 2.650 0.125 ;
        RECT  2.040 -0.115 2.530 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.060 -0.115 1.920 0.115 ;
        RECT  0.940 -0.115 1.060 0.125 ;
        RECT  0.340 -0.115 0.940 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 1.145 4.340 1.375 ;
        RECT  4.190 0.765 4.270 1.375 ;
        RECT  3.815 1.145 4.190 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 1.030 2.630 1.375 ;
        RECT  2.050 1.145 2.510 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.705 0.395 3.775 0.765 ;
        RECT  3.635 0.395 3.705 0.465 ;
        RECT  3.635 0.695 3.705 0.765 ;
        RECT  3.565 0.330 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.870 0.195 3.110 0.265 ;
        RECT  2.950 0.340 3.020 0.930 ;
        RECT  2.800 0.195 2.870 0.930 ;
        RECT  1.680 0.195 2.800 0.265 ;
        RECT  2.315 0.860 2.800 0.930 ;
        RECT  2.145 0.475 2.720 0.545 ;
        RECT  1.990 0.335 2.245 0.405 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.475 2.145 0.635 ;
        RECT  1.920 0.335 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQND2BWP40

MACRO SDFNQND4BWP40
    CLASS CORE ;
    FOREIGN SDFNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.195 4.820 0.440 ;
        RECT  4.725 0.705 4.820 1.010 ;
        RECT  4.655 0.355 4.725 0.440 ;
        RECT  4.655 0.705 4.725 0.805 ;
        RECT  4.445 0.355 4.655 0.805 ;
        RECT  4.415 0.355 4.445 0.485 ;
        RECT  4.420 0.710 4.445 0.805 ;
        RECT  4.345 0.710 4.420 0.970 ;
        RECT  4.345 0.210 4.415 0.485 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.018800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.100 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.540 0.495 2.905 0.630 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.990 0.465 ;
        RECT  4.630 -0.115 4.915 0.115 ;
        RECT  4.510 -0.115 4.630 0.225 ;
        RECT  4.225 -0.115 4.510 0.115 ;
        RECT  4.155 -0.115 4.225 0.315 ;
        RECT  3.860 -0.115 4.155 0.115 ;
        RECT  3.790 -0.115 3.860 0.315 ;
        RECT  2.785 -0.115 3.790 0.115 ;
        RECT  2.665 -0.115 2.785 0.125 ;
        RECT  2.430 -0.115 2.665 0.115 ;
        RECT  2.310 -0.115 2.430 0.130 ;
        RECT  2.040 -0.115 2.310 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.060 -0.115 1.920 0.115 ;
        RECT  0.940 -0.115 1.060 0.125 ;
        RECT  0.340 -0.115 0.940 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.990 1.145 5.040 1.375 ;
        RECT  4.915 0.710 4.990 1.375 ;
        RECT  4.630 1.145 4.915 1.375 ;
        RECT  4.510 0.875 4.630 1.375 ;
        RECT  4.225 1.145 4.510 1.375 ;
        RECT  4.155 0.845 4.225 1.375 ;
        RECT  3.860 1.145 4.155 1.375 ;
        RECT  3.730 1.130 3.860 1.375 ;
        RECT  2.835 1.145 3.730 1.375 ;
        RECT  2.715 1.025 2.835 1.375 ;
        RECT  2.405 1.145 2.715 1.375 ;
        RECT  2.335 0.995 2.405 1.375 ;
        RECT  2.050 1.145 2.335 1.375 ;
        RECT  1.930 0.900 2.050 1.375 ;
        RECT  1.120 1.145 1.930 1.375 ;
        RECT  1.000 1.130 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.195 4.820 0.440 ;
        RECT  4.725 0.705 4.820 1.010 ;
        RECT  4.345 0.210 4.375 0.485 ;
        RECT  4.345 0.710 4.375 0.970 ;
        RECT  4.195 0.395 4.265 0.765 ;
        RECT  4.045 0.395 4.195 0.465 ;
        RECT  4.050 0.695 4.195 0.765 ;
        RECT  3.900 0.545 4.070 0.615 ;
        RECT  3.980 0.695 4.050 0.980 ;
        RECT  3.975 0.330 4.045 0.465 ;
        RECT  3.750 0.395 3.975 0.465 ;
        RECT  3.830 0.545 3.900 0.930 ;
        RECT  3.425 0.860 3.830 0.930 ;
        RECT  3.680 0.395 3.750 0.600 ;
        RECT  3.530 0.200 3.605 0.780 ;
        RECT  3.285 0.200 3.530 0.270 ;
        RECT  3.355 0.350 3.425 0.930 ;
        RECT  3.215 0.200 3.285 0.625 ;
        RECT  2.500 0.885 3.245 0.955 ;
        RECT  2.260 0.200 3.215 0.270 ;
        RECT  3.060 0.555 3.215 0.625 ;
        RECT  3.070 0.355 3.145 0.475 ;
        RECT  2.500 0.355 3.070 0.425 ;
        RECT  2.990 0.555 3.060 0.805 ;
        RECT  2.910 0.735 2.990 0.805 ;
        RECT  2.145 0.480 2.305 0.550 ;
        RECT  2.175 0.195 2.260 0.270 ;
        RECT  1.990 0.340 2.250 0.410 ;
        RECT  2.150 0.745 2.225 0.950 ;
        RECT  1.680 0.195 2.175 0.265 ;
        RECT  1.990 0.745 2.150 0.815 ;
        RECT  2.075 0.480 2.145 0.660 ;
        RECT  1.920 0.340 1.990 0.815 ;
        RECT  1.900 0.620 1.920 0.740 ;
        RECT  1.795 0.345 1.850 0.570 ;
        RECT  1.795 0.810 1.825 0.915 ;
        RECT  1.770 0.345 1.795 0.915 ;
        RECT  1.725 0.500 1.770 0.915 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.655 0.355 1.690 0.435 ;
        RECT  1.575 0.355 1.655 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.690 1.575 0.760 ;
        RECT  1.450 0.845 1.530 0.915 ;
        RECT  1.450 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.470 0.265 ;
        RECT  1.360 0.345 1.450 0.915 ;
        RECT  0.585 0.985 1.450 1.055 ;
        RECT  1.150 0.345 1.360 0.415 ;
        RECT  1.145 0.845 1.360 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.610 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.075 0.525 2.145 0.595 ;
        RECT  1.585 0.525 1.655 0.595 ;
        LAYER M2 ;
        RECT  1.535 0.525 2.195 0.595 ;
    END
END SDFNQND4BWP40

MACRO SDFNSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.315 4.725 0.925 ;
        RECT  4.635 0.315 4.655 0.435 ;
        RECT  4.635 0.795 4.655 0.925 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.610 2.835 0.680 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.115 4.760 0.115 ;
        RECT  4.440 -0.115 4.520 0.425 ;
        RECT  4.125 -0.115 4.440 0.115 ;
        RECT  4.055 -0.115 4.125 0.280 ;
        RECT  3.740 -0.115 4.055 0.115 ;
        RECT  3.620 -0.115 3.740 0.280 ;
        RECT  2.805 -0.115 3.620 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.760 1.375 ;
        RECT  4.420 1.080 4.540 1.375 ;
        RECT  3.740 1.145 4.420 1.375 ;
        RECT  3.620 0.860 3.740 1.375 ;
        RECT  2.900 1.145 3.620 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.115 1.145 2.395 1.375 ;
        RECT  1.995 1.050 2.115 1.375 ;
        RECT  1.125 1.145 1.995 1.375 ;
        RECT  0.995 1.120 1.125 1.375 ;
        RECT  0.340 1.145 0.995 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.525 4.585 0.635 ;
        RECT  4.490 0.525 4.565 1.010 ;
        RECT  4.120 0.940 4.490 1.010 ;
        RECT  4.255 0.325 4.325 0.870 ;
        RECT  4.190 0.580 4.255 0.700 ;
        RECT  4.050 0.350 4.120 1.010 ;
        RECT  3.590 0.350 4.050 0.420 ;
        RECT  3.910 0.615 3.980 0.780 ;
        RECT  3.325 0.710 3.910 0.780 ;
        RECT  3.520 0.350 3.590 0.610 ;
        RECT  3.350 0.995 3.460 1.075 ;
        RECT  3.135 0.995 3.350 1.065 ;
        RECT  3.285 0.710 3.325 0.925 ;
        RECT  3.215 0.335 3.285 0.925 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.685 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.775 2.685 0.980 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.980 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  1.820 0.910 2.555 0.980 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.830 ;
        RECT  1.750 0.910 1.820 1.065 ;
        RECT  1.750 0.760 1.795 0.830 ;
        RECT  1.610 0.995 1.750 1.065 ;
        RECT  1.605 0.195 1.675 0.910 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.565 0.840 1.605 0.910 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.350 0.960 0.420 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.350 0.865 0.910 ;
        RECT  0.645 0.875 0.715 1.050 ;
        RECT  0.555 0.530 0.610 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQD0BWP40

MACRO SDFNSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.075 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.685 4.655 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.115 4.760 0.115 ;
        RECT  4.440 -0.115 4.520 0.420 ;
        RECT  4.125 -0.115 4.440 0.115 ;
        RECT  4.055 -0.115 4.125 0.280 ;
        RECT  3.740 -0.115 4.055 0.115 ;
        RECT  3.620 -0.115 3.740 0.280 ;
        RECT  2.805 -0.115 3.620 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.760 1.375 ;
        RECT  4.420 1.080 4.540 1.375 ;
        RECT  3.740 1.145 4.420 1.375 ;
        RECT  3.620 0.860 3.740 1.375 ;
        RECT  2.900 1.145 3.620 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.115 1.145 2.395 1.375 ;
        RECT  1.995 1.050 2.115 1.375 ;
        RECT  1.120 1.145 1.995 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.525 4.585 0.635 ;
        RECT  4.490 0.525 4.565 1.010 ;
        RECT  4.120 0.940 4.490 1.010 ;
        RECT  4.255 0.370 4.325 0.870 ;
        RECT  4.190 0.580 4.255 0.700 ;
        RECT  4.050 0.350 4.120 1.010 ;
        RECT  3.590 0.350 4.050 0.420 ;
        RECT  3.910 0.615 3.980 0.780 ;
        RECT  3.325 0.710 3.910 0.780 ;
        RECT  3.520 0.350 3.590 0.610 ;
        RECT  3.350 0.995 3.460 1.075 ;
        RECT  3.135 0.995 3.350 1.065 ;
        RECT  3.285 0.710 3.325 0.925 ;
        RECT  3.215 0.335 3.285 0.925 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.685 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.775 2.685 0.980 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.980 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  1.820 0.910 2.555 0.980 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.830 ;
        RECT  1.750 0.910 1.820 1.065 ;
        RECT  1.750 0.760 1.795 0.830 ;
        RECT  1.610 0.995 1.750 1.065 ;
        RECT  1.605 0.195 1.675 0.910 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.565 0.840 1.605 0.910 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQD1BWP40

MACRO SDFNSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.660 0.370 4.725 0.880 ;
        RECT  4.655 0.195 4.660 1.075 ;
        RECT  4.585 0.195 4.655 0.445 ;
        RECT  4.585 0.805 4.655 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.680 0.605 2.835 0.675 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.255 ;
        RECT  4.470 -0.115 4.775 0.115 ;
        RECT  4.395 -0.115 4.470 0.420 ;
        RECT  4.070 -0.115 4.395 0.115 ;
        RECT  3.980 -0.115 4.070 0.280 ;
        RECT  3.700 -0.115 3.980 0.115 ;
        RECT  3.570 -0.115 3.700 0.280 ;
        RECT  2.780 -0.115 3.570 0.115 ;
        RECT  2.660 -0.115 2.780 0.190 ;
        RECT  2.065 -0.115 2.660 0.115 ;
        RECT  1.935 -0.115 2.065 0.125 ;
        RECT  1.145 -0.115 1.935 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.950 4.845 1.375 ;
        RECT  4.490 1.145 4.775 1.375 ;
        RECT  4.370 1.080 4.490 1.375 ;
        RECT  3.705 1.145 4.370 1.375 ;
        RECT  3.635 0.995 3.705 1.375 ;
        RECT  2.875 1.145 3.635 1.375 ;
        RECT  2.745 1.050 2.875 1.375 ;
        RECT  2.485 1.145 2.745 1.375 ;
        RECT  2.355 1.050 2.485 1.375 ;
        RECT  2.220 1.145 2.355 1.375 ;
        RECT  2.090 1.070 2.220 1.375 ;
        RECT  1.120 1.145 2.090 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.515 0.525 4.585 0.635 ;
        RECT  4.440 0.525 4.515 0.985 ;
        RECT  4.070 0.915 4.440 0.985 ;
        RECT  4.210 0.330 4.300 0.405 ;
        RECT  4.210 0.775 4.300 0.845 ;
        RECT  4.140 0.330 4.210 0.845 ;
        RECT  4.000 0.350 4.070 0.985 ;
        RECT  3.575 0.350 4.000 0.420 ;
        RECT  3.860 0.500 3.930 0.915 ;
        RECT  3.265 0.845 3.860 0.915 ;
        RECT  3.505 0.350 3.575 0.610 ;
        RECT  3.340 0.995 3.450 1.075 ;
        RECT  3.115 0.995 3.340 1.065 ;
        RECT  3.195 0.335 3.265 0.915 ;
        RECT  3.115 0.195 3.175 0.265 ;
        RECT  3.045 0.195 3.115 1.065 ;
        RECT  3.020 0.870 3.045 1.065 ;
        RECT  2.590 0.870 3.020 0.940 ;
        RECT  2.855 0.185 2.965 0.330 ;
        RECT  2.590 0.260 2.855 0.330 ;
        RECT  2.590 0.410 2.690 0.480 ;
        RECT  2.520 0.195 2.590 0.330 ;
        RECT  2.520 0.410 2.590 0.940 ;
        RECT  1.670 0.195 2.520 0.265 ;
        RECT  2.020 0.870 2.520 0.940 ;
        RECT  2.370 0.345 2.440 0.765 ;
        RECT  1.985 0.695 2.370 0.765 ;
        RECT  1.950 0.870 2.020 1.065 ;
        RECT  1.915 0.575 1.985 0.765 ;
        RECT  1.610 0.995 1.950 1.065 ;
        RECT  1.820 0.335 1.890 0.405 ;
        RECT  1.820 0.830 1.870 0.900 ;
        RECT  1.750 0.335 1.820 0.900 ;
        RECT  1.600 0.195 1.670 0.925 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.585 0.815 1.600 0.925 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQD2BWP40

MACRO SDFNSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.185 5.380 0.460 ;
        RECT  5.285 0.785 5.370 1.075 ;
        RECT  5.215 0.330 5.285 0.460 ;
        RECT  5.215 0.785 5.285 0.905 ;
        RECT  5.005 0.330 5.215 0.905 ;
        RECT  4.995 0.330 5.005 0.460 ;
        RECT  4.995 0.785 5.005 0.905 ;
        RECT  4.905 0.185 4.995 0.460 ;
        RECT  4.905 0.785 4.995 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.495 2.905 0.765 ;
        RECT  2.830 0.495 2.835 0.680 ;
        RECT  2.670 0.610 2.830 0.680 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 -0.115 5.600 0.115 ;
        RECT  5.475 -0.115 5.545 0.410 ;
        RECT  5.165 -0.115 5.475 0.115 ;
        RECT  5.095 -0.115 5.165 0.255 ;
        RECT  4.790 -0.115 5.095 0.115 ;
        RECT  4.715 -0.115 4.790 0.420 ;
        RECT  4.055 -0.115 4.715 0.115 ;
        RECT  3.925 -0.115 4.055 0.250 ;
        RECT  3.670 -0.115 3.925 0.115 ;
        RECT  3.540 -0.115 3.670 0.250 ;
        RECT  2.770 -0.115 3.540 0.115 ;
        RECT  2.650 -0.115 2.770 0.190 ;
        RECT  2.065 -0.115 2.650 0.115 ;
        RECT  1.935 -0.115 2.065 0.125 ;
        RECT  1.145 -0.115 1.935 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 1.145 5.600 1.375 ;
        RECT  5.475 0.725 5.545 1.375 ;
        RECT  5.165 1.145 5.475 1.375 ;
        RECT  5.095 0.995 5.165 1.375 ;
        RECT  4.820 1.145 5.095 1.375 ;
        RECT  4.690 1.030 4.820 1.375 ;
        RECT  4.445 1.145 4.690 1.375 ;
        RECT  4.310 1.030 4.445 1.375 ;
        RECT  3.675 1.145 4.310 1.375 ;
        RECT  3.605 0.995 3.675 1.375 ;
        RECT  2.865 1.145 3.605 1.375 ;
        RECT  2.735 1.050 2.865 1.375 ;
        RECT  2.480 1.145 2.735 1.375 ;
        RECT  2.355 1.050 2.480 1.375 ;
        RECT  2.220 1.145 2.355 1.375 ;
        RECT  2.090 1.070 2.220 1.375 ;
        RECT  1.120 1.145 2.090 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.185 5.380 0.460 ;
        RECT  5.285 0.785 5.370 1.075 ;
        RECT  4.905 0.185 4.935 0.460 ;
        RECT  4.905 0.785 4.935 1.075 ;
        RECT  4.835 0.545 4.935 0.615 ;
        RECT  4.750 0.545 4.835 0.920 ;
        RECT  4.255 0.850 4.750 0.920 ;
        RECT  4.505 0.695 4.620 0.765 ;
        RECT  4.505 0.395 4.615 0.465 ;
        RECT  4.435 0.395 4.505 0.765 ;
        RECT  4.335 0.575 4.435 0.685 ;
        RECT  4.185 0.340 4.255 0.920 ;
        RECT  3.545 0.340 4.185 0.410 ;
        RECT  3.955 0.850 4.185 0.920 ;
        RECT  3.880 0.550 4.085 0.620 ;
        RECT  3.810 0.550 3.880 0.915 ;
        RECT  3.245 0.845 3.810 0.915 ;
        RECT  3.475 0.340 3.545 0.640 ;
        RECT  3.310 0.995 3.420 1.075 ;
        RECT  3.095 0.995 3.310 1.065 ;
        RECT  3.175 0.335 3.245 0.915 ;
        RECT  3.095 0.195 3.170 0.265 ;
        RECT  3.025 0.195 3.095 1.065 ;
        RECT  2.990 0.870 3.025 1.065 ;
        RECT  2.580 0.870 2.990 0.940 ;
        RECT  2.845 0.185 2.955 0.330 ;
        RECT  2.580 0.260 2.845 0.330 ;
        RECT  2.580 0.410 2.670 0.480 ;
        RECT  2.510 0.195 2.580 0.330 ;
        RECT  2.510 0.410 2.580 0.940 ;
        RECT  1.670 0.195 2.510 0.265 ;
        RECT  2.020 0.870 2.510 0.940 ;
        RECT  2.370 0.345 2.440 0.765 ;
        RECT  1.985 0.695 2.370 0.765 ;
        RECT  1.950 0.870 2.020 1.065 ;
        RECT  1.915 0.575 1.985 0.765 ;
        RECT  1.610 0.995 1.950 1.065 ;
        RECT  1.820 0.335 1.890 0.405 ;
        RECT  1.820 0.830 1.870 0.900 ;
        RECT  1.750 0.335 1.820 0.900 ;
        RECT  1.600 0.195 1.670 0.925 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.585 0.815 1.600 0.925 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQD4BWP40

MACRO SDFNSNQND0BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.055 ;
        RECT  4.635 0.185 4.655 0.300 ;
        RECT  4.635 0.915 4.655 1.055 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.610 2.835 0.680 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.180 ;
        RECT  4.150 -0.115 4.420 0.115 ;
        RECT  4.030 -0.115 4.150 0.210 ;
        RECT  3.730 -0.115 4.030 0.115 ;
        RECT  3.610 -0.115 3.730 0.210 ;
        RECT  2.805 -0.115 3.610 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.145 4.760 1.375 ;
        RECT  4.445 0.915 4.520 1.375 ;
        RECT  3.770 1.145 4.445 1.375 ;
        RECT  3.650 0.985 3.770 1.375 ;
        RECT  2.900 1.145 3.650 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.115 1.145 2.395 1.375 ;
        RECT  1.995 1.050 2.115 1.375 ;
        RECT  1.125 1.145 1.995 1.375 ;
        RECT  0.995 1.120 1.125 1.375 ;
        RECT  0.340 1.145 0.995 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.505 0.525 4.585 0.635 ;
        RECT  4.430 0.280 4.505 0.635 ;
        RECT  3.475 0.280 4.430 0.350 ;
        RECT  4.300 0.420 4.350 0.490 ;
        RECT  4.300 1.005 4.350 1.075 ;
        RECT  4.230 0.420 4.300 1.075 ;
        RECT  4.055 0.585 4.230 0.695 ;
        RECT  3.985 0.920 4.145 0.990 ;
        RECT  3.915 0.430 3.985 0.990 ;
        RECT  3.625 0.430 3.915 0.500 ;
        RECT  3.775 0.645 3.845 0.915 ;
        RECT  3.275 0.845 3.775 0.915 ;
        RECT  3.555 0.430 3.625 0.620 ;
        RECT  3.475 0.705 3.570 0.775 ;
        RECT  3.405 0.280 3.475 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.205 0.350 3.275 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.685 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.775 2.685 0.980 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.980 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  1.820 0.910 2.555 0.980 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.830 ;
        RECT  1.750 0.910 1.820 1.065 ;
        RECT  1.750 0.760 1.795 0.830 ;
        RECT  1.610 0.995 1.750 1.065 ;
        RECT  1.605 0.195 1.675 0.910 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.565 0.840 1.605 0.910 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.350 0.960 0.420 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.350 0.865 0.910 ;
        RECT  0.645 0.875 0.715 1.050 ;
        RECT  0.555 0.530 0.610 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQND0BWP40

MACRO SDFNSNQND1BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.075 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.685 4.655 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.210 ;
        RECT  4.150 -0.115 4.420 0.115 ;
        RECT  4.030 -0.115 4.150 0.210 ;
        RECT  3.730 -0.115 4.030 0.115 ;
        RECT  3.610 -0.115 3.730 0.210 ;
        RECT  2.805 -0.115 3.610 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.145 4.760 1.375 ;
        RECT  4.445 0.720 4.520 1.375 ;
        RECT  3.770 1.145 4.445 1.375 ;
        RECT  3.640 1.020 3.770 1.375 ;
        RECT  2.900 1.145 3.640 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.115 1.145 2.395 1.375 ;
        RECT  1.995 1.050 2.115 1.375 ;
        RECT  1.120 1.145 1.995 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.505 0.525 4.585 0.635 ;
        RECT  4.430 0.280 4.505 0.635 ;
        RECT  3.475 0.280 4.430 0.350 ;
        RECT  4.300 0.420 4.350 0.490 ;
        RECT  4.300 1.000 4.350 1.070 ;
        RECT  4.230 0.420 4.300 1.070 ;
        RECT  4.055 0.585 4.230 0.695 ;
        RECT  4.055 0.805 4.125 1.065 ;
        RECT  3.985 0.805 4.055 0.875 ;
        RECT  3.915 0.430 3.985 0.875 ;
        RECT  3.625 0.430 3.915 0.500 ;
        RECT  3.775 0.645 3.845 0.915 ;
        RECT  3.285 0.845 3.775 0.915 ;
        RECT  3.555 0.430 3.625 0.620 ;
        RECT  3.475 0.705 3.570 0.775 ;
        RECT  3.405 0.280 3.475 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.215 0.335 3.285 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.685 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.775 2.685 0.980 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.980 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  1.820 0.910 2.555 0.980 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.830 ;
        RECT  1.750 0.910 1.820 1.065 ;
        RECT  1.750 0.760 1.795 0.830 ;
        RECT  1.610 0.995 1.750 1.065 ;
        RECT  1.605 0.195 1.675 0.910 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.565 0.840 1.605 0.910 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQND1BWP40

MACRO SDFNSNQND2BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.115 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.660 0.370 4.725 0.880 ;
        RECT  4.655 0.195 4.660 1.075 ;
        RECT  4.585 0.195 4.655 0.445 ;
        RECT  4.585 0.805 4.655 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.680 0.605 2.835 0.675 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.275 ;
        RECT  4.490 -0.115 4.775 0.115 ;
        RECT  4.370 -0.115 4.490 0.180 ;
        RECT  4.095 -0.115 4.370 0.115 ;
        RECT  3.975 -0.115 4.095 0.210 ;
        RECT  3.695 -0.115 3.975 0.115 ;
        RECT  3.555 -0.115 3.695 0.210 ;
        RECT  2.780 -0.115 3.555 0.115 ;
        RECT  2.660 -0.115 2.780 0.190 ;
        RECT  2.065 -0.115 2.660 0.115 ;
        RECT  1.935 -0.115 2.065 0.125 ;
        RECT  1.145 -0.115 1.935 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.950 4.845 1.375 ;
        RECT  4.465 1.145 4.775 1.375 ;
        RECT  4.395 0.725 4.465 1.375 ;
        RECT  3.720 1.145 4.395 1.375 ;
        RECT  3.640 0.985 3.720 1.375 ;
        RECT  2.875 1.145 3.640 1.375 ;
        RECT  2.745 1.050 2.875 1.375 ;
        RECT  2.485 1.145 2.745 1.375 ;
        RECT  2.355 1.050 2.485 1.375 ;
        RECT  2.220 1.145 2.355 1.375 ;
        RECT  2.090 1.070 2.220 1.375 ;
        RECT  1.120 1.145 2.090 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.495 0.525 4.585 0.635 ;
        RECT  4.420 0.280 4.495 0.635 ;
        RECT  3.490 0.280 4.420 0.350 ;
        RECT  4.255 0.810 4.300 0.880 ;
        RECT  4.080 0.420 4.295 0.495 ;
        RECT  4.185 0.690 4.255 0.880 ;
        RECT  4.080 0.690 4.185 0.770 ;
        RECT  3.940 0.855 4.115 0.925 ;
        RECT  4.010 0.420 4.080 0.770 ;
        RECT  3.870 0.430 3.940 0.925 ;
        RECT  3.650 0.430 3.870 0.500 ;
        RECT  3.720 0.635 3.790 0.915 ;
        RECT  3.265 0.845 3.720 0.915 ;
        RECT  3.580 0.430 3.650 0.605 ;
        RECT  3.500 0.535 3.580 0.605 ;
        RECT  3.415 0.705 3.555 0.775 ;
        RECT  3.415 0.280 3.490 0.395 ;
        RECT  3.340 0.995 3.450 1.075 ;
        RECT  3.345 0.280 3.415 0.775 ;
        RECT  3.115 0.995 3.340 1.065 ;
        RECT  3.195 0.335 3.265 0.915 ;
        RECT  3.115 0.195 3.175 0.265 ;
        RECT  3.045 0.195 3.115 1.065 ;
        RECT  3.020 0.870 3.045 1.065 ;
        RECT  2.590 0.870 3.020 0.940 ;
        RECT  2.855 0.185 2.965 0.330 ;
        RECT  2.590 0.260 2.855 0.330 ;
        RECT  2.590 0.410 2.690 0.480 ;
        RECT  2.520 0.195 2.590 0.330 ;
        RECT  2.520 0.410 2.590 0.940 ;
        RECT  1.670 0.195 2.520 0.265 ;
        RECT  2.020 0.870 2.520 0.940 ;
        RECT  2.370 0.345 2.440 0.765 ;
        RECT  1.985 0.695 2.370 0.765 ;
        RECT  1.950 0.870 2.020 1.065 ;
        RECT  1.915 0.575 1.985 0.765 ;
        RECT  1.610 0.995 1.950 1.065 ;
        RECT  1.820 0.335 1.890 0.405 ;
        RECT  1.820 0.830 1.870 0.900 ;
        RECT  1.750 0.335 1.820 0.900 ;
        RECT  1.600 0.195 1.670 0.925 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.585 0.815 1.600 0.925 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQND2BWP40

MACRO SDFNSNQND4BWP40
    CLASS CORE ;
    FOREIGN SDFNSNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.425 0.190 5.520 0.440 ;
        RECT  5.425 0.745 5.520 1.005 ;
        RECT  5.355 0.355 5.425 0.440 ;
        RECT  5.355 0.745 5.425 0.830 ;
        RECT  5.145 0.355 5.355 0.830 ;
        RECT  5.120 0.355 5.145 0.475 ;
        RECT  5.120 0.710 5.145 0.830 ;
        RECT  5.050 0.205 5.120 0.475 ;
        RECT  5.050 0.710 5.120 1.020 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.430 ;
        RECT  5.310 -0.115 5.610 0.115 ;
        RECT  5.235 -0.115 5.310 0.270 ;
        RECT  4.950 -0.115 5.235 0.115 ;
        RECT  4.830 -0.115 4.950 0.210 ;
        RECT  4.560 -0.115 4.830 0.115 ;
        RECT  4.440 -0.115 4.560 0.210 ;
        RECT  4.130 -0.115 4.440 0.115 ;
        RECT  4.005 -0.115 4.130 0.210 ;
        RECT  3.760 -0.115 4.005 0.115 ;
        RECT  3.635 -0.115 3.760 0.210 ;
        RECT  2.805 -0.115 3.635 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.600 0.705 5.690 1.375 ;
        RECT  5.325 1.145 5.600 1.375 ;
        RECT  5.215 0.905 5.325 1.375 ;
        RECT  4.930 1.145 5.215 1.375 ;
        RECT  4.855 0.725 4.930 1.375 ;
        RECT  4.165 1.145 4.855 1.375 ;
        RECT  4.035 1.040 4.165 1.375 ;
        RECT  3.760 1.145 4.035 1.375 ;
        RECT  3.620 1.050 3.760 1.375 ;
        RECT  2.900 1.145 3.620 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.115 1.145 2.395 1.375 ;
        RECT  1.995 1.050 2.115 1.375 ;
        RECT  1.120 1.145 1.995 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.190 5.520 0.440 ;
        RECT  5.425 0.745 5.520 1.005 ;
        RECT  5.050 0.205 5.075 0.475 ;
        RECT  5.050 0.710 5.075 1.020 ;
        RECT  4.915 0.545 5.065 0.620 ;
        RECT  4.840 0.280 4.915 0.620 ;
        RECT  3.950 0.280 4.840 0.350 ;
        RECT  4.710 0.420 4.760 0.490 ;
        RECT  4.710 0.810 4.760 0.880 ;
        RECT  4.640 0.420 4.710 0.880 ;
        RECT  4.485 0.585 4.640 0.695 ;
        RECT  4.465 0.805 4.535 1.065 ;
        RECT  4.405 0.805 4.465 0.875 ;
        RECT  4.335 0.430 4.405 0.875 ;
        RECT  4.090 0.430 4.335 0.500 ;
        RECT  4.185 0.645 4.255 0.915 ;
        RECT  3.285 0.845 4.185 0.915 ;
        RECT  4.020 0.430 4.090 0.565 ;
        RECT  3.765 0.495 4.020 0.565 ;
        RECT  3.830 0.280 3.950 0.400 ;
        RECT  3.575 0.705 3.950 0.775 ;
        RECT  3.575 0.280 3.830 0.350 ;
        RECT  3.655 0.495 3.765 0.625 ;
        RECT  3.505 0.280 3.575 0.775 ;
        RECT  3.450 0.280 3.505 0.415 ;
        RECT  3.445 0.705 3.505 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.215 0.335 3.285 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.685 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.775 2.685 0.980 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.980 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  1.820 0.910 2.555 0.980 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.830 ;
        RECT  1.750 0.910 1.820 1.065 ;
        RECT  1.750 0.760 1.795 0.830 ;
        RECT  1.610 0.995 1.750 1.065 ;
        RECT  1.605 0.195 1.675 0.910 ;
        RECT  1.490 0.995 1.610 1.075 ;
        RECT  1.565 0.840 1.605 0.910 ;
        RECT  1.415 0.200 1.485 0.405 ;
        RECT  1.335 0.565 1.485 0.635 ;
        RECT  1.320 0.855 1.485 0.925 ;
        RECT  0.640 0.200 1.415 0.270 ;
        RECT  1.265 0.350 1.335 0.785 ;
        RECT  1.250 0.855 1.320 1.050 ;
        RECT  1.200 0.350 1.265 0.420 ;
        RECT  1.190 0.715 1.265 0.785 ;
        RECT  0.715 0.980 1.250 1.050 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFNSNQND4BWP40

MACRO SDFQD0BWP40
    CLASS CORE ;
    FOREIGN SDFQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.630 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.255 ;
        RECT  2.655 -0.115 3.375 0.115 ;
        RECT  2.535 -0.115 2.655 0.125 ;
        RECT  2.040 -0.115 2.535 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.130 -0.115 1.920 0.115 ;
        RECT  1.000 -0.115 1.130 0.125 ;
        RECT  0.340 -0.115 1.000 0.115 ;
        RECT  0.220 -0.115 0.340 0.260 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.640 1.145 3.310 1.375 ;
        RECT  2.520 0.970 2.640 1.375 ;
        RECT  2.060 1.145 2.520 1.375 ;
        RECT  1.940 0.855 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.980 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.810 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.740 3.785 0.810 ;
        RECT  3.565 0.195 3.635 0.465 ;
        RECT  3.565 0.740 3.635 0.960 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.335 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.005 0.860 3.415 0.930 ;
        RECT  3.265 0.395 3.335 0.600 ;
        RECT  3.115 0.195 3.195 0.780 ;
        RECT  2.930 0.195 3.115 0.265 ;
        RECT  2.935 0.345 3.005 0.930 ;
        RECT  2.900 0.345 2.935 0.465 ;
        RECT  2.830 0.185 2.930 0.265 ;
        RECT  2.800 0.185 2.830 0.875 ;
        RECT  2.760 0.195 2.800 0.875 ;
        RECT  2.420 0.195 2.760 0.265 ;
        RECT  2.430 0.785 2.760 0.875 ;
        RECT  2.610 0.520 2.690 0.640 ;
        RECT  2.155 0.520 2.610 0.610 ;
        RECT  2.345 0.785 2.430 1.015 ;
        RECT  2.350 0.195 2.420 0.415 ;
        RECT  1.680 0.195 2.350 0.265 ;
        RECT  2.000 0.370 2.260 0.440 ;
        RECT  2.165 0.690 2.235 0.945 ;
        RECT  2.000 0.690 2.165 0.760 ;
        RECT  1.930 0.370 2.000 0.760 ;
        RECT  1.880 0.620 1.930 0.760 ;
        RECT  1.810 0.370 1.860 0.490 ;
        RECT  1.810 0.830 1.860 0.925 ;
        RECT  1.740 0.370 1.810 0.925 ;
        RECT  1.605 0.995 1.770 1.065 ;
        RECT  1.600 0.350 1.670 0.775 ;
        RECT  1.535 0.845 1.605 1.065 ;
        RECT  1.530 0.705 1.600 0.775 ;
        RECT  1.440 0.845 1.535 0.915 ;
        RECT  1.440 0.345 1.505 0.505 ;
        RECT  0.585 0.195 1.485 0.265 ;
        RECT  0.590 0.985 1.455 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.150 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.910 ;
        RECT  0.125 0.840 0.525 0.910 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.105 0.840 0.125 1.070 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.210 0.525 2.280 0.595 ;
        RECT  1.600 0.525 1.670 0.595 ;
        LAYER M2 ;
        RECT  1.550 0.525 2.330 0.595 ;
    END
END SDFQD0BWP40

MACRO SDFQD1BWP40
    CLASS CORE ;
    FOREIGN SDFQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.605 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.025 1.065 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.605 -0.115 3.375 0.115 ;
        RECT  2.535 -0.115 2.605 0.290 ;
        RECT  2.040 -0.115 2.535 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.110 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 0.890 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 0.855 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.765 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.695 3.785 0.765 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.485 0.545 3.590 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.950 0.350 3.020 0.930 ;
        RECT  2.790 0.195 2.860 0.810 ;
        RECT  2.430 0.360 2.790 0.430 ;
        RECT  2.430 0.720 2.790 0.810 ;
        RECT  2.330 0.535 2.710 0.615 ;
        RECT  2.350 0.195 2.430 0.430 ;
        RECT  2.345 0.720 2.430 0.920 ;
        RECT  1.680 0.195 2.350 0.265 ;
        RECT  2.100 0.525 2.330 0.615 ;
        RECT  2.030 0.375 2.270 0.445 ;
        RECT  2.155 0.695 2.250 0.945 ;
        RECT  2.030 0.695 2.155 0.765 ;
        RECT  1.960 0.375 2.030 0.765 ;
        RECT  1.890 0.620 1.960 0.765 ;
        RECT  1.820 0.380 1.880 0.480 ;
        RECT  1.820 0.845 1.840 0.925 ;
        RECT  1.750 0.380 1.820 0.925 ;
        RECT  1.600 0.995 1.770 1.065 ;
        RECT  1.610 0.350 1.680 0.760 ;
        RECT  1.530 0.690 1.610 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.440 0.345 1.540 0.505 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  0.575 0.195 1.485 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.210 0.525 2.280 0.595 ;
        RECT  1.610 0.525 1.680 0.595 ;
        LAYER M2 ;
        RECT  1.560 0.525 2.330 0.595 ;
    END
END SDFQD1BWP40

MACRO SDFQD2BWP40
    CLASS CORE ;
    FOREIGN SDFQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.605 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.120000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.195 4.040 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.023600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 -0.115 4.340 0.115 ;
        RECT  4.195 -0.115 4.270 0.455 ;
        RECT  3.815 -0.115 4.195 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.605 -0.115 3.375 0.115 ;
        RECT  2.535 -0.115 2.605 0.255 ;
        RECT  2.040 -0.115 2.535 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.110 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.275 1.145 4.340 1.375 ;
        RECT  4.205 0.705 4.275 1.375 ;
        RECT  3.815 1.145 4.205 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 0.890 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 0.855 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.785 0.395 3.855 0.765 ;
        RECT  3.635 0.395 3.785 0.465 ;
        RECT  3.635 0.695 3.785 0.765 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 0.980 ;
        RECT  3.485 0.545 3.600 0.615 ;
        RECT  3.340 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.270 0.395 3.340 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.950 0.350 3.020 0.930 ;
        RECT  2.790 0.195 2.860 0.810 ;
        RECT  2.430 0.350 2.790 0.430 ;
        RECT  2.430 0.720 2.790 0.810 ;
        RECT  2.330 0.535 2.710 0.615 ;
        RECT  2.350 0.195 2.430 0.430 ;
        RECT  2.345 0.720 2.430 0.910 ;
        RECT  1.680 0.195 2.350 0.265 ;
        RECT  2.100 0.525 2.330 0.615 ;
        RECT  2.030 0.375 2.270 0.445 ;
        RECT  2.155 0.695 2.250 0.945 ;
        RECT  2.030 0.695 2.155 0.765 ;
        RECT  1.960 0.375 2.030 0.765 ;
        RECT  1.890 0.620 1.960 0.765 ;
        RECT  1.820 0.380 1.880 0.480 ;
        RECT  1.820 0.845 1.840 0.925 ;
        RECT  1.750 0.380 1.820 0.925 ;
        RECT  1.600 0.995 1.770 1.065 ;
        RECT  1.610 0.350 1.680 0.760 ;
        RECT  1.530 0.690 1.610 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.440 0.345 1.540 0.505 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  0.575 0.195 1.485 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.210 0.525 2.280 0.595 ;
        RECT  1.610 0.525 1.680 0.595 ;
        LAYER M2 ;
        RECT  1.560 0.525 2.330 0.595 ;
    END
END SDFQD2BWP40

MACRO SDFQD4BWP40
    CLASS CORE ;
    FOREIGN SDFQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.605 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.740 4.405 1.040 ;
        RECT  4.305 0.195 4.390 0.455 ;
        RECT  4.235 0.370 4.305 0.455 ;
        RECT  4.235 0.740 4.305 0.825 ;
        RECT  4.025 0.370 4.235 0.825 ;
        RECT  4.000 0.370 4.025 0.465 ;
        RECT  4.005 0.725 4.025 0.825 ;
        RECT  3.920 0.725 4.005 1.055 ;
        RECT  3.920 0.195 4.000 0.465 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.290 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.565 -0.115 4.620 0.115 ;
        RECT  4.485 -0.115 4.565 0.455 ;
        RECT  4.190 -0.115 4.485 0.115 ;
        RECT  4.115 -0.115 4.190 0.285 ;
        RECT  3.805 -0.115 4.115 0.115 ;
        RECT  3.735 -0.115 3.805 0.315 ;
        RECT  3.415 -0.115 3.735 0.115 ;
        RECT  3.345 -0.115 3.415 0.315 ;
        RECT  2.595 -0.115 3.345 0.115 ;
        RECT  2.525 -0.115 2.595 0.255 ;
        RECT  2.030 -0.115 2.525 0.115 ;
        RECT  1.910 -0.115 2.030 0.125 ;
        RECT  1.110 -0.115 1.910 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.565 1.145 4.620 1.375 ;
        RECT  4.485 0.690 4.565 1.375 ;
        RECT  4.210 1.145 4.485 1.375 ;
        RECT  4.090 0.905 4.210 1.375 ;
        RECT  3.805 1.145 4.090 1.375 ;
        RECT  3.735 0.845 3.805 1.375 ;
        RECT  3.420 1.145 3.735 1.375 ;
        RECT  3.290 1.130 3.420 1.375 ;
        RECT  2.620 1.145 3.290 1.375 ;
        RECT  2.500 0.890 2.620 1.375 ;
        RECT  2.050 1.145 2.500 1.375 ;
        RECT  1.930 0.855 2.050 1.375 ;
        RECT  1.110 1.145 1.930 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.740 4.405 1.040 ;
        RECT  4.305 0.195 4.390 0.455 ;
        RECT  3.920 0.195 3.955 0.465 ;
        RECT  3.920 0.725 3.955 1.055 ;
        RECT  3.835 0.545 3.950 0.615 ;
        RECT  3.765 0.395 3.835 0.765 ;
        RECT  3.615 0.395 3.765 0.465 ;
        RECT  3.615 0.695 3.765 0.765 ;
        RECT  3.545 0.185 3.615 0.465 ;
        RECT  3.475 0.545 3.615 0.615 ;
        RECT  3.545 0.695 3.615 1.025 ;
        RECT  3.315 0.395 3.545 0.465 ;
        RECT  3.395 0.545 3.475 0.930 ;
        RECT  3.000 0.860 3.395 0.930 ;
        RECT  3.245 0.395 3.315 0.600 ;
        RECT  3.095 0.195 3.175 0.780 ;
        RECT  2.850 0.195 3.095 0.265 ;
        RECT  2.930 0.350 3.000 0.930 ;
        RECT  2.780 0.195 2.850 0.820 ;
        RECT  2.420 0.350 2.780 0.430 ;
        RECT  2.420 0.745 2.780 0.820 ;
        RECT  2.070 0.525 2.700 0.610 ;
        RECT  2.340 0.195 2.420 0.430 ;
        RECT  2.335 0.745 2.420 0.910 ;
        RECT  1.670 0.195 2.340 0.265 ;
        RECT  2.000 0.375 2.250 0.445 ;
        RECT  2.150 0.690 2.225 0.945 ;
        RECT  2.000 0.690 2.150 0.760 ;
        RECT  1.930 0.375 2.000 0.760 ;
        RECT  1.870 0.620 1.930 0.760 ;
        RECT  1.800 0.365 1.850 0.485 ;
        RECT  1.800 0.830 1.850 0.900 ;
        RECT  1.730 0.365 1.800 0.900 ;
        RECT  1.595 0.995 1.760 1.065 ;
        RECT  1.590 0.345 1.660 0.760 ;
        RECT  1.525 0.845 1.595 1.065 ;
        RECT  1.520 0.690 1.590 0.760 ;
        RECT  1.440 0.845 1.525 0.915 ;
        RECT  1.440 0.345 1.495 0.505 ;
        RECT  0.575 0.195 1.475 0.265 ;
        RECT  0.595 0.985 1.445 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.200 0.525 2.270 0.595 ;
        RECT  1.590 0.525 1.660 0.595 ;
        LAYER M2 ;
        RECT  1.540 0.525 2.320 0.595 ;
    END
END SDFQD4BWP40

MACRO SDFQND0BWP40
    CLASS CORE ;
    FOREIGN SDFQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.620 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.185 4.025 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.885 0.640 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.705 -0.115 3.375 0.115 ;
        RECT  2.560 -0.115 2.705 0.125 ;
        RECT  2.040 -0.115 2.560 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.120 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.120 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.895 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.640 1.145 3.310 1.375 ;
        RECT  2.520 0.970 2.640 1.375 ;
        RECT  2.060 1.145 2.520 1.375 ;
        RECT  1.940 0.855 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.810 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.740 3.775 0.810 ;
        RECT  3.485 0.545 3.670 0.615 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.740 3.635 1.025 ;
        RECT  3.325 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.005 0.860 3.415 0.930 ;
        RECT  3.255 0.395 3.325 0.600 ;
        RECT  3.105 0.195 3.185 0.780 ;
        RECT  2.930 0.195 3.105 0.265 ;
        RECT  2.935 0.350 3.005 0.930 ;
        RECT  2.900 0.350 2.935 0.470 ;
        RECT  2.830 0.185 2.930 0.265 ;
        RECT  2.800 0.185 2.830 0.850 ;
        RECT  2.760 0.195 2.800 0.850 ;
        RECT  1.680 0.195 2.760 0.265 ;
        RECT  2.415 0.770 2.760 0.850 ;
        RECT  2.590 0.520 2.690 0.640 ;
        RECT  2.355 0.545 2.590 0.615 ;
        RECT  2.345 0.770 2.415 0.910 ;
        RECT  2.105 0.525 2.355 0.615 ;
        RECT  2.035 0.355 2.260 0.425 ;
        RECT  2.150 0.715 2.250 0.865 ;
        RECT  2.035 0.715 2.150 0.785 ;
        RECT  1.960 0.355 2.035 0.785 ;
        RECT  1.870 0.605 1.960 0.740 ;
        RECT  1.800 0.390 1.880 0.465 ;
        RECT  1.800 0.805 1.815 0.925 ;
        RECT  1.730 0.390 1.800 0.925 ;
        RECT  1.600 0.995 1.750 1.065 ;
        RECT  1.590 0.350 1.660 0.765 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.520 0.695 1.590 0.765 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  1.440 0.345 1.495 0.505 ;
        RECT  0.585 0.195 1.460 0.265 ;
        RECT  0.580 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.140 0.845 1.370 0.915 ;
        RECT  0.805 0.335 0.910 0.405 ;
        RECT  0.805 0.845 0.910 0.915 ;
        RECT  0.735 0.335 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.220 0.525 2.290 0.595 ;
        RECT  1.590 0.525 1.660 0.595 ;
        LAYER M2 ;
        RECT  1.540 0.525 2.340 0.595 ;
    END
END SDFQND0BWP40

MACRO SDFQND1BWP40
    CLASS CORE ;
    FOREIGN SDFQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.060 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.605 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.185 4.025 1.065 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 -0.115 4.060 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.605 -0.115 3.375 0.115 ;
        RECT  2.535 -0.115 2.605 0.255 ;
        RECT  2.040 -0.115 2.535 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.110 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.815 1.145 4.060 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 0.890 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 0.870 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.765 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.695 3.775 0.765 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 1.025 ;
        RECT  3.485 0.545 3.630 0.615 ;
        RECT  3.330 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.260 0.395 3.330 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.950 0.350 3.020 0.930 ;
        RECT  2.790 0.195 2.860 0.800 ;
        RECT  2.430 0.350 2.790 0.430 ;
        RECT  2.430 0.710 2.790 0.800 ;
        RECT  2.330 0.535 2.710 0.615 ;
        RECT  2.350 0.195 2.430 0.430 ;
        RECT  2.345 0.710 2.430 0.910 ;
        RECT  1.680 0.195 2.350 0.265 ;
        RECT  2.100 0.525 2.330 0.615 ;
        RECT  2.030 0.375 2.270 0.445 ;
        RECT  2.155 0.695 2.250 0.940 ;
        RECT  2.030 0.695 2.155 0.765 ;
        RECT  1.960 0.375 2.030 0.765 ;
        RECT  1.880 0.575 1.960 0.700 ;
        RECT  1.810 0.380 1.880 0.480 ;
        RECT  1.810 0.805 1.825 0.925 ;
        RECT  1.740 0.380 1.810 0.925 ;
        RECT  1.600 0.995 1.770 1.065 ;
        RECT  1.600 0.370 1.670 0.760 ;
        RECT  1.530 0.690 1.600 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.440 0.345 1.530 0.505 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  0.575 0.195 1.485 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.210 0.525 2.280 0.595 ;
        RECT  1.600 0.525 1.670 0.595 ;
        LAYER M2 ;
        RECT  1.550 0.525 2.330 0.595 ;
    END
END SDFQND1BWP40

MACRO SDFQND2BWP40
    CLASS CORE ;
    FOREIGN SDFQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.605 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.124000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.935 0.185 4.050 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 -0.115 4.340 0.115 ;
        RECT  4.165 -0.115 4.270 0.480 ;
        RECT  3.815 -0.115 4.165 0.115 ;
        RECT  3.745 -0.115 3.815 0.315 ;
        RECT  3.445 -0.115 3.745 0.115 ;
        RECT  3.375 -0.115 3.445 0.315 ;
        RECT  2.605 -0.115 3.375 0.115 ;
        RECT  2.535 -0.115 2.605 0.255 ;
        RECT  2.040 -0.115 2.535 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.110 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.255 1.145 4.340 1.375 ;
        RECT  4.145 0.715 4.255 1.375 ;
        RECT  3.815 1.145 4.145 1.375 ;
        RECT  3.745 0.845 3.815 1.375 ;
        RECT  3.440 1.145 3.745 1.375 ;
        RECT  3.310 1.130 3.440 1.375 ;
        RECT  2.630 1.145 3.310 1.375 ;
        RECT  2.510 0.890 2.630 1.375 ;
        RECT  2.060 1.145 2.510 1.375 ;
        RECT  1.940 0.870 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.775 0.395 3.845 0.765 ;
        RECT  3.635 0.395 3.775 0.465 ;
        RECT  3.635 0.695 3.775 0.765 ;
        RECT  3.485 0.545 3.650 0.615 ;
        RECT  3.565 0.185 3.635 0.465 ;
        RECT  3.565 0.695 3.635 1.025 ;
        RECT  3.330 0.395 3.565 0.465 ;
        RECT  3.415 0.545 3.485 0.930 ;
        RECT  3.020 0.860 3.415 0.930 ;
        RECT  3.260 0.395 3.330 0.600 ;
        RECT  3.110 0.195 3.190 0.780 ;
        RECT  2.860 0.195 3.110 0.265 ;
        RECT  2.950 0.350 3.020 0.930 ;
        RECT  2.790 0.195 2.860 0.800 ;
        RECT  2.430 0.350 2.790 0.430 ;
        RECT  2.430 0.710 2.790 0.800 ;
        RECT  2.330 0.535 2.710 0.615 ;
        RECT  2.350 0.195 2.430 0.430 ;
        RECT  2.345 0.710 2.430 0.910 ;
        RECT  1.680 0.195 2.350 0.265 ;
        RECT  2.100 0.525 2.330 0.615 ;
        RECT  2.030 0.375 2.270 0.445 ;
        RECT  2.155 0.695 2.250 0.940 ;
        RECT  2.030 0.695 2.155 0.765 ;
        RECT  1.960 0.375 2.030 0.765 ;
        RECT  1.880 0.575 1.960 0.700 ;
        RECT  1.810 0.380 1.880 0.480 ;
        RECT  1.810 0.805 1.825 0.925 ;
        RECT  1.740 0.380 1.810 0.925 ;
        RECT  1.600 0.995 1.770 1.065 ;
        RECT  1.600 0.370 1.670 0.760 ;
        RECT  1.530 0.690 1.600 0.760 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.440 0.345 1.530 0.505 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  0.575 0.195 1.485 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.140 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.900 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.210 0.525 2.280 0.595 ;
        RECT  1.600 0.525 1.670 0.595 ;
        LAYER M2 ;
        RECT  1.550 0.525 2.330 0.595 ;
    END
END SDFQND2BWP40

MACRO SDFQND4BWP40
    CLASS CORE ;
    FOREIGN SDFQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.495 0.665 0.625 ;
        RECT  0.360 0.495 0.445 0.705 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.350 0.600 0.425 ;
        RECT  0.175 0.350 0.260 0.765 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 0.210 4.820 0.470 ;
        RECT  4.725 0.705 4.820 1.015 ;
        RECT  4.655 0.370 4.725 0.470 ;
        RECT  4.655 0.705 4.725 0.815 ;
        RECT  4.445 0.370 4.655 0.815 ;
        RECT  4.420 0.370 4.445 0.475 ;
        RECT  4.420 0.695 4.445 0.815 ;
        RECT  4.350 0.205 4.420 0.475 ;
        RECT  4.350 0.695 4.420 1.005 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.023800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.085 0.765 ;
        RECT  0.890 0.635 1.010 0.765 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.300 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 -0.115 5.040 0.115 ;
        RECT  4.915 -0.115 4.985 0.410 ;
        RECT  4.630 -0.115 4.915 0.115 ;
        RECT  4.510 -0.115 4.630 0.290 ;
        RECT  4.225 -0.115 4.510 0.115 ;
        RECT  4.155 -0.115 4.225 0.305 ;
        RECT  3.855 -0.115 4.155 0.115 ;
        RECT  3.785 -0.115 3.855 0.305 ;
        RECT  3.000 -0.115 3.785 0.115 ;
        RECT  2.910 -0.115 3.000 0.170 ;
        RECT  2.615 -0.115 2.910 0.115 ;
        RECT  2.540 -0.115 2.615 0.280 ;
        RECT  2.040 -0.115 2.540 0.115 ;
        RECT  1.920 -0.115 2.040 0.125 ;
        RECT  1.110 -0.115 1.920 0.115 ;
        RECT  0.990 -0.115 1.110 0.125 ;
        RECT  0.340 -0.115 0.990 0.115 ;
        RECT  0.220 -0.115 0.340 0.270 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.985 1.145 5.040 1.375 ;
        RECT  4.915 0.695 4.985 1.375 ;
        RECT  4.630 1.145 4.915 1.375 ;
        RECT  4.510 0.885 4.630 1.375 ;
        RECT  4.225 1.145 4.510 1.375 ;
        RECT  4.155 0.845 4.225 1.375 ;
        RECT  3.850 1.145 4.155 1.375 ;
        RECT  3.720 1.130 3.850 1.375 ;
        RECT  3.040 1.145 3.720 1.375 ;
        RECT  2.920 0.970 3.040 1.375 ;
        RECT  2.650 1.145 2.920 1.375 ;
        RECT  2.530 0.860 2.650 1.375 ;
        RECT  2.060 1.145 2.530 1.375 ;
        RECT  1.940 1.040 2.060 1.375 ;
        RECT  1.110 1.145 1.940 1.375 ;
        RECT  0.990 1.130 1.110 1.375 ;
        RECT  0.340 1.145 0.990 1.375 ;
        RECT  0.220 0.990 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.725 0.210 4.820 0.470 ;
        RECT  4.725 0.705 4.820 1.015 ;
        RECT  4.350 0.205 4.375 0.475 ;
        RECT  4.350 0.695 4.375 1.005 ;
        RECT  4.210 0.385 4.280 0.765 ;
        RECT  4.045 0.385 4.210 0.455 ;
        RECT  4.045 0.695 4.210 0.765 ;
        RECT  3.895 0.545 4.095 0.615 ;
        RECT  3.975 0.195 4.045 0.455 ;
        RECT  3.975 0.695 4.045 0.980 ;
        RECT  3.735 0.385 3.975 0.455 ;
        RECT  3.825 0.545 3.895 0.930 ;
        RECT  3.430 0.860 3.825 0.930 ;
        RECT  3.665 0.385 3.735 0.600 ;
        RECT  3.515 0.195 3.595 0.780 ;
        RECT  3.290 0.195 3.515 0.265 ;
        RECT  3.360 0.345 3.430 0.930 ;
        RECT  3.220 0.195 3.290 0.490 ;
        RECT  3.130 0.830 3.225 0.950 ;
        RECT  3.090 0.420 3.220 0.490 ;
        RECT  3.080 0.210 3.150 0.330 ;
        RECT  2.840 0.830 3.130 0.900 ;
        RECT  3.010 0.420 3.090 0.685 ;
        RECT  2.700 0.250 3.080 0.330 ;
        RECT  2.460 0.420 3.010 0.490 ;
        RECT  2.740 0.830 2.840 0.960 ;
        RECT  2.650 0.560 2.805 0.760 ;
        RECT  2.390 0.195 2.460 0.945 ;
        RECT  1.690 0.195 2.390 0.265 ;
        RECT  2.365 0.805 2.390 0.945 ;
        RECT  2.040 0.865 2.275 0.935 ;
        RECT  2.040 0.335 2.255 0.405 ;
        RECT  2.110 0.520 2.210 0.790 ;
        RECT  1.970 0.335 2.040 0.935 ;
        RECT  1.880 0.535 1.970 0.655 ;
        RECT  1.810 0.375 1.890 0.445 ;
        RECT  1.810 0.805 1.825 0.925 ;
        RECT  1.740 0.375 1.810 0.925 ;
        RECT  1.600 0.995 1.770 1.065 ;
        RECT  1.600 0.350 1.670 0.765 ;
        RECT  1.530 0.690 1.600 0.765 ;
        RECT  1.530 0.845 1.600 1.065 ;
        RECT  1.440 0.845 1.530 0.915 ;
        RECT  1.440 0.345 1.520 0.505 ;
        RECT  0.585 0.195 1.480 0.265 ;
        RECT  0.595 0.985 1.450 1.055 ;
        RECT  1.370 0.345 1.440 0.915 ;
        RECT  1.145 0.345 1.370 0.415 ;
        RECT  1.135 0.845 1.370 0.915 ;
        RECT  0.805 0.845 0.910 0.915 ;
        RECT  0.810 0.335 0.880 0.525 ;
        RECT  0.805 0.455 0.810 0.525 ;
        RECT  0.735 0.455 0.805 0.915 ;
        RECT  0.525 0.695 0.600 0.915 ;
        RECT  0.140 0.845 0.525 0.915 ;
        RECT  0.105 0.845 0.140 1.070 ;
        RECT  0.105 0.185 0.125 0.300 ;
        RECT  0.035 0.185 0.105 1.070 ;
        LAYER VIA1 ;
        RECT  2.685 0.665 2.755 0.735 ;
        RECT  2.125 0.665 2.195 0.735 ;
        RECT  1.600 0.665 1.670 0.735 ;
        LAYER M2 ;
        RECT  1.550 0.665 2.805 0.735 ;
    END
END SDFQND4BWP40

MACRO SDFSNQD0BWP40
    CLASS CORE ;
    FOREIGN SDFSNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.315 4.725 0.925 ;
        RECT  4.635 0.315 4.655 0.435 ;
        RECT  4.635 0.795 4.655 0.925 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.610 2.835 0.680 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 -0.115 4.760 0.115 ;
        RECT  4.440 -0.115 4.520 0.425 ;
        RECT  4.125 -0.115 4.440 0.115 ;
        RECT  4.055 -0.115 4.125 0.280 ;
        RECT  3.740 -0.115 4.055 0.115 ;
        RECT  3.620 -0.115 3.740 0.280 ;
        RECT  2.805 -0.115 3.620 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.760 1.375 ;
        RECT  4.420 1.080 4.540 1.375 ;
        RECT  3.740 1.145 4.420 1.375 ;
        RECT  3.620 0.860 3.740 1.375 ;
        RECT  2.900 1.145 3.620 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.205 1.145 2.395 1.375 ;
        RECT  2.085 1.070 2.205 1.375 ;
        RECT  1.120 1.145 2.085 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.525 4.585 0.635 ;
        RECT  4.490 0.525 4.565 1.010 ;
        RECT  4.120 0.940 4.490 1.010 ;
        RECT  4.255 0.325 4.325 0.870 ;
        RECT  4.190 0.580 4.255 0.700 ;
        RECT  4.050 0.350 4.120 1.010 ;
        RECT  3.590 0.350 4.050 0.420 ;
        RECT  3.910 0.615 3.980 0.780 ;
        RECT  3.325 0.710 3.910 0.780 ;
        RECT  3.520 0.350 3.590 0.610 ;
        RECT  3.350 0.995 3.460 1.075 ;
        RECT  3.135 0.995 3.350 1.065 ;
        RECT  3.285 0.710 3.325 0.925 ;
        RECT  3.215 0.345 3.285 0.925 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.015 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.760 2.720 0.830 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.830 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.945 0.910 2.015 1.050 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.650 0.980 1.945 1.050 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.910 ;
        RECT  1.750 0.840 1.795 0.910 ;
        RECT  1.605 0.195 1.675 0.770 ;
        RECT  1.580 0.840 1.650 1.050 ;
        RECT  1.565 0.700 1.605 0.770 ;
        RECT  1.405 0.840 1.580 0.910 ;
        RECT  0.640 0.200 1.510 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.340 1.405 0.910 ;
        RECT  1.200 0.340 1.335 0.410 ;
        RECT  1.180 0.840 1.335 0.910 ;
        RECT  0.865 0.340 0.960 0.410 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.340 0.865 0.910 ;
        RECT  0.645 0.875 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFSNQD0BWP40

MACRO SDFSNQD1BWP40
    CLASS CORE ;
    FOREIGN SDFSNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.075 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.685 4.655 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.610 2.835 0.680 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.515 -0.115 4.760 0.115 ;
        RECT  4.445 -0.115 4.515 0.440 ;
        RECT  4.125 -0.115 4.445 0.115 ;
        RECT  4.055 -0.115 4.125 0.280 ;
        RECT  3.740 -0.115 4.055 0.115 ;
        RECT  3.620 -0.115 3.740 0.280 ;
        RECT  2.805 -0.115 3.620 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 1.145 4.760 1.375 ;
        RECT  4.420 1.080 4.540 1.375 ;
        RECT  3.740 1.145 4.420 1.375 ;
        RECT  3.620 0.860 3.740 1.375 ;
        RECT  2.900 1.145 3.620 1.375 ;
        RECT  2.780 1.050 2.900 1.375 ;
        RECT  2.515 1.145 2.780 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.205 1.145 2.395 1.375 ;
        RECT  2.085 1.070 2.205 1.375 ;
        RECT  1.120 1.145 2.085 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.565 0.525 4.585 0.635 ;
        RECT  4.490 0.525 4.565 1.010 ;
        RECT  4.120 0.940 4.490 1.010 ;
        RECT  4.255 0.255 4.325 0.870 ;
        RECT  4.190 0.580 4.255 0.700 ;
        RECT  4.050 0.350 4.120 1.010 ;
        RECT  3.590 0.350 4.050 0.420 ;
        RECT  3.910 0.615 3.980 0.780 ;
        RECT  3.325 0.710 3.910 0.780 ;
        RECT  3.520 0.350 3.590 0.610 ;
        RECT  3.350 0.995 3.460 1.075 ;
        RECT  3.135 0.995 3.350 1.065 ;
        RECT  3.285 0.710 3.325 0.925 ;
        RECT  3.215 0.335 3.285 0.925 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.015 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.720 0.480 ;
        RECT  2.625 0.760 2.720 0.830 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.830 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.945 0.910 2.015 1.050 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.650 0.980 1.945 1.050 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.910 ;
        RECT  1.750 0.840 1.795 0.910 ;
        RECT  1.605 0.195 1.675 0.770 ;
        RECT  1.580 0.840 1.650 1.050 ;
        RECT  1.565 0.700 1.605 0.770 ;
        RECT  1.405 0.840 1.580 0.910 ;
        RECT  0.640 0.200 1.510 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.350 1.405 0.910 ;
        RECT  1.200 0.350 1.335 0.420 ;
        RECT  1.190 0.840 1.335 0.910 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFSNQD1BWP40

MACRO SDFSNQD2BWP40
    CLASS CORE ;
    FOREIGN SDFSNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.185 0.385 4.410 0.455 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.660 0.370 4.725 0.880 ;
        RECT  4.655 0.195 4.660 1.075 ;
        RECT  4.585 0.195 4.655 0.445 ;
        RECT  4.585 0.805 4.655 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.670 0.610 2.835 0.680 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.275 ;
        RECT  4.470 -0.115 4.775 0.115 ;
        RECT  4.395 -0.115 4.470 0.260 ;
        RECT  4.060 -0.115 4.395 0.115 ;
        RECT  3.970 -0.115 4.060 0.280 ;
        RECT  3.700 -0.115 3.970 0.115 ;
        RECT  3.580 -0.115 3.700 0.280 ;
        RECT  2.775 -0.115 3.580 0.115 ;
        RECT  2.655 -0.115 2.775 0.190 ;
        RECT  2.025 -0.115 2.655 0.115 ;
        RECT  1.905 -0.115 2.025 0.190 ;
        RECT  1.145 -0.115 1.905 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.950 4.845 1.375 ;
        RECT  4.490 1.145 4.775 1.375 ;
        RECT  4.370 1.080 4.490 1.375 ;
        RECT  3.700 1.145 4.370 1.375 ;
        RECT  3.580 0.865 3.700 1.375 ;
        RECT  2.835 1.145 3.580 1.375 ;
        RECT  2.765 0.855 2.835 1.375 ;
        RECT  2.495 1.145 2.765 1.375 ;
        RECT  2.365 1.050 2.495 1.375 ;
        RECT  2.070 1.145 2.365 1.375 ;
        RECT  1.945 1.050 2.070 1.375 ;
        RECT  1.120 1.145 1.945 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.515 0.520 4.585 0.635 ;
        RECT  4.440 0.520 4.515 0.985 ;
        RECT  4.070 0.915 4.440 0.985 ;
        RECT  4.280 0.365 4.370 0.620 ;
        RECT  4.210 0.225 4.300 0.295 ;
        RECT  4.210 0.775 4.300 0.845 ;
        RECT  4.140 0.225 4.210 0.845 ;
        RECT  4.000 0.350 4.070 0.985 ;
        RECT  3.550 0.350 4.000 0.420 ;
        RECT  3.860 0.615 3.930 0.795 ;
        RECT  3.300 0.725 3.860 0.795 ;
        RECT  3.480 0.350 3.550 0.610 ;
        RECT  3.285 0.995 3.395 1.075 ;
        RECT  3.245 0.725 3.300 0.885 ;
        RECT  3.095 0.995 3.285 1.065 ;
        RECT  3.175 0.335 3.245 0.885 ;
        RECT  3.095 0.195 3.165 0.265 ;
        RECT  3.025 0.195 3.095 1.065 ;
        RECT  2.845 0.185 2.955 0.330 ;
        RECT  2.580 0.260 2.845 0.330 ;
        RECT  2.585 0.410 2.685 0.480 ;
        RECT  2.585 0.825 2.680 0.895 ;
        RECT  2.515 0.410 2.585 0.895 ;
        RECT  2.510 0.195 2.580 0.330 ;
        RECT  2.165 0.195 2.510 0.265 ;
        RECT  2.375 0.365 2.445 0.805 ;
        RECT  2.235 0.735 2.375 0.805 ;
        RECT  2.235 0.355 2.305 0.605 ;
        RECT  2.035 0.535 2.235 0.605 ;
        RECT  2.165 0.735 2.235 0.935 ;
        RECT  2.095 0.195 2.165 0.330 ;
        RECT  1.940 0.735 2.165 0.805 ;
        RECT  1.650 0.260 2.095 0.330 ;
        RECT  1.865 0.680 1.940 0.805 ;
        RECT  1.790 0.400 1.885 0.470 ;
        RECT  1.790 0.885 1.865 0.955 ;
        RECT  1.720 0.400 1.790 0.955 ;
        RECT  1.575 0.260 1.650 0.815 ;
        RECT  0.640 0.200 1.505 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.350 1.405 0.910 ;
        RECT  1.200 0.350 1.335 0.420 ;
        RECT  1.190 0.840 1.335 0.910 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.290 0.385 4.360 0.455 ;
        RECT  2.235 0.385 2.305 0.455 ;
    END
END SDFSNQD2BWP40

MACRO SDFSNQD4BWP40
    CLASS CORE ;
    FOREIGN SDFSNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.185 0.385 4.710 0.455 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.285 0.185 5.380 0.460 ;
        RECT  5.285 0.785 5.370 1.075 ;
        RECT  5.215 0.330 5.285 0.460 ;
        RECT  5.215 0.785 5.285 0.905 ;
        RECT  5.005 0.330 5.215 0.905 ;
        RECT  4.995 0.330 5.005 0.460 ;
        RECT  4.995 0.785 5.005 0.905 ;
        RECT  4.905 0.185 4.995 0.460 ;
        RECT  4.905 0.785 4.995 1.075 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.670 0.605 2.835 0.675 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 -0.115 5.600 0.115 ;
        RECT  5.475 -0.115 5.545 0.410 ;
        RECT  5.165 -0.115 5.475 0.115 ;
        RECT  5.095 -0.115 5.165 0.255 ;
        RECT  4.790 -0.115 5.095 0.115 ;
        RECT  4.715 -0.115 4.790 0.305 ;
        RECT  4.055 -0.115 4.715 0.115 ;
        RECT  3.925 -0.115 4.055 0.250 ;
        RECT  3.670 -0.115 3.925 0.115 ;
        RECT  3.540 -0.115 3.670 0.250 ;
        RECT  2.775 -0.115 3.540 0.115 ;
        RECT  2.655 -0.115 2.775 0.190 ;
        RECT  2.025 -0.115 2.655 0.115 ;
        RECT  1.905 -0.115 2.025 0.190 ;
        RECT  1.145 -0.115 1.905 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.545 1.145 5.600 1.375 ;
        RECT  5.475 0.725 5.545 1.375 ;
        RECT  5.165 1.145 5.475 1.375 ;
        RECT  5.095 0.995 5.165 1.375 ;
        RECT  4.820 1.145 5.095 1.375 ;
        RECT  4.690 1.030 4.820 1.375 ;
        RECT  4.445 1.145 4.690 1.375 ;
        RECT  4.310 1.030 4.445 1.375 ;
        RECT  3.700 1.145 4.310 1.375 ;
        RECT  3.580 0.885 3.700 1.375 ;
        RECT  2.835 1.145 3.580 1.375 ;
        RECT  2.765 0.855 2.835 1.375 ;
        RECT  2.495 1.145 2.765 1.375 ;
        RECT  2.365 1.050 2.495 1.375 ;
        RECT  2.070 1.145 2.365 1.375 ;
        RECT  1.945 1.050 2.070 1.375 ;
        RECT  1.120 1.145 1.945 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.285 0.185 5.380 0.460 ;
        RECT  5.285 0.785 5.370 1.075 ;
        RECT  4.905 0.185 4.935 0.460 ;
        RECT  4.905 0.785 4.935 1.075 ;
        RECT  4.835 0.545 4.935 0.615 ;
        RECT  4.750 0.545 4.835 0.960 ;
        RECT  4.255 0.890 4.750 0.960 ;
        RECT  4.580 0.365 4.670 0.620 ;
        RECT  4.505 0.750 4.620 0.820 ;
        RECT  4.505 0.215 4.615 0.285 ;
        RECT  4.435 0.215 4.505 0.820 ;
        RECT  4.335 0.575 4.435 0.685 ;
        RECT  4.185 0.340 4.255 0.960 ;
        RECT  3.545 0.340 4.185 0.410 ;
        RECT  3.955 0.890 4.185 0.960 ;
        RECT  3.880 0.550 4.085 0.620 ;
        RECT  3.810 0.550 3.880 0.795 ;
        RECT  3.300 0.725 3.810 0.795 ;
        RECT  3.475 0.340 3.545 0.635 ;
        RECT  3.285 0.995 3.395 1.075 ;
        RECT  3.245 0.725 3.300 0.885 ;
        RECT  3.095 0.995 3.285 1.065 ;
        RECT  3.175 0.335 3.245 0.885 ;
        RECT  3.095 0.195 3.165 0.265 ;
        RECT  3.025 0.195 3.095 1.065 ;
        RECT  2.845 0.185 2.955 0.330 ;
        RECT  2.580 0.260 2.845 0.330 ;
        RECT  2.585 0.410 2.685 0.480 ;
        RECT  2.585 0.825 2.680 0.895 ;
        RECT  2.515 0.410 2.585 0.895 ;
        RECT  2.510 0.195 2.580 0.330 ;
        RECT  2.165 0.195 2.510 0.265 ;
        RECT  2.375 0.365 2.445 0.805 ;
        RECT  2.235 0.735 2.375 0.805 ;
        RECT  2.235 0.355 2.305 0.605 ;
        RECT  2.035 0.535 2.235 0.605 ;
        RECT  2.165 0.735 2.235 0.935 ;
        RECT  2.095 0.195 2.165 0.330 ;
        RECT  1.940 0.735 2.165 0.805 ;
        RECT  1.650 0.260 2.095 0.330 ;
        RECT  1.865 0.680 1.940 0.805 ;
        RECT  1.790 0.400 1.885 0.470 ;
        RECT  1.790 0.885 1.865 0.955 ;
        RECT  1.720 0.400 1.790 0.955 ;
        RECT  1.575 0.260 1.650 0.815 ;
        RECT  0.640 0.200 1.505 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.350 1.405 0.910 ;
        RECT  1.200 0.350 1.335 0.420 ;
        RECT  1.190 0.840 1.335 0.910 ;
        RECT  0.865 0.355 0.960 0.425 ;
        RECT  0.865 0.835 0.940 0.910 ;
        RECT  0.795 0.355 0.865 0.910 ;
        RECT  0.645 0.795 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.590 0.385 4.660 0.455 ;
        RECT  2.235 0.385 2.305 0.455 ;
    END
END SDFSNQD4BWP40

MACRO SDFSNQND0BWP40
    CLASS CORE ;
    FOREIGN SDFSNQND0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.055 ;
        RECT  4.635 0.185 4.655 0.300 ;
        RECT  4.635 0.915 4.655 1.055 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.180 ;
        RECT  4.150 -0.115 4.420 0.115 ;
        RECT  4.030 -0.115 4.150 0.210 ;
        RECT  3.730 -0.115 4.030 0.115 ;
        RECT  3.610 -0.115 3.730 0.210 ;
        RECT  2.805 -0.115 3.610 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.145 4.760 1.375 ;
        RECT  4.445 0.915 4.520 1.375 ;
        RECT  3.770 1.145 4.445 1.375 ;
        RECT  3.650 1.020 3.770 1.375 ;
        RECT  2.905 1.145 3.650 1.375 ;
        RECT  2.775 1.050 2.905 1.375 ;
        RECT  2.515 1.145 2.775 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.205 1.145 2.395 1.375 ;
        RECT  2.085 1.070 2.205 1.375 ;
        RECT  1.120 1.145 2.085 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.505 0.525 4.585 0.635 ;
        RECT  4.430 0.280 4.505 0.635 ;
        RECT  3.475 0.280 4.430 0.350 ;
        RECT  4.300 0.420 4.350 0.490 ;
        RECT  4.300 1.005 4.350 1.075 ;
        RECT  4.230 0.420 4.300 1.075 ;
        RECT  4.055 0.585 4.230 0.695 ;
        RECT  3.985 0.900 4.145 0.970 ;
        RECT  3.915 0.430 3.985 0.970 ;
        RECT  3.625 0.430 3.915 0.500 ;
        RECT  3.775 0.645 3.845 0.915 ;
        RECT  3.275 0.845 3.775 0.915 ;
        RECT  3.555 0.430 3.625 0.620 ;
        RECT  3.475 0.705 3.570 0.775 ;
        RECT  3.405 0.280 3.475 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.205 0.350 3.275 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.015 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.725 0.480 ;
        RECT  2.625 0.760 2.720 0.830 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.830 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.945 0.910 2.015 1.050 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.650 0.980 1.945 1.050 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.910 ;
        RECT  1.750 0.840 1.795 0.910 ;
        RECT  1.605 0.195 1.675 0.770 ;
        RECT  1.580 0.840 1.650 1.050 ;
        RECT  1.565 0.700 1.605 0.770 ;
        RECT  1.405 0.840 1.580 0.910 ;
        RECT  0.640 0.200 1.510 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.340 1.405 0.910 ;
        RECT  1.200 0.340 1.335 0.410 ;
        RECT  1.180 0.840 1.335 0.910 ;
        RECT  0.865 0.340 0.960 0.410 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.340 0.865 0.910 ;
        RECT  0.645 0.875 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFSNQND0BWP40

MACRO SDFSNQND1BWP40
    CLASS CORE ;
    FOREIGN SDFSNQND1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.655 0.185 4.725 1.075 ;
        RECT  4.635 0.185 4.655 0.465 ;
        RECT  4.635 0.685 4.655 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.540 -0.115 4.760 0.115 ;
        RECT  4.420 -0.115 4.540 0.180 ;
        RECT  4.150 -0.115 4.420 0.115 ;
        RECT  4.030 -0.115 4.150 0.210 ;
        RECT  3.730 -0.115 4.030 0.115 ;
        RECT  3.610 -0.115 3.730 0.210 ;
        RECT  2.805 -0.115 3.610 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.145 4.760 1.375 ;
        RECT  4.445 0.720 4.520 1.375 ;
        RECT  3.770 1.145 4.445 1.375 ;
        RECT  3.640 1.020 3.770 1.375 ;
        RECT  2.905 1.145 3.640 1.375 ;
        RECT  2.775 1.050 2.905 1.375 ;
        RECT  2.515 1.145 2.775 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.205 1.145 2.395 1.375 ;
        RECT  2.085 1.070 2.205 1.375 ;
        RECT  1.120 1.145 2.085 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.505 0.525 4.585 0.635 ;
        RECT  4.430 0.280 4.505 0.635 ;
        RECT  3.475 0.280 4.430 0.350 ;
        RECT  4.300 0.420 4.350 0.490 ;
        RECT  4.300 0.810 4.350 0.880 ;
        RECT  4.230 0.420 4.300 0.880 ;
        RECT  4.055 0.585 4.230 0.695 ;
        RECT  4.055 0.805 4.125 1.065 ;
        RECT  3.985 0.805 4.055 0.875 ;
        RECT  3.915 0.430 3.985 0.875 ;
        RECT  3.625 0.430 3.915 0.500 ;
        RECT  3.775 0.645 3.845 0.915 ;
        RECT  3.285 0.845 3.775 0.915 ;
        RECT  3.555 0.430 3.625 0.620 ;
        RECT  3.475 0.705 3.570 0.775 ;
        RECT  3.405 0.280 3.475 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.215 0.335 3.285 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.015 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.725 0.480 ;
        RECT  2.625 0.760 2.720 0.830 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.830 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.945 0.910 2.015 1.050 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.650 0.980 1.945 1.050 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.910 ;
        RECT  1.750 0.840 1.795 0.910 ;
        RECT  1.605 0.195 1.675 0.770 ;
        RECT  1.580 0.840 1.650 1.050 ;
        RECT  1.565 0.700 1.605 0.770 ;
        RECT  1.405 0.840 1.580 0.910 ;
        RECT  0.640 0.200 1.510 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.340 1.405 0.910 ;
        RECT  1.200 0.340 1.335 0.410 ;
        RECT  1.180 0.840 1.335 0.910 ;
        RECT  0.865 0.340 0.960 0.410 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.340 0.865 0.910 ;
        RECT  0.645 0.790 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFSNQND1BWP40

MACRO SDFSNQND2BWP40
    CLASS CORE ;
    FOREIGN SDFSNQND2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.900 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M2 ;
        RECT  2.080 0.665 4.360 0.735 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.660 0.370 4.725 0.795 ;
        RECT  4.655 0.195 4.660 1.075 ;
        RECT  4.585 0.195 4.655 0.445 ;
        RECT  4.585 0.720 4.655 1.075 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.490 2.910 0.905 ;
        RECT  2.670 0.605 2.835 0.675 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.115 4.900 0.115 ;
        RECT  4.775 -0.115 4.845 0.275 ;
        RECT  4.490 -0.115 4.775 0.115 ;
        RECT  4.370 -0.115 4.490 0.180 ;
        RECT  4.095 -0.115 4.370 0.115 ;
        RECT  3.975 -0.115 4.095 0.210 ;
        RECT  3.695 -0.115 3.975 0.115 ;
        RECT  3.555 -0.115 3.695 0.210 ;
        RECT  2.775 -0.115 3.555 0.115 ;
        RECT  2.655 -0.115 2.775 0.190 ;
        RECT  2.025 -0.115 2.655 0.115 ;
        RECT  1.905 -0.115 2.025 0.190 ;
        RECT  1.145 -0.115 1.905 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 1.145 4.900 1.375 ;
        RECT  4.775 0.865 4.845 1.375 ;
        RECT  4.465 1.145 4.775 1.375 ;
        RECT  4.395 0.865 4.465 1.375 ;
        RECT  3.720 1.145 4.395 1.375 ;
        RECT  3.640 0.985 3.720 1.375 ;
        RECT  2.835 1.145 3.640 1.375 ;
        RECT  2.765 0.985 2.835 1.375 ;
        RECT  2.495 1.145 2.765 1.375 ;
        RECT  2.365 1.050 2.495 1.375 ;
        RECT  2.070 1.145 2.365 1.375 ;
        RECT  1.945 1.050 2.070 1.375 ;
        RECT  1.120 1.145 1.945 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.495 0.525 4.585 0.635 ;
        RECT  4.420 0.280 4.495 0.635 ;
        RECT  3.455 0.280 4.420 0.350 ;
        RECT  4.210 0.620 4.340 0.790 ;
        RECT  4.080 0.865 4.300 0.935 ;
        RECT  4.080 0.420 4.295 0.495 ;
        RECT  3.940 1.005 4.115 1.075 ;
        RECT  4.010 0.420 4.080 0.935 ;
        RECT  3.870 0.430 3.940 1.075 ;
        RECT  3.595 0.430 3.870 0.500 ;
        RECT  3.720 0.635 3.790 0.915 ;
        RECT  3.245 0.845 3.720 0.915 ;
        RECT  3.525 0.430 3.595 0.625 ;
        RECT  3.455 0.705 3.545 0.775 ;
        RECT  3.385 0.280 3.455 0.775 ;
        RECT  3.285 0.995 3.395 1.075 ;
        RECT  3.095 0.995 3.285 1.065 ;
        RECT  3.175 0.335 3.245 0.915 ;
        RECT  3.095 0.195 3.165 0.265 ;
        RECT  3.025 0.195 3.095 1.065 ;
        RECT  2.845 0.185 2.955 0.330 ;
        RECT  2.580 0.260 2.845 0.330 ;
        RECT  2.585 0.410 2.685 0.480 ;
        RECT  2.585 0.865 2.680 0.935 ;
        RECT  2.515 0.410 2.585 0.935 ;
        RECT  2.510 0.195 2.580 0.330 ;
        RECT  2.165 0.195 2.510 0.265 ;
        RECT  2.375 0.365 2.445 0.935 ;
        RECT  2.030 0.865 2.375 0.935 ;
        RECT  2.100 0.620 2.230 0.790 ;
        RECT  2.095 0.195 2.165 0.330 ;
        RECT  1.650 0.260 2.095 0.330 ;
        RECT  1.960 0.695 2.030 0.935 ;
        RECT  1.905 0.695 1.960 0.805 ;
        RECT  1.790 0.400 1.885 0.470 ;
        RECT  1.790 0.865 1.865 0.935 ;
        RECT  1.720 0.400 1.790 0.935 ;
        RECT  1.575 0.260 1.650 0.815 ;
        RECT  0.640 0.200 1.505 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.340 1.405 0.910 ;
        RECT  1.200 0.340 1.335 0.410 ;
        RECT  1.180 0.840 1.335 0.910 ;
        RECT  0.865 0.340 0.960 0.410 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.340 0.865 0.910 ;
        RECT  0.645 0.790 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
        LAYER VIA1 ;
        RECT  4.240 0.665 4.310 0.735 ;
        RECT  2.130 0.665 2.200 0.735 ;
    END
END SDFSNQND2BWP40

MACRO SDFSNQND4BWP40
    CLASS CORE ;
    FOREIGN SDFSNQND4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.395 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.027600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.035 0.495 0.195 0.765 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.019200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.355 2.205 0.625 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.425 0.190 5.520 0.440 ;
        RECT  5.425 0.745 5.520 1.005 ;
        RECT  5.355 0.355 5.425 0.440 ;
        RECT  5.355 0.745 5.425 0.830 ;
        RECT  5.145 0.355 5.355 0.830 ;
        RECT  5.120 0.355 5.145 0.475 ;
        RECT  5.120 0.710 5.145 0.830 ;
        RECT  5.050 0.205 5.120 0.475 ;
        RECT  5.050 0.710 5.120 1.020 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.026400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.085 0.765 ;
        RECT  0.945 0.495 1.015 0.640 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 0.465 2.910 0.765 ;
        RECT  2.710 0.605 2.835 0.675 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.115 5.740 0.115 ;
        RECT  5.610 -0.115 5.690 0.430 ;
        RECT  5.305 -0.115 5.610 0.115 ;
        RECT  5.235 -0.115 5.305 0.270 ;
        RECT  4.950 -0.115 5.235 0.115 ;
        RECT  4.830 -0.115 4.950 0.210 ;
        RECT  4.560 -0.115 4.830 0.115 ;
        RECT  4.440 -0.115 4.560 0.210 ;
        RECT  4.130 -0.115 4.440 0.115 ;
        RECT  4.005 -0.115 4.130 0.210 ;
        RECT  3.760 -0.115 4.005 0.115 ;
        RECT  3.635 -0.115 3.760 0.210 ;
        RECT  2.805 -0.115 3.635 0.115 ;
        RECT  2.695 -0.115 2.805 0.195 ;
        RECT  2.095 -0.115 2.695 0.115 ;
        RECT  1.975 -0.115 2.095 0.125 ;
        RECT  1.145 -0.115 1.975 0.115 ;
        RECT  1.015 -0.115 1.145 0.130 ;
        RECT  0.340 -0.115 1.015 0.115 ;
        RECT  0.220 -0.115 0.340 0.280 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 1.145 5.740 1.375 ;
        RECT  5.610 0.705 5.690 1.375 ;
        RECT  5.325 1.145 5.610 1.375 ;
        RECT  5.215 0.905 5.325 1.375 ;
        RECT  4.930 1.145 5.215 1.375 ;
        RECT  4.855 0.720 4.930 1.375 ;
        RECT  4.165 1.145 4.855 1.375 ;
        RECT  4.035 1.005 4.165 1.375 ;
        RECT  3.760 1.145 4.035 1.375 ;
        RECT  3.620 1.050 3.760 1.375 ;
        RECT  2.905 1.145 3.620 1.375 ;
        RECT  2.775 1.050 2.905 1.375 ;
        RECT  2.515 1.145 2.775 1.375 ;
        RECT  2.395 1.050 2.515 1.375 ;
        RECT  2.205 1.145 2.395 1.375 ;
        RECT  2.085 1.070 2.205 1.375 ;
        RECT  1.120 1.145 2.085 1.375 ;
        RECT  1.000 1.120 1.120 1.375 ;
        RECT  0.340 1.145 1.000 1.375 ;
        RECT  0.220 0.985 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.425 0.190 5.520 0.440 ;
        RECT  5.425 0.745 5.520 1.005 ;
        RECT  5.050 0.205 5.075 0.475 ;
        RECT  5.050 0.710 5.075 1.020 ;
        RECT  4.915 0.545 5.065 0.620 ;
        RECT  4.840 0.280 4.915 0.620 ;
        RECT  3.950 0.280 4.840 0.350 ;
        RECT  4.670 0.420 4.760 0.495 ;
        RECT  4.670 0.815 4.760 0.885 ;
        RECT  4.600 0.420 4.670 0.885 ;
        RECT  4.435 0.585 4.600 0.695 ;
        RECT  4.460 0.800 4.530 1.065 ;
        RECT  4.355 0.800 4.460 0.870 ;
        RECT  4.285 0.425 4.355 0.870 ;
        RECT  4.235 0.425 4.285 0.565 ;
        RECT  3.765 0.495 4.235 0.565 ;
        RECT  4.145 0.645 4.215 0.915 ;
        RECT  3.285 0.845 4.145 0.915 ;
        RECT  3.830 0.280 3.950 0.400 ;
        RECT  3.515 0.705 3.950 0.775 ;
        RECT  3.515 0.280 3.830 0.350 ;
        RECT  3.655 0.495 3.765 0.625 ;
        RECT  3.445 0.280 3.515 0.775 ;
        RECT  3.360 0.995 3.470 1.075 ;
        RECT  3.135 0.995 3.360 1.065 ;
        RECT  3.215 0.335 3.285 0.915 ;
        RECT  3.135 0.195 3.200 0.265 ;
        RECT  3.065 0.195 3.135 1.065 ;
        RECT  2.015 0.910 3.065 0.980 ;
        RECT  2.885 0.185 2.995 0.340 ;
        RECT  2.625 0.270 2.885 0.340 ;
        RECT  2.625 0.410 2.725 0.480 ;
        RECT  2.625 0.760 2.720 0.830 ;
        RECT  2.555 0.195 2.625 0.340 ;
        RECT  2.555 0.410 2.625 0.830 ;
        RECT  2.345 0.195 2.555 0.265 ;
        RECT  2.415 0.345 2.485 0.830 ;
        RECT  2.010 0.760 2.415 0.830 ;
        RECT  2.275 0.195 2.345 0.610 ;
        RECT  1.675 0.195 2.275 0.265 ;
        RECT  1.945 0.910 2.015 1.050 ;
        RECT  1.940 0.610 2.010 0.830 ;
        RECT  1.650 0.980 1.945 1.050 ;
        RECT  1.870 0.335 1.915 0.405 ;
        RECT  1.795 0.335 1.870 0.910 ;
        RECT  1.750 0.840 1.795 0.910 ;
        RECT  1.605 0.195 1.675 0.770 ;
        RECT  1.580 0.840 1.650 1.050 ;
        RECT  1.565 0.700 1.605 0.770 ;
        RECT  1.405 0.840 1.580 0.910 ;
        RECT  0.640 0.200 1.510 0.270 ;
        RECT  0.715 0.980 1.490 1.050 ;
        RECT  1.335 0.340 1.405 0.910 ;
        RECT  1.200 0.340 1.335 0.410 ;
        RECT  1.180 0.840 1.335 0.910 ;
        RECT  0.865 0.340 0.960 0.410 ;
        RECT  0.865 0.840 0.940 0.910 ;
        RECT  0.795 0.340 0.865 0.910 ;
        RECT  0.645 0.790 0.715 1.050 ;
        RECT  0.555 0.530 0.615 0.650 ;
        RECT  0.485 0.350 0.555 0.915 ;
        RECT  0.125 0.350 0.485 0.420 ;
        RECT  0.125 0.845 0.485 0.915 ;
        RECT  0.055 0.300 0.125 0.420 ;
        RECT  0.055 0.845 0.125 1.075 ;
    END
END SDFSNQND4BWP40

MACRO SEDFCNQD0BWP40
    CLASS CORE ;
    FOREIGN SEDFCNQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.195 5.985 1.065 ;
        RECT  5.895 0.195 5.915 0.315 ;
        RECT  5.895 0.935 5.915 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.021400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.014600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.355 3.645 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.805 -0.115 6.020 0.115 ;
        RECT  5.675 -0.115 5.805 0.160 ;
        RECT  5.435 -0.115 5.675 0.115 ;
        RECT  5.305 -0.115 5.435 0.160 ;
        RECT  4.345 -0.115 5.305 0.115 ;
        RECT  4.225 -0.115 4.345 0.345 ;
        RECT  3.515 -0.115 4.225 0.115 ;
        RECT  3.395 -0.115 3.515 0.125 ;
        RECT  2.520 -0.115 3.395 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.780 1.145 6.020 1.375 ;
        RECT  5.705 1.005 5.780 1.375 ;
        RECT  5.215 1.145 5.705 1.375 ;
        RECT  5.145 1.005 5.215 1.375 ;
        RECT  4.385 1.145 5.145 1.375 ;
        RECT  4.265 0.890 4.385 1.375 ;
        RECT  3.995 1.145 4.265 1.375 ;
        RECT  3.875 1.015 3.995 1.375 ;
        RECT  3.560 1.145 3.875 1.375 ;
        RECT  3.440 1.030 3.560 1.375 ;
        RECT  2.395 1.145 3.440 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.825 0.520 5.840 0.640 ;
        RECT  5.755 0.240 5.825 0.925 ;
        RECT  5.035 0.240 5.755 0.310 ;
        RECT  5.055 0.855 5.755 0.925 ;
        RECT  5.615 0.380 5.685 0.775 ;
        RECT  5.210 0.380 5.615 0.450 ;
        RECT  5.490 0.695 5.615 0.775 ;
        RECT  5.405 0.540 5.505 0.615 ;
        RECT  5.330 0.540 5.405 0.760 ;
        RECT  4.795 0.690 5.330 0.760 ;
        RECT  5.140 0.380 5.210 0.600 ;
        RECT  4.895 0.530 5.140 0.600 ;
        RECT  4.930 0.830 5.055 0.925 ;
        RECT  4.965 0.240 5.035 0.425 ;
        RECT  4.615 0.995 4.935 1.065 ;
        RECT  4.825 0.200 4.895 0.600 ;
        RECT  4.755 0.690 4.795 0.890 ;
        RECT  4.685 0.350 4.755 0.890 ;
        RECT  4.545 0.425 4.615 1.065 ;
        RECT  4.135 0.425 4.545 0.495 ;
        RECT  4.175 0.740 4.545 0.810 ;
        RECT  3.945 0.565 4.465 0.650 ;
        RECT  4.105 0.740 4.175 0.900 ;
        RECT  4.055 0.195 4.135 0.495 ;
        RECT  3.285 0.195 4.055 0.265 ;
        RECT  3.795 0.335 3.955 0.405 ;
        RECT  3.875 0.565 3.945 0.925 ;
        RECT  3.165 0.855 3.875 0.925 ;
        RECT  3.725 0.335 3.795 0.765 ;
        RECT  3.455 0.695 3.725 0.765 ;
        RECT  3.385 0.660 3.455 0.765 ;
        RECT  3.315 0.360 3.360 0.430 ;
        RECT  3.235 0.360 3.315 0.775 ;
        RECT  3.165 0.190 3.285 0.265 ;
        RECT  3.025 0.995 3.215 1.065 ;
        RECT  3.105 0.685 3.165 0.925 ;
        RECT  3.105 0.335 3.150 0.410 ;
        RECT  3.095 0.335 3.105 0.925 ;
        RECT  3.030 0.335 3.095 0.760 ;
        RECT  2.965 0.690 3.030 0.760 ;
        RECT  2.955 0.845 3.025 1.065 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.955 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.675 0.985 2.835 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.675 1.055 ;
        RECT  2.255 0.200 2.335 0.345 ;
        RECT  1.925 0.200 2.255 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.720 ;
        RECT  1.680 0.640 2.045 0.720 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.675 0.640 1.680 0.765 ;
        RECT  1.600 0.505 1.675 0.765 ;
        RECT  0.455 0.205 1.610 0.275 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.100 0.685 1.220 0.765 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  4.825 0.245 4.895 0.315 ;
        RECT  2.260 0.245 2.330 0.315 ;
        LAYER M2 ;
        RECT  2.210 0.245 4.945 0.315 ;
    END
END SEDFCNQD0BWP40

MACRO SEDFCNQD1BWP40
    CLASS CORE ;
    FOREIGN SEDFCNQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.020 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.195 5.985 1.065 ;
        RECT  5.895 0.195 5.915 0.475 ;
        RECT  5.895 0.730 5.915 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.040400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.355 3.645 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.805 -0.115 6.020 0.115 ;
        RECT  5.675 -0.115 5.805 0.160 ;
        RECT  5.435 -0.115 5.675 0.115 ;
        RECT  5.305 -0.115 5.435 0.160 ;
        RECT  4.345 -0.115 5.305 0.115 ;
        RECT  4.225 -0.115 4.345 0.345 ;
        RECT  3.515 -0.115 4.225 0.115 ;
        RECT  3.395 -0.115 3.515 0.125 ;
        RECT  2.520 -0.115 3.395 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.780 1.145 6.020 1.375 ;
        RECT  5.705 1.005 5.780 1.375 ;
        RECT  5.215 1.145 5.705 1.375 ;
        RECT  5.145 1.005 5.215 1.375 ;
        RECT  4.385 1.145 5.145 1.375 ;
        RECT  4.265 0.890 4.385 1.375 ;
        RECT  3.995 1.145 4.265 1.375 ;
        RECT  3.875 1.015 3.995 1.375 ;
        RECT  3.560 1.145 3.875 1.375 ;
        RECT  3.440 1.030 3.560 1.375 ;
        RECT  2.395 1.145 3.440 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.825 0.520 5.840 0.640 ;
        RECT  5.755 0.240 5.825 0.925 ;
        RECT  5.035 0.240 5.755 0.310 ;
        RECT  5.055 0.855 5.755 0.925 ;
        RECT  5.615 0.380 5.685 0.775 ;
        RECT  5.210 0.380 5.615 0.450 ;
        RECT  5.490 0.695 5.615 0.775 ;
        RECT  5.405 0.540 5.505 0.615 ;
        RECT  5.330 0.540 5.405 0.760 ;
        RECT  4.795 0.690 5.330 0.760 ;
        RECT  5.140 0.380 5.210 0.600 ;
        RECT  4.895 0.530 5.140 0.600 ;
        RECT  4.930 0.830 5.055 0.925 ;
        RECT  4.965 0.240 5.035 0.425 ;
        RECT  4.615 0.995 4.935 1.065 ;
        RECT  4.825 0.200 4.895 0.600 ;
        RECT  4.755 0.690 4.795 0.890 ;
        RECT  4.685 0.350 4.755 0.890 ;
        RECT  4.545 0.425 4.615 1.065 ;
        RECT  4.135 0.425 4.545 0.495 ;
        RECT  4.175 0.740 4.545 0.810 ;
        RECT  3.945 0.565 4.465 0.650 ;
        RECT  4.105 0.740 4.175 0.955 ;
        RECT  4.055 0.195 4.135 0.495 ;
        RECT  3.285 0.195 4.055 0.265 ;
        RECT  3.795 0.335 3.955 0.405 ;
        RECT  3.875 0.565 3.945 0.925 ;
        RECT  3.165 0.855 3.875 0.925 ;
        RECT  3.725 0.335 3.795 0.765 ;
        RECT  3.455 0.695 3.725 0.765 ;
        RECT  3.385 0.660 3.455 0.765 ;
        RECT  3.305 0.360 3.360 0.430 ;
        RECT  3.305 0.655 3.315 0.775 ;
        RECT  3.235 0.360 3.305 0.775 ;
        RECT  3.165 0.190 3.285 0.265 ;
        RECT  3.025 0.995 3.215 1.065 ;
        RECT  3.105 0.685 3.165 0.925 ;
        RECT  3.105 0.335 3.150 0.410 ;
        RECT  3.095 0.335 3.105 0.925 ;
        RECT  3.030 0.335 3.095 0.760 ;
        RECT  2.965 0.690 3.030 0.760 ;
        RECT  2.955 0.845 3.025 1.065 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.955 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.675 0.985 2.835 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.675 1.055 ;
        RECT  2.255 0.200 2.335 0.345 ;
        RECT  1.925 0.200 2.255 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.720 ;
        RECT  1.680 0.640 2.045 0.720 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.675 0.640 1.680 0.765 ;
        RECT  1.600 0.505 1.675 0.765 ;
        RECT  0.455 0.205 1.610 0.275 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.100 0.685 1.220 0.765 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  4.825 0.245 4.895 0.315 ;
        RECT  2.260 0.245 2.330 0.315 ;
        LAYER M2 ;
        RECT  2.210 0.245 4.945 0.315 ;
    END
END SEDFCNQD1BWP40

MACRO SEDFCNQD2BWP40
    CLASS CORE ;
    FOREIGN SEDFCNQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.300 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.148200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.195 5.985 1.065 ;
        RECT  5.895 0.195 5.915 0.475 ;
        RECT  5.895 0.730 5.915 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.040400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.355 3.645 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.215 -0.115 6.300 0.115 ;
        RECT  6.140 -0.115 6.215 0.490 ;
        RECT  5.805 -0.115 6.140 0.115 ;
        RECT  5.675 -0.115 5.805 0.160 ;
        RECT  5.435 -0.115 5.675 0.115 ;
        RECT  5.305 -0.115 5.435 0.160 ;
        RECT  4.345 -0.115 5.305 0.115 ;
        RECT  4.225 -0.115 4.345 0.345 ;
        RECT  3.515 -0.115 4.225 0.115 ;
        RECT  3.395 -0.115 3.515 0.125 ;
        RECT  2.520 -0.115 3.395 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.215 1.145 6.300 1.375 ;
        RECT  6.140 0.670 6.215 1.375 ;
        RECT  5.780 1.145 6.140 1.375 ;
        RECT  5.705 1.005 5.780 1.375 ;
        RECT  5.215 1.145 5.705 1.375 ;
        RECT  5.145 1.005 5.215 1.375 ;
        RECT  4.385 1.145 5.145 1.375 ;
        RECT  4.265 0.890 4.385 1.375 ;
        RECT  3.995 1.145 4.265 1.375 ;
        RECT  3.875 1.015 3.995 1.375 ;
        RECT  3.560 1.145 3.875 1.375 ;
        RECT  3.440 1.030 3.560 1.375 ;
        RECT  2.395 1.145 3.440 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.825 0.520 5.840 0.640 ;
        RECT  5.755 0.240 5.825 0.925 ;
        RECT  5.035 0.240 5.755 0.310 ;
        RECT  5.430 0.855 5.755 0.925 ;
        RECT  5.615 0.380 5.685 0.775 ;
        RECT  5.210 0.380 5.615 0.450 ;
        RECT  5.490 0.695 5.615 0.775 ;
        RECT  5.405 0.540 5.505 0.615 ;
        RECT  5.310 0.855 5.430 1.065 ;
        RECT  5.330 0.540 5.405 0.760 ;
        RECT  4.795 0.690 5.330 0.760 ;
        RECT  5.055 0.855 5.310 0.925 ;
        RECT  5.140 0.380 5.210 0.600 ;
        RECT  4.895 0.530 5.140 0.600 ;
        RECT  4.930 0.830 5.055 0.925 ;
        RECT  4.965 0.240 5.035 0.425 ;
        RECT  4.615 0.995 4.935 1.065 ;
        RECT  4.825 0.200 4.895 0.600 ;
        RECT  4.755 0.690 4.795 0.890 ;
        RECT  4.685 0.350 4.755 0.890 ;
        RECT  4.545 0.425 4.615 1.065 ;
        RECT  4.135 0.425 4.545 0.495 ;
        RECT  4.175 0.740 4.545 0.810 ;
        RECT  3.945 0.565 4.465 0.650 ;
        RECT  4.105 0.740 4.175 0.955 ;
        RECT  4.055 0.195 4.135 0.495 ;
        RECT  3.285 0.195 4.055 0.265 ;
        RECT  3.795 0.335 3.955 0.405 ;
        RECT  3.875 0.565 3.945 0.925 ;
        RECT  3.165 0.855 3.875 0.925 ;
        RECT  3.725 0.335 3.795 0.765 ;
        RECT  3.455 0.695 3.725 0.765 ;
        RECT  3.385 0.660 3.455 0.765 ;
        RECT  3.305 0.360 3.360 0.430 ;
        RECT  3.305 0.655 3.315 0.775 ;
        RECT  3.235 0.360 3.305 0.775 ;
        RECT  3.165 0.190 3.285 0.265 ;
        RECT  3.025 0.995 3.215 1.065 ;
        RECT  3.105 0.685 3.165 0.925 ;
        RECT  3.105 0.335 3.150 0.410 ;
        RECT  3.095 0.335 3.105 0.925 ;
        RECT  3.030 0.335 3.095 0.760 ;
        RECT  2.965 0.690 3.030 0.760 ;
        RECT  2.955 0.845 3.025 1.065 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.955 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.675 0.985 2.835 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.675 1.055 ;
        RECT  2.255 0.200 2.335 0.345 ;
        RECT  1.925 0.200 2.255 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.720 ;
        RECT  1.680 0.640 2.045 0.720 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.675 0.640 1.680 0.765 ;
        RECT  1.600 0.505 1.675 0.765 ;
        RECT  0.455 0.205 1.610 0.275 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.100 0.685 1.220 0.765 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  4.825 0.245 4.895 0.315 ;
        RECT  2.260 0.245 2.330 0.315 ;
        LAYER M2 ;
        RECT  2.210 0.245 4.945 0.315 ;
    END
END SEDFCNQD2BWP40

MACRO SEDFCNQD4BWP40
    CLASS CORE ;
    FOREIGN SEDFCNQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.237000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.685 0.195 6.780 0.475 ;
        RECT  6.685 0.710 6.780 1.010 ;
        RECT  6.615 0.355 6.685 0.475 ;
        RECT  6.615 0.710 6.685 0.830 ;
        RECT  6.405 0.355 6.615 0.830 ;
        RECT  6.380 0.355 6.405 0.475 ;
        RECT  6.380 0.710 6.405 0.830 ;
        RECT  6.310 0.195 6.380 0.475 ;
        RECT  6.310 0.710 6.380 1.010 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.019800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.052800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.355 3.645 0.625 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.945 -0.115 7.000 0.115 ;
        RECT  6.870 -0.115 6.945 0.450 ;
        RECT  6.590 -0.115 6.870 0.115 ;
        RECT  6.465 -0.115 6.590 0.235 ;
        RECT  6.215 -0.115 6.465 0.115 ;
        RECT  6.085 -0.115 6.215 0.160 ;
        RECT  5.405 -0.115 6.085 0.115 ;
        RECT  5.305 -0.115 5.405 0.270 ;
        RECT  4.345 -0.115 5.305 0.115 ;
        RECT  4.225 -0.115 4.345 0.345 ;
        RECT  3.515 -0.115 4.225 0.115 ;
        RECT  3.395 -0.115 3.515 0.125 ;
        RECT  2.520 -0.115 3.395 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.950 1.145 7.000 1.375 ;
        RECT  6.875 0.700 6.950 1.375 ;
        RECT  6.590 1.145 6.875 1.375 ;
        RECT  6.465 0.905 6.590 1.375 ;
        RECT  6.215 1.145 6.465 1.375 ;
        RECT  6.090 1.025 6.215 1.375 ;
        RECT  5.625 1.145 6.090 1.375 ;
        RECT  5.500 1.025 5.625 1.375 ;
        RECT  5.240 1.145 5.500 1.375 ;
        RECT  5.120 1.025 5.240 1.375 ;
        RECT  4.385 1.145 5.120 1.375 ;
        RECT  4.265 0.890 4.385 1.375 ;
        RECT  3.995 1.145 4.265 1.375 ;
        RECT  3.875 1.015 3.995 1.375 ;
        RECT  3.560 1.145 3.875 1.375 ;
        RECT  3.440 1.030 3.560 1.375 ;
        RECT  2.395 1.145 3.440 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.685 0.195 6.780 0.475 ;
        RECT  6.685 0.710 6.780 1.010 ;
        RECT  6.310 0.195 6.335 0.475 ;
        RECT  6.310 0.710 6.335 1.010 ;
        RECT  6.240 0.545 6.325 0.615 ;
        RECT  6.170 0.240 6.240 0.930 ;
        RECT  5.545 0.240 6.170 0.310 ;
        RECT  5.820 0.860 6.170 0.930 ;
        RECT  6.030 0.380 6.100 0.780 ;
        RECT  5.685 0.380 6.030 0.450 ;
        RECT  5.900 0.710 6.030 0.780 ;
        RECT  5.830 0.530 5.950 0.630 ;
        RECT  5.755 0.530 5.830 0.760 ;
        RECT  5.700 0.860 5.820 1.060 ;
        RECT  4.795 0.690 5.755 0.760 ;
        RECT  5.430 0.860 5.700 0.930 ;
        RECT  5.615 0.380 5.685 0.600 ;
        RECT  4.895 0.530 5.615 0.600 ;
        RECT  5.475 0.240 5.545 0.425 ;
        RECT  5.035 0.355 5.475 0.425 ;
        RECT  5.310 0.860 5.430 1.060 ;
        RECT  5.085 0.860 5.310 0.930 ;
        RECT  5.045 0.830 5.085 0.930 ;
        RECT  4.930 0.830 5.045 0.925 ;
        RECT  4.965 0.305 5.035 0.425 ;
        RECT  4.615 0.995 4.935 1.065 ;
        RECT  4.825 0.200 4.895 0.600 ;
        RECT  4.755 0.690 4.795 0.890 ;
        RECT  4.685 0.350 4.755 0.890 ;
        RECT  4.545 0.425 4.615 1.065 ;
        RECT  4.135 0.425 4.545 0.495 ;
        RECT  4.175 0.740 4.545 0.810 ;
        RECT  3.945 0.565 4.465 0.650 ;
        RECT  4.105 0.740 4.175 0.955 ;
        RECT  4.055 0.195 4.135 0.495 ;
        RECT  3.285 0.195 4.055 0.265 ;
        RECT  3.795 0.335 3.955 0.405 ;
        RECT  3.875 0.565 3.945 0.925 ;
        RECT  3.165 0.855 3.875 0.925 ;
        RECT  3.725 0.335 3.795 0.765 ;
        RECT  3.455 0.695 3.725 0.765 ;
        RECT  3.385 0.660 3.455 0.765 ;
        RECT  3.305 0.360 3.360 0.430 ;
        RECT  3.305 0.655 3.315 0.775 ;
        RECT  3.235 0.360 3.305 0.775 ;
        RECT  3.165 0.190 3.285 0.265 ;
        RECT  3.025 0.995 3.215 1.065 ;
        RECT  3.105 0.685 3.165 0.925 ;
        RECT  3.105 0.335 3.150 0.410 ;
        RECT  3.095 0.335 3.105 0.925 ;
        RECT  3.030 0.335 3.095 0.760 ;
        RECT  2.965 0.690 3.030 0.760 ;
        RECT  2.955 0.845 3.025 1.065 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.955 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.675 0.985 2.835 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.675 1.055 ;
        RECT  2.255 0.200 2.335 0.345 ;
        RECT  1.925 0.200 2.255 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.720 ;
        RECT  1.680 0.640 2.045 0.720 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.675 0.640 1.680 0.765 ;
        RECT  1.600 0.505 1.675 0.765 ;
        RECT  0.455 0.205 1.610 0.275 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.100 0.685 1.220 0.765 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  4.825 0.245 4.895 0.315 ;
        RECT  2.260 0.245 2.330 0.315 ;
        LAYER M2 ;
        RECT  2.210 0.245 4.945 0.315 ;
    END
END SEDFCNQD4BWP40

MACRO SEDFQD0BWP40
    CLASS CORE ;
    FOREIGN SEDFQD0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.023400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.045 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.021400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 -0.115 5.600 0.115 ;
        RECT  5.285 -0.115 5.355 0.315 ;
        RECT  4.985 -0.115 5.285 0.115 ;
        RECT  4.915 -0.115 4.985 0.285 ;
        RECT  4.170 -0.115 4.915 0.115 ;
        RECT  4.030 -0.115 4.170 0.130 ;
        RECT  3.550 -0.115 4.030 0.115 ;
        RECT  3.430 -0.115 3.550 0.125 ;
        RECT  2.520 -0.115 3.430 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 1.145 5.600 1.375 ;
        RECT  5.285 0.895 5.355 1.375 ;
        RECT  4.980 1.145 5.285 1.375 ;
        RECT  4.850 1.130 4.980 1.375 ;
        RECT  4.150 1.145 4.850 1.375 ;
        RECT  4.030 0.970 4.150 1.375 ;
        RECT  3.545 1.145 4.030 1.375 ;
        RECT  3.425 1.000 3.545 1.375 ;
        RECT  2.395 1.145 3.425 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.245 0.395 5.315 0.810 ;
        RECT  5.200 0.395 5.245 0.465 ;
        RECT  5.175 0.740 5.245 0.810 ;
        RECT  5.080 0.190 5.200 0.465 ;
        RECT  5.105 0.740 5.175 0.900 ;
        RECT  5.025 0.545 5.155 0.615 ;
        RECT  4.865 0.395 5.080 0.465 ;
        RECT  4.955 0.545 5.025 0.920 ;
        RECT  4.550 0.850 4.955 0.920 ;
        RECT  4.775 0.395 4.865 0.600 ;
        RECT  4.400 0.995 4.730 1.065 ;
        RECT  4.480 0.235 4.550 0.920 ;
        RECT  4.330 0.200 4.400 1.065 ;
        RECT  3.265 0.200 4.330 0.270 ;
        RECT  4.315 0.785 4.330 1.065 ;
        RECT  3.935 0.785 4.315 0.855 ;
        RECT  3.800 0.540 4.235 0.660 ;
        RECT  3.860 0.785 3.935 0.930 ;
        RECT  3.730 0.340 3.760 0.420 ;
        RECT  3.660 0.340 3.730 0.930 ;
        RECT  3.640 0.340 3.660 0.600 ;
        RECT  3.385 0.485 3.640 0.600 ;
        RECT  3.500 0.670 3.590 0.930 ;
        RECT  3.160 0.860 3.500 0.930 ;
        RECT  3.315 0.350 3.340 0.430 ;
        RECT  3.230 0.350 3.315 0.780 ;
        RECT  3.145 0.190 3.265 0.270 ;
        RECT  3.020 1.000 3.215 1.070 ;
        RECT  3.110 0.690 3.160 0.930 ;
        RECT  3.110 0.350 3.150 0.420 ;
        RECT  3.090 0.350 3.110 0.930 ;
        RECT  3.030 0.350 3.090 0.760 ;
        RECT  2.980 0.690 3.030 0.760 ;
        RECT  2.950 0.845 3.020 1.070 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.950 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.695 0.985 2.855 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.695 1.055 ;
        RECT  2.275 0.200 2.345 0.345 ;
        RECT  1.925 0.200 2.275 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.755 ;
        RECT  1.675 0.685 2.045 0.755 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.650 0.505 1.675 0.755 ;
        RECT  1.600 0.505 1.650 0.765 ;
        RECT  1.085 0.195 1.610 0.265 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.095 0.685 1.220 0.765 ;
        RECT  1.015 0.195 1.085 0.275 ;
        RECT  0.455 0.205 1.015 0.275 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  5.110 0.245 5.180 0.315 ;
        RECT  2.275 0.245 2.345 0.315 ;
        LAYER M2 ;
        RECT  2.225 0.245 5.230 0.315 ;
    END
END SEDFQD0BWP40

MACRO SEDFQD1BWP40
    CLASS CORE ;
    FOREIGN SEDFQD1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.065 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 -0.115 5.600 0.115 ;
        RECT  5.285 -0.115 5.355 0.315 ;
        RECT  4.985 -0.115 5.285 0.115 ;
        RECT  4.915 -0.115 4.985 0.300 ;
        RECT  4.170 -0.115 4.915 0.115 ;
        RECT  4.030 -0.115 4.170 0.130 ;
        RECT  3.540 -0.115 4.030 0.115 ;
        RECT  3.420 -0.115 3.540 0.125 ;
        RECT  2.520 -0.115 3.420 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 1.145 5.600 1.375 ;
        RECT  5.285 0.895 5.355 1.375 ;
        RECT  4.980 1.145 5.285 1.375 ;
        RECT  4.850 1.130 4.980 1.375 ;
        RECT  4.150 1.145 4.850 1.375 ;
        RECT  4.030 0.890 4.150 1.375 ;
        RECT  3.545 1.145 4.030 1.375 ;
        RECT  3.425 1.000 3.545 1.375 ;
        RECT  2.395 1.145 3.425 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.245 0.395 5.315 0.810 ;
        RECT  5.185 0.395 5.245 0.465 ;
        RECT  5.175 0.740 5.245 0.810 ;
        RECT  5.095 0.195 5.185 0.465 ;
        RECT  5.105 0.740 5.175 1.025 ;
        RECT  5.025 0.545 5.155 0.615 ;
        RECT  4.865 0.395 5.095 0.465 ;
        RECT  4.955 0.545 5.025 0.920 ;
        RECT  4.550 0.850 4.955 0.920 ;
        RECT  4.775 0.395 4.865 0.600 ;
        RECT  4.400 0.995 4.730 1.065 ;
        RECT  4.480 0.350 4.550 0.920 ;
        RECT  4.330 0.200 4.400 1.065 ;
        RECT  3.265 0.200 4.330 0.270 ;
        RECT  4.315 0.740 4.330 1.065 ;
        RECT  3.935 0.740 4.315 0.810 ;
        RECT  3.800 0.540 4.235 0.660 ;
        RECT  3.860 0.740 3.935 0.930 ;
        RECT  3.730 0.340 3.760 0.420 ;
        RECT  3.660 0.340 3.730 0.930 ;
        RECT  3.640 0.340 3.660 0.600 ;
        RECT  3.385 0.485 3.640 0.600 ;
        RECT  3.500 0.670 3.590 0.930 ;
        RECT  3.160 0.860 3.500 0.930 ;
        RECT  3.315 0.350 3.340 0.430 ;
        RECT  3.230 0.350 3.315 0.780 ;
        RECT  3.145 0.190 3.265 0.270 ;
        RECT  3.020 1.000 3.215 1.070 ;
        RECT  3.110 0.690 3.160 0.930 ;
        RECT  3.110 0.350 3.150 0.420 ;
        RECT  3.090 0.350 3.110 0.930 ;
        RECT  3.030 0.350 3.090 0.760 ;
        RECT  2.980 0.690 3.030 0.760 ;
        RECT  2.950 0.845 3.020 1.070 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.950 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.695 0.985 2.855 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.695 1.055 ;
        RECT  2.275 0.200 2.345 0.345 ;
        RECT  1.925 0.200 2.275 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.755 ;
        RECT  1.675 0.685 2.045 0.755 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.650 0.505 1.675 0.755 ;
        RECT  1.600 0.505 1.650 0.765 ;
        RECT  1.085 0.195 1.610 0.265 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.095 0.685 1.220 0.765 ;
        RECT  1.015 0.195 1.085 0.275 ;
        RECT  0.455 0.205 1.015 0.275 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  5.110 0.245 5.180 0.315 ;
        RECT  2.275 0.245 2.345 0.315 ;
        LAYER M2 ;
        RECT  2.225 0.245 5.230 0.315 ;
    END
END SEDFQD1BWP40

MACRO SEDFQD2BWP40
    CLASS CORE ;
    FOREIGN SEDFQD2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.164000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.195 5.565 1.070 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 -0.115 5.880 0.115 ;
        RECT  5.730 -0.115 5.810 0.475 ;
        RECT  5.355 -0.115 5.730 0.115 ;
        RECT  5.285 -0.115 5.355 0.315 ;
        RECT  4.985 -0.115 5.285 0.115 ;
        RECT  4.915 -0.115 4.985 0.270 ;
        RECT  4.170 -0.115 4.915 0.115 ;
        RECT  4.030 -0.115 4.170 0.130 ;
        RECT  3.540 -0.115 4.030 0.115 ;
        RECT  3.420 -0.115 3.540 0.125 ;
        RECT  2.520 -0.115 3.420 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.810 1.145 5.880 1.375 ;
        RECT  5.730 0.680 5.810 1.375 ;
        RECT  5.355 1.145 5.730 1.375 ;
        RECT  5.285 0.895 5.355 1.375 ;
        RECT  4.980 1.145 5.285 1.375 ;
        RECT  4.850 1.130 4.980 1.375 ;
        RECT  4.150 1.145 4.850 1.375 ;
        RECT  4.030 0.890 4.150 1.375 ;
        RECT  3.545 1.145 4.030 1.375 ;
        RECT  3.425 1.000 3.545 1.375 ;
        RECT  2.395 1.145 3.425 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.245 0.395 5.315 0.810 ;
        RECT  5.185 0.395 5.245 0.465 ;
        RECT  5.175 0.740 5.245 0.810 ;
        RECT  5.095 0.195 5.185 0.465 ;
        RECT  5.105 0.740 5.175 0.900 ;
        RECT  5.025 0.545 5.155 0.615 ;
        RECT  4.865 0.395 5.095 0.465 ;
        RECT  4.955 0.545 5.025 0.920 ;
        RECT  4.550 0.850 4.955 0.920 ;
        RECT  4.775 0.395 4.865 0.600 ;
        RECT  4.400 0.995 4.730 1.065 ;
        RECT  4.480 0.350 4.550 0.920 ;
        RECT  4.330 0.200 4.400 1.065 ;
        RECT  3.265 0.200 4.330 0.270 ;
        RECT  4.315 0.740 4.330 1.065 ;
        RECT  3.935 0.740 4.315 0.810 ;
        RECT  3.800 0.540 4.235 0.660 ;
        RECT  3.860 0.740 3.935 0.930 ;
        RECT  3.730 0.340 3.760 0.420 ;
        RECT  3.660 0.340 3.730 0.930 ;
        RECT  3.640 0.340 3.660 0.600 ;
        RECT  3.385 0.485 3.640 0.600 ;
        RECT  3.500 0.670 3.590 0.930 ;
        RECT  3.160 0.860 3.500 0.930 ;
        RECT  3.315 0.350 3.340 0.430 ;
        RECT  3.230 0.350 3.315 0.780 ;
        RECT  3.145 0.190 3.265 0.270 ;
        RECT  3.020 1.000 3.215 1.070 ;
        RECT  3.110 0.690 3.160 0.930 ;
        RECT  3.110 0.350 3.150 0.420 ;
        RECT  3.090 0.350 3.110 0.930 ;
        RECT  3.030 0.350 3.090 0.760 ;
        RECT  2.980 0.690 3.030 0.760 ;
        RECT  2.950 0.845 3.020 1.070 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.950 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.695 0.985 2.855 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.695 1.055 ;
        RECT  2.275 0.200 2.345 0.345 ;
        RECT  1.925 0.200 2.275 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.755 ;
        RECT  1.675 0.685 2.045 0.755 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.650 0.505 1.675 0.755 ;
        RECT  1.600 0.505 1.650 0.765 ;
        RECT  1.085 0.195 1.610 0.265 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.095 0.685 1.220 0.765 ;
        RECT  1.015 0.195 1.085 0.275 ;
        RECT  0.455 0.205 1.015 0.275 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  5.105 0.245 5.175 0.315 ;
        RECT  2.275 0.245 2.345 0.315 ;
        LAYER M2 ;
        RECT  2.225 0.245 5.225 0.315 ;
    END
END SEDFQD2BWP40

MACRO SEDFQD4BWP40
    CLASS CORE ;
    FOREIGN SEDFQD4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN SI
        ANTENNAGATEAREA 0.009600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.495 0.290 0.765 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.024800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.835 0.630 0.950 0.915 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.240000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.125 0.195 6.220 0.470 ;
        RECT  6.125 0.710 6.220 1.010 ;
        RECT  6.055 0.355 6.125 0.470 ;
        RECT  6.055 0.710 6.125 0.830 ;
        RECT  5.845 0.355 6.055 0.830 ;
        RECT  5.815 0.355 5.845 0.470 ;
        RECT  5.820 0.710 5.845 0.830 ;
        RECT  5.745 0.710 5.820 1.010 ;
        RECT  5.745 0.195 5.815 0.470 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.025200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.495 2.425 0.765 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.018400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 0.495 1.505 0.625 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.505 0.495 2.740 0.765 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.390 -0.115 6.440 0.115 ;
        RECT  6.310 -0.115 6.390 0.470 ;
        RECT  6.030 -0.115 6.310 0.115 ;
        RECT  5.910 -0.115 6.030 0.250 ;
        RECT  5.625 -0.115 5.910 0.115 ;
        RECT  5.555 -0.115 5.625 0.315 ;
        RECT  4.565 -0.115 5.555 0.115 ;
        RECT  4.455 -0.115 4.565 0.345 ;
        RECT  4.180 -0.115 4.455 0.115 ;
        RECT  4.110 -0.115 4.180 0.290 ;
        RECT  3.500 -0.115 4.110 0.115 ;
        RECT  3.380 -0.115 3.500 0.125 ;
        RECT  2.520 -0.115 3.380 0.115 ;
        RECT  2.400 -0.115 2.520 0.125 ;
        RECT  0.945 -0.115 2.400 0.115 ;
        RECT  0.815 -0.115 0.945 0.135 ;
        RECT  0.190 -0.115 0.815 0.115 ;
        RECT  0.070 -0.115 0.190 0.260 ;
        RECT  0.000 -0.115 0.070 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.385 1.145 6.440 1.375 ;
        RECT  6.315 0.715 6.385 1.375 ;
        RECT  6.030 1.145 6.315 1.375 ;
        RECT  5.910 0.905 6.030 1.375 ;
        RECT  5.625 1.145 5.910 1.375 ;
        RECT  5.555 0.970 5.625 1.375 ;
        RECT  4.150 1.145 5.555 1.375 ;
        RECT  4.030 1.050 4.150 1.375 ;
        RECT  3.545 1.145 4.030 1.375 ;
        RECT  3.425 1.000 3.545 1.375 ;
        RECT  2.395 1.145 3.425 1.375 ;
        RECT  2.275 1.130 2.395 1.375 ;
        RECT  0.950 1.145 2.275 1.375 ;
        RECT  0.810 1.125 0.950 1.375 ;
        RECT  0.190 1.145 0.810 1.375 ;
        RECT  0.070 0.990 0.190 1.375 ;
        RECT  0.000 1.145 0.070 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.125 0.195 6.220 0.470 ;
        RECT  6.125 0.710 6.220 1.010 ;
        RECT  5.745 0.195 5.775 0.470 ;
        RECT  5.745 0.710 5.775 1.010 ;
        RECT  5.670 0.545 5.765 0.615 ;
        RECT  5.600 0.545 5.670 0.880 ;
        RECT  5.245 0.780 5.600 0.880 ;
        RECT  5.470 0.465 5.500 0.600 ;
        RECT  5.400 0.200 5.470 0.600 ;
        RECT  4.730 0.200 5.400 0.270 ;
        RECT  5.100 0.995 5.385 1.065 ;
        RECT  5.170 0.340 5.245 0.880 ;
        RECT  4.895 0.340 5.170 0.410 ;
        RECT  5.030 0.480 5.100 1.065 ;
        RECT  4.970 0.480 5.030 0.610 ;
        RECT  4.345 0.995 5.030 1.065 ;
        RECT  4.885 0.805 4.960 0.925 ;
        RECT  4.825 0.340 4.895 0.640 ;
        RECT  4.545 0.855 4.885 0.925 ;
        RECT  4.785 0.520 4.825 0.640 ;
        RECT  4.715 0.715 4.775 0.785 ;
        RECT  4.715 0.200 4.730 0.465 ;
        RECT  4.645 0.200 4.715 0.785 ;
        RECT  4.470 0.715 4.545 0.925 ;
        RECT  4.220 0.715 4.470 0.785 ;
        RECT  4.270 0.900 4.345 1.065 ;
        RECT  3.900 0.900 4.270 0.970 ;
        RECT  3.825 0.200 3.900 0.970 ;
        RECT  3.265 0.200 3.825 0.270 ;
        RECT  3.680 0.340 3.750 0.790 ;
        RECT  3.615 0.340 3.680 0.595 ;
        RECT  3.380 0.485 3.615 0.595 ;
        RECT  3.500 0.670 3.590 0.930 ;
        RECT  3.155 0.860 3.500 0.930 ;
        RECT  3.300 0.355 3.340 0.425 ;
        RECT  3.300 0.680 3.330 0.785 ;
        RECT  3.230 0.355 3.300 0.785 ;
        RECT  3.145 0.190 3.265 0.270 ;
        RECT  3.005 1.000 3.215 1.070 ;
        RECT  3.110 0.690 3.155 0.930 ;
        RECT  3.110 0.350 3.150 0.420 ;
        RECT  3.085 0.350 3.110 0.930 ;
        RECT  3.030 0.350 3.085 0.760 ;
        RECT  2.965 0.690 3.030 0.760 ;
        RECT  2.935 0.845 3.005 1.070 ;
        RECT  2.890 0.355 2.960 0.505 ;
        RECT  2.890 0.845 2.935 0.915 ;
        RECT  2.820 0.355 2.890 0.915 ;
        RECT  2.695 0.985 2.855 1.075 ;
        RECT  2.425 0.355 2.820 0.425 ;
        RECT  2.420 0.845 2.820 0.915 ;
        RECT  0.455 0.985 2.695 1.055 ;
        RECT  2.275 0.200 2.345 0.345 ;
        RECT  1.925 0.200 2.275 0.270 ;
        RECT  2.120 0.845 2.195 0.915 ;
        RECT  2.120 0.355 2.175 0.425 ;
        RECT  2.050 0.355 2.120 0.915 ;
        RECT  2.045 0.355 2.050 0.755 ;
        RECT  1.675 0.685 2.045 0.755 ;
        RECT  1.845 0.345 1.975 0.435 ;
        RECT  1.845 0.825 1.960 0.915 ;
        RECT  1.055 0.345 1.845 0.415 ;
        RECT  1.030 0.840 1.845 0.915 ;
        RECT  1.650 0.505 1.675 0.755 ;
        RECT  1.600 0.505 1.650 0.765 ;
        RECT  1.085 0.195 1.610 0.265 ;
        RECT  1.220 0.695 1.600 0.765 ;
        RECT  1.095 0.685 1.220 0.765 ;
        RECT  1.015 0.195 1.085 0.275 ;
        RECT  0.455 0.205 1.015 0.275 ;
        RECT  0.735 0.480 1.015 0.550 ;
        RECT  0.730 0.480 0.735 0.915 ;
        RECT  0.645 0.360 0.730 0.915 ;
        RECT  0.630 0.360 0.645 0.695 ;
        RECT  0.560 0.575 0.630 0.695 ;
        RECT  0.380 0.205 0.455 1.055 ;
        LAYER VIA1 ;
        RECT  4.655 0.245 4.725 0.315 ;
        RECT  2.275 0.245 2.345 0.315 ;
        LAYER M2 ;
        RECT  2.225 0.245 4.775 0.315 ;
    END
END SEDFQD4BWP40

MACRO TAPCELLBWP40
    CLASS CORE ;
    FOREIGN TAPCELLBWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 -0.115 0.560 0.115 ;
        RECT  0.220 -0.115 0.340 0.410 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.145 0.560 1.375 ;
        RECT  0.220 0.780 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
END TAPCELLBWP40

MACRO TIEHBWP40
    CLASS CORE ;
    FOREIGN TIEHBWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.051750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.735 0.385 1.045 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.175 -0.115 0.420 0.115 ;
        RECT  0.085 -0.115 0.175 0.465 ;
        RECT  0.000 -0.115 0.085 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.175 1.145 0.420 1.375 ;
        RECT  0.085 0.745 0.175 1.375 ;
        RECT  0.000 1.145 0.085 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 0.185 0.365 0.615 ;
        RECT  0.190 0.545 0.295 0.615 ;
    END
END TIEHBWP40

MACRO TIELBWP40
    CLASS CORE ;
    FOREIGN TIELBWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.420 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.040250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 0.185 0.385 0.485 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.175 -0.115 0.420 0.115 ;
        RECT  0.085 -0.115 0.175 0.465 ;
        RECT  0.000 -0.115 0.085 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.175 1.145 0.420 1.375 ;
        RECT  0.085 0.745 0.175 1.375 ;
        RECT  0.000 1.145 0.085 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.295 0.555 0.365 1.045 ;
        RECT  0.190 0.555 0.295 0.625 ;
    END
END TIELBWP40

MACRO XNR2D0BWP40
    CLASS CORE ;
    FOREIGN XNR2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.195 1.365 1.065 ;
        RECT  1.280 0.195 1.295 0.470 ;
        RECT  1.255 0.980 1.295 1.065 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 0.350 1.085 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.155 -0.115 1.400 0.115 ;
        RECT  1.055 -0.115 1.155 0.230 ;
        RECT  0.260 -0.115 1.055 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.145 1.400 1.375 ;
        RECT  1.045 0.995 1.145 1.375 ;
        RECT  0.340 1.145 1.045 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.160 0.515 1.225 0.830 ;
        RECT  1.155 0.515 1.160 0.925 ;
        RECT  1.090 0.760 1.155 0.925 ;
        RECT  0.710 0.855 1.090 0.925 ;
        RECT  0.850 0.705 0.970 0.775 ;
        RECT  0.850 0.200 0.945 0.270 ;
        RECT  0.725 0.995 0.905 1.075 ;
        RECT  0.780 0.200 0.850 0.775 ;
        RECT  0.330 0.200 0.780 0.270 ;
        RECT  0.510 0.995 0.725 1.065 ;
        RECT  0.620 0.350 0.710 0.925 ;
        RECT  0.425 0.350 0.525 0.790 ;
        RECT  0.440 0.860 0.510 1.065 ;
        RECT  0.125 0.860 0.440 0.930 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR2D0BWP40

MACRO XNR2D1BWP40
    CLASS CORE ;
    FOREIGN XNR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.092000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.195 1.365 1.075 ;
        RECT  1.280 0.195 1.295 0.470 ;
        RECT  1.255 0.990 1.295 1.075 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 0.350 1.085 0.630 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.145 -0.115 1.400 0.115 ;
        RECT  1.045 -0.115 1.145 0.230 ;
        RECT  0.260 -0.115 1.045 0.115 ;
        RECT  0.260 0.355 0.350 0.425 ;
        RECT  0.190 -0.115 0.260 0.425 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.145 1.400 1.375 ;
        RECT  1.045 0.995 1.145 1.375 ;
        RECT  0.340 1.145 1.045 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.155 0.515 1.225 0.925 ;
        RECT  0.710 0.855 1.155 0.925 ;
        RECT  0.850 0.705 0.970 0.775 ;
        RECT  0.850 0.200 0.945 0.270 ;
        RECT  0.725 0.995 0.905 1.075 ;
        RECT  0.780 0.200 0.850 0.775 ;
        RECT  0.330 0.200 0.780 0.270 ;
        RECT  0.510 0.995 0.725 1.065 ;
        RECT  0.620 0.350 0.710 0.925 ;
        RECT  0.425 0.350 0.525 0.790 ;
        RECT  0.440 0.860 0.510 1.065 ;
        RECT  0.125 0.860 0.440 0.930 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.275 0.120 0.435 ;
        RECT  0.035 0.275 0.105 1.040 ;
    END
END XNR2D1BWP40

MACRO XNR2D2BWP40
    CLASS CORE ;
    FOREIGN XNR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 0.355 1.925 0.770 ;
        RECT  1.695 0.355 1.845 0.480 ;
        RECT  1.695 0.700 1.845 0.770 ;
        RECT  1.625 0.195 1.695 0.480 ;
        RECT  1.625 0.700 1.695 1.055 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.155 0.495 1.405 0.625 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 -0.115 1.960 0.115 ;
        RECT  1.800 -0.115 1.900 0.275 ;
        RECT  1.530 -0.115 1.800 0.115 ;
        RECT  1.410 -0.115 1.530 0.130 ;
        RECT  0.335 -0.115 1.410 0.115 ;
        RECT  0.225 -0.115 0.335 0.235 ;
        RECT  0.000 -0.115 0.225 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.895 1.145 1.960 1.375 ;
        RECT  1.810 0.850 1.895 1.375 ;
        RECT  1.530 1.145 1.810 1.375 ;
        RECT  1.440 0.840 1.530 1.375 ;
        RECT  0.340 1.145 1.440 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.545 0.550 1.745 0.620 ;
        RECT  1.475 0.200 1.545 0.620 ;
        RECT  0.685 0.200 1.475 0.270 ;
        RECT  1.085 0.785 1.360 0.855 ;
        RECT  1.085 0.350 1.305 0.420 ;
        RECT  1.015 0.350 1.085 0.855 ;
        RECT  0.825 0.340 0.905 0.980 ;
        RECT  0.385 0.910 0.825 0.980 ;
        RECT  0.685 0.770 0.735 0.840 ;
        RECT  0.615 0.200 0.685 0.840 ;
        RECT  0.455 0.290 0.525 0.830 ;
        RECT  0.315 0.305 0.385 0.980 ;
        RECT  0.140 0.305 0.315 0.375 ;
        RECT  0.035 0.910 0.315 0.980 ;
        RECT  0.050 0.185 0.140 0.375 ;
    END
END XNR2D2BWP40

MACRO XNR2D3BWP40
    CLASS CORE ;
    FOREIGN XNR2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.222300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.260 0.200 2.345 0.480 ;
        RECT  2.260 0.775 2.345 1.055 ;
        RECT  2.240 0.200 2.260 1.055 ;
        RECT  2.100 0.355 2.240 0.885 ;
        RECT  1.905 0.355 2.100 0.470 ;
        RECT  1.925 0.775 2.100 0.885 ;
        RECT  1.835 0.775 1.925 1.055 ;
        RECT  1.810 0.195 1.905 0.470 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.465 0.280 0.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.525 0.495 1.590 0.620 ;
        RECT  1.435 0.495 1.525 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.020 -0.115 2.120 0.275 ;
        RECT  1.730 -0.115 2.020 0.115 ;
        RECT  1.610 -0.115 1.730 0.130 ;
        RECT  0.545 -0.115 1.610 0.115 ;
        RECT  0.435 -0.115 0.545 0.235 ;
        RECT  0.160 -0.115 0.435 0.115 ;
        RECT  0.060 -0.115 0.160 0.370 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.020 0.985 2.120 1.375 ;
        RECT  1.705 1.145 2.020 1.375 ;
        RECT  1.635 0.695 1.705 1.375 ;
        RECT  0.560 1.145 1.635 1.375 ;
        RECT  0.440 1.120 0.560 1.375 ;
        RECT  0.160 1.145 0.440 1.375 ;
        RECT  0.060 0.890 0.160 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 0.540 1.965 0.615 ;
        RECT  1.670 0.200 1.740 0.615 ;
        RECT  0.890 0.200 1.670 0.270 ;
        RECT  1.365 0.340 1.540 0.410 ;
        RECT  1.365 0.840 1.530 0.910 ;
        RECT  1.275 0.340 1.365 0.910 ;
        RECT  1.100 0.345 1.180 1.050 ;
        RECT  1.050 0.345 1.100 0.485 ;
        RECT  0.665 0.290 0.680 0.460 ;
        RECT  0.665 0.700 0.680 0.870 ;
        RECT  0.575 0.520 0.610 0.650 ;
        RECT  0.505 0.305 0.575 1.050 ;
        RECT  0.360 0.305 0.505 0.375 ;
        RECT  0.265 0.890 0.505 1.050 ;
        RECT  0.270 0.185 0.360 0.375 ;
        RECT  0.575 0.980 1.100 1.050 ;
        RECT  0.890 0.790 0.980 0.860 ;
        RECT  0.820 0.200 0.890 0.860 ;
        RECT  0.680 0.290 0.750 0.870 ;
    END
END XNR2D3BWP40

MACRO XNR2D4BWP40
    CLASS CORE ;
    FOREIGN XNR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.195 2.695 1.055 ;
        RECT  2.615 0.195 2.625 0.905 ;
        RECT  2.485 0.355 2.615 0.905 ;
        RECT  2.315 0.355 2.485 0.480 ;
        RECT  2.315 0.775 2.485 0.905 ;
        RECT  2.245 0.195 2.315 0.480 ;
        RECT  2.245 0.775 2.315 1.055 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 0.495 0.385 0.765 ;
        RECT  0.035 0.495 0.305 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.785 0.495 2.020 0.625 ;
        RECT  1.715 0.495 1.785 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 -0.115 2.940 0.115 ;
        RECT  2.800 -0.115 2.900 0.460 ;
        RECT  2.520 -0.115 2.800 0.115 ;
        RECT  2.420 -0.115 2.520 0.275 ;
        RECT  2.140 -0.115 2.420 0.115 ;
        RECT  2.020 -0.115 2.140 0.130 ;
        RECT  0.905 -0.115 2.020 0.115 ;
        RECT  0.795 -0.115 0.905 0.280 ;
        RECT  0.525 -0.115 0.795 0.115 ;
        RECT  0.415 -0.115 0.525 0.235 ;
        RECT  0.135 -0.115 0.415 0.115 ;
        RECT  0.050 -0.115 0.135 0.405 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.720 2.900 1.375 ;
        RECT  2.520 1.145 2.800 1.375 ;
        RECT  2.420 0.985 2.520 1.375 ;
        RECT  2.120 1.145 2.420 1.375 ;
        RECT  2.040 0.760 2.120 1.375 ;
        RECT  0.910 1.145 2.040 1.375 ;
        RECT  0.790 1.120 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 1.120 0.530 1.375 ;
        RECT  0.135 1.145 0.410 1.375 ;
        RECT  0.050 0.735 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.315 0.355 2.415 0.480 ;
        RECT  2.315 0.775 2.415 0.905 ;
        RECT  2.245 0.195 2.315 0.480 ;
        RECT  2.245 0.775 2.315 1.055 ;
        RECT  2.165 0.550 2.305 0.620 ;
        RECT  2.095 0.200 2.165 0.620 ;
        RECT  1.215 0.200 2.095 0.270 ;
        RECT  1.640 0.340 1.960 0.410 ;
        RECT  1.640 0.945 1.960 1.015 ;
        RECT  1.570 0.340 1.640 1.015 ;
        RECT  1.405 0.345 1.490 1.050 ;
        RECT  0.545 0.980 1.405 1.050 ;
        RECT  1.215 0.790 1.300 0.860 ;
        RECT  1.145 0.200 1.215 0.860 ;
        RECT  0.985 0.195 1.075 0.450 ;
        RECT  0.965 0.720 1.070 0.910 ;
        RECT  0.835 0.380 0.985 0.450 ;
        RECT  0.835 0.720 0.965 0.795 ;
        RECT  0.750 0.380 0.835 0.795 ;
        RECT  0.715 0.380 0.750 0.450 ;
        RECT  0.715 0.720 0.750 0.795 ;
        RECT  0.615 0.245 0.715 0.450 ;
        RECT  0.615 0.720 0.715 0.900 ;
        RECT  0.545 0.520 0.680 0.650 ;
        RECT  0.475 0.305 0.545 1.050 ;
        RECT  0.330 0.305 0.475 0.375 ;
        RECT  0.240 0.185 0.330 0.375 ;
        RECT  0.240 0.890 0.475 1.050 ;
    END
END XNR2D4BWP40

MACRO XNR2D6BWP40
    CLASS CORE ;
    FOREIGN XNR2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.357000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.175 0.195 3.265 0.485 ;
        RECT  3.180 0.775 3.260 1.060 ;
        RECT  2.975 0.775 3.180 0.905 ;
        RECT  2.975 0.355 3.175 0.485 ;
        RECT  2.885 0.355 2.975 0.905 ;
        RECT  2.880 0.195 2.885 0.905 ;
        RECT  2.795 0.195 2.880 1.055 ;
        RECT  2.765 0.355 2.795 0.905 ;
        RECT  2.500 0.355 2.765 0.480 ;
        RECT  2.500 0.775 2.765 0.905 ;
        RECT  2.425 0.195 2.500 0.480 ;
        RECT  2.420 0.775 2.500 1.055 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.093600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.390 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.495 2.205 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.115 3.500 0.115 ;
        RECT  3.360 -0.115 3.460 0.480 ;
        RECT  3.090 -0.115 3.360 0.115 ;
        RECT  2.970 -0.115 3.090 0.255 ;
        RECT  2.700 -0.115 2.970 0.115 ;
        RECT  2.600 -0.115 2.700 0.275 ;
        RECT  2.320 -0.115 2.600 0.115 ;
        RECT  2.200 -0.115 2.320 0.130 ;
        RECT  1.100 -0.115 2.200 0.115 ;
        RECT  0.980 -0.115 1.100 0.230 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.210 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.210 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 1.145 3.500 1.375 ;
        RECT  3.360 0.720 3.460 1.375 ;
        RECT  3.085 1.145 3.360 1.375 ;
        RECT  2.975 0.985 3.085 1.375 ;
        RECT  2.700 1.145 2.975 1.375 ;
        RECT  2.600 0.985 2.700 1.375 ;
        RECT  2.320 1.145 2.600 1.375 ;
        RECT  2.200 0.880 2.320 1.375 ;
        RECT  1.100 1.145 2.200 1.375 ;
        RECT  0.980 1.120 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 1.120 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.175 0.195 3.265 0.485 ;
        RECT  3.180 0.775 3.260 1.060 ;
        RECT  3.045 0.775 3.180 0.905 ;
        RECT  3.045 0.355 3.175 0.485 ;
        RECT  2.500 0.355 2.695 0.480 ;
        RECT  2.500 0.775 2.695 0.905 ;
        RECT  2.425 0.195 2.500 0.480 ;
        RECT  2.420 0.775 2.500 1.055 ;
        RECT  2.345 0.550 2.650 0.620 ;
        RECT  2.275 0.200 2.345 0.620 ;
        RECT  1.455 0.200 2.275 0.270 ;
        RECT  1.980 0.340 2.140 0.410 ;
        RECT  1.980 0.960 2.090 1.030 ;
        RECT  1.910 0.340 1.980 1.030 ;
        RECT  1.700 0.360 1.770 1.040 ;
        RECT  1.615 0.360 1.700 0.440 ;
        RECT  0.660 0.970 1.700 1.040 ;
        RECT  1.455 0.790 1.570 0.860 ;
        RECT  1.385 0.200 1.455 0.860 ;
        RECT  1.210 0.330 1.290 0.900 ;
        RECT  0.785 0.330 1.210 0.410 ;
        RECT  0.035 0.845 0.590 0.915 ;
        RECT  0.785 0.820 1.210 0.900 ;
        RECT  0.660 0.520 0.890 0.650 ;
        RECT  0.590 0.280 0.660 1.040 ;
        RECT  0.035 0.280 0.590 0.375 ;
    END
END XNR2D6BWP40

MACRO XNR2D8BWP40
    CLASS CORE ;
    FOREIGN XNR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.468000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.205 4.375 0.485 ;
        RECT  4.305 0.780 4.375 1.065 ;
        RECT  3.995 0.355 4.305 0.485 ;
        RECT  4.005 0.780 4.305 0.905 ;
        RECT  3.925 0.780 4.005 1.065 ;
        RECT  3.925 0.205 3.995 0.485 ;
        RECT  3.815 0.355 3.925 0.485 ;
        RECT  3.815 0.780 3.925 0.905 ;
        RECT  3.610 0.355 3.815 0.905 ;
        RECT  3.605 0.205 3.610 1.065 ;
        RECT  3.540 0.205 3.605 0.480 ;
        RECT  3.535 0.780 3.605 1.065 ;
        RECT  3.230 0.355 3.540 0.480 ;
        RECT  3.230 0.780 3.535 0.905 ;
        RECT  3.160 0.195 3.230 0.480 ;
        RECT  3.160 0.780 3.230 1.065 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.128000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.385 0.495 0.665 0.625 ;
        RECT  0.315 0.495 0.385 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.495 2.915 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 -0.115 4.620 0.115 ;
        RECT  4.480 -0.115 4.580 0.485 ;
        RECT  4.200 -0.115 4.480 0.115 ;
        RECT  4.100 -0.115 4.200 0.275 ;
        RECT  3.820 -0.115 4.100 0.115 ;
        RECT  3.720 -0.115 3.820 0.275 ;
        RECT  3.435 -0.115 3.720 0.115 ;
        RECT  3.335 -0.115 3.435 0.275 ;
        RECT  3.035 -0.115 3.335 0.115 ;
        RECT  2.960 -0.115 3.035 0.415 ;
        RECT  1.650 -0.115 2.960 0.115 ;
        RECT  1.580 -0.115 1.650 0.275 ;
        RECT  1.295 -0.115 1.580 0.115 ;
        RECT  1.170 -0.115 1.295 0.245 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.215 ;
        RECT  0.535 -0.115 0.790 0.115 ;
        RECT  0.405 -0.115 0.535 0.240 ;
        RECT  0.135 -0.115 0.405 0.115 ;
        RECT  0.050 -0.115 0.135 0.495 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 1.145 4.620 1.375 ;
        RECT  4.480 0.705 4.580 1.375 ;
        RECT  4.200 1.145 4.480 1.375 ;
        RECT  4.100 0.985 4.200 1.375 ;
        RECT  3.820 1.145 4.100 1.375 ;
        RECT  3.720 0.985 3.820 1.375 ;
        RECT  3.435 1.145 3.720 1.375 ;
        RECT  3.335 0.985 3.435 1.375 ;
        RECT  3.055 1.145 3.335 1.375 ;
        RECT  2.935 1.130 3.055 1.375 ;
        RECT  1.670 1.145 2.935 1.375 ;
        RECT  1.560 0.980 1.670 1.375 ;
        RECT  1.285 1.145 1.560 1.375 ;
        RECT  1.175 0.980 1.285 1.375 ;
        RECT  0.905 1.145 1.175 1.375 ;
        RECT  0.795 1.025 0.905 1.375 ;
        RECT  0.535 1.145 0.795 1.375 ;
        RECT  0.405 1.045 0.535 1.375 ;
        RECT  0.135 1.145 0.405 1.375 ;
        RECT  0.050 0.720 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.205 4.375 0.485 ;
        RECT  4.305 0.780 4.375 1.065 ;
        RECT  3.995 0.355 4.305 0.485 ;
        RECT  4.005 0.780 4.305 0.905 ;
        RECT  3.925 0.780 4.005 1.065 ;
        RECT  3.925 0.205 3.995 0.485 ;
        RECT  3.885 0.355 3.925 0.485 ;
        RECT  3.885 0.780 3.925 0.905 ;
        RECT  3.230 0.355 3.535 0.480 ;
        RECT  3.230 0.780 3.535 0.905 ;
        RECT  3.160 0.195 3.230 0.480 ;
        RECT  3.160 0.780 3.230 1.065 ;
        RECT  3.080 0.550 3.495 0.625 ;
        RECT  3.010 0.550 3.080 1.060 ;
        RECT  2.555 0.990 3.010 1.060 ;
        RECT  2.705 0.850 2.875 0.920 ;
        RECT  2.705 0.350 2.860 0.420 ;
        RECT  2.635 0.350 2.705 0.920 ;
        RECT  2.555 0.195 2.685 0.265 ;
        RECT  2.485 0.195 2.555 1.060 ;
        RECT  1.735 0.195 2.485 0.265 ;
        RECT  1.740 0.990 2.485 1.060 ;
        RECT  2.325 0.340 2.405 0.920 ;
        RECT  1.350 0.545 2.325 0.615 ;
        RECT  1.230 0.360 2.045 0.430 ;
        RECT  1.230 0.810 2.045 0.880 ;
        RECT  1.145 0.360 1.230 0.880 ;
        RECT  0.975 0.360 1.145 0.430 ;
        RECT  0.975 0.810 1.145 0.880 ;
        RECT  0.855 0.530 1.065 0.620 ;
        RECT  0.775 0.310 0.855 0.955 ;
        RECT  0.320 0.310 0.775 0.380 ;
        RECT  0.220 0.885 0.775 0.955 ;
        RECT  0.250 0.220 0.320 0.380 ;
    END
END XNR2D8BWP40

MACRO XNR3D0BWP40
    CLASS CORE ;
    FOREIGN XNR3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.625 1.045 ;
        RECT  2.535 0.185 2.555 0.315 ;
        RECT  2.540 0.895 2.555 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.295 0.215 2.345 0.485 ;
        RECT  2.215 0.215 2.295 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.033000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.115 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 -0.115 2.660 0.115 ;
        RECT  2.290 -0.115 2.410 0.140 ;
        RECT  1.505 -0.115 2.290 0.115 ;
        RECT  1.435 -0.115 1.505 0.465 ;
        RECT  1.140 -0.115 1.435 0.115 ;
        RECT  1.060 -0.115 1.140 0.280 ;
        RECT  0.320 -0.115 1.060 0.115 ;
        RECT  0.240 -0.115 0.320 0.355 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.145 2.660 1.375 ;
        RECT  2.290 1.120 2.410 1.375 ;
        RECT  1.580 1.145 2.290 1.375 ;
        RECT  1.510 0.835 1.580 1.375 ;
        RECT  1.410 0.835 1.510 0.905 ;
        RECT  1.190 1.145 1.510 1.375 ;
        RECT  1.070 1.135 1.190 1.375 ;
        RECT  0.340 1.145 1.070 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.470 0.535 2.485 0.655 ;
        RECT  2.395 0.535 2.470 1.050 ;
        RECT  1.940 0.980 2.395 1.050 ;
        RECT  2.110 0.840 2.180 0.910 ;
        RECT  2.040 0.205 2.110 0.910 ;
        RECT  1.645 0.205 2.040 0.275 ;
        RECT  1.870 0.350 1.940 1.050 ;
        RECT  1.825 0.350 1.870 0.450 ;
        RECT  1.715 0.520 1.785 0.765 ;
        RECT  1.320 0.695 1.715 0.765 ;
        RECT  1.575 0.205 1.645 0.615 ;
        RECT  1.480 0.545 1.575 0.615 ;
        RECT  0.795 0.995 1.440 1.065 ;
        RECT  1.240 0.330 1.320 0.900 ;
        RECT  0.875 0.195 0.945 0.915 ;
        RECT  0.505 0.195 0.875 0.265 ;
        RECT  0.725 0.340 0.795 1.065 ;
        RECT  0.610 0.340 0.725 0.410 ;
        RECT  0.655 0.920 0.725 1.065 ;
        RECT  0.575 0.490 0.655 0.800 ;
        RECT  0.465 0.730 0.575 0.800 ;
        RECT  0.435 0.195 0.505 0.620 ;
        RECT  0.385 0.730 0.465 0.930 ;
        RECT  0.335 0.540 0.435 0.620 ;
        RECT  0.130 0.860 0.385 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D0BWP40

MACRO XNR3D1BWP40
    CLASS CORE ;
    FOREIGN XNR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.086825 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.185 2.625 1.045 ;
        RECT  2.535 0.185 2.555 0.465 ;
        RECT  2.540 0.730 2.555 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.030200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.295 0.215 2.345 0.485 ;
        RECT  2.215 0.215 2.295 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.033000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.115 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 -0.115 2.660 0.115 ;
        RECT  2.290 -0.115 2.410 0.140 ;
        RECT  1.505 -0.115 2.290 0.115 ;
        RECT  1.435 -0.115 1.505 0.465 ;
        RECT  1.140 -0.115 1.435 0.115 ;
        RECT  1.060 -0.115 1.140 0.405 ;
        RECT  0.320 -0.115 1.060 0.115 ;
        RECT  0.240 -0.115 0.320 0.355 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.145 2.660 1.375 ;
        RECT  2.290 1.120 2.410 1.375 ;
        RECT  1.580 1.145 2.290 1.375 ;
        RECT  1.510 0.835 1.580 1.375 ;
        RECT  1.410 0.835 1.510 0.905 ;
        RECT  1.190 1.145 1.510 1.375 ;
        RECT  1.070 1.135 1.190 1.375 ;
        RECT  0.340 1.145 1.070 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.470 0.535 2.485 0.655 ;
        RECT  2.395 0.535 2.470 1.050 ;
        RECT  1.940 0.980 2.395 1.050 ;
        RECT  2.110 0.840 2.180 0.910 ;
        RECT  2.040 0.205 2.110 0.910 ;
        RECT  1.645 0.205 2.040 0.275 ;
        RECT  1.870 0.350 1.940 1.050 ;
        RECT  1.825 0.350 1.870 0.450 ;
        RECT  1.715 0.520 1.785 0.765 ;
        RECT  1.320 0.695 1.715 0.765 ;
        RECT  1.575 0.205 1.645 0.615 ;
        RECT  1.480 0.545 1.575 0.615 ;
        RECT  0.795 0.995 1.440 1.065 ;
        RECT  1.240 0.330 1.320 0.900 ;
        RECT  0.875 0.195 0.945 0.915 ;
        RECT  0.505 0.195 0.875 0.265 ;
        RECT  0.725 0.340 0.795 1.065 ;
        RECT  0.610 0.340 0.725 0.410 ;
        RECT  0.655 0.915 0.725 1.065 ;
        RECT  0.575 0.490 0.655 0.800 ;
        RECT  0.465 0.730 0.575 0.800 ;
        RECT  0.435 0.195 0.505 0.620 ;
        RECT  0.385 0.730 0.465 0.930 ;
        RECT  0.335 0.540 0.435 0.620 ;
        RECT  0.130 0.860 0.385 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D1BWP40

MACRO XNR3D2BWP40
    CLASS CORE ;
    FOREIGN XNR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.113250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.680 0.355 2.765 0.795 ;
        RECT  2.590 0.355 2.680 0.465 ;
        RECT  2.590 0.715 2.680 0.795 ;
        RECT  2.490 0.185 2.590 0.465 ;
        RECT  2.490 0.715 2.590 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.030200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.215 2.345 0.485 ;
        RECT  2.190 0.215 2.270 0.655 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.033000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.115 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.280 ;
        RECT  2.385 -0.115 2.670 0.115 ;
        RECT  2.265 -0.115 2.385 0.140 ;
        RECT  1.505 -0.115 2.265 0.115 ;
        RECT  1.435 -0.115 1.505 0.465 ;
        RECT  1.140 -0.115 1.435 0.115 ;
        RECT  1.060 -0.115 1.140 0.405 ;
        RECT  0.320 -0.115 1.060 0.115 ;
        RECT  0.240 -0.115 0.320 0.355 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.905 2.750 1.375 ;
        RECT  2.385 1.145 2.670 1.375 ;
        RECT  2.265 1.120 2.385 1.375 ;
        RECT  1.580 1.145 2.265 1.375 ;
        RECT  1.510 0.835 1.580 1.375 ;
        RECT  1.410 0.835 1.510 0.905 ;
        RECT  1.190 1.145 1.510 1.375 ;
        RECT  1.070 1.135 1.190 1.375 ;
        RECT  0.340 1.145 1.070 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.420 0.555 2.540 0.635 ;
        RECT  2.345 0.555 2.420 1.050 ;
        RECT  1.940 0.980 2.345 1.050 ;
        RECT  2.110 0.840 2.180 0.910 ;
        RECT  2.040 0.205 2.110 0.910 ;
        RECT  1.645 0.205 2.040 0.275 ;
        RECT  1.870 0.350 1.940 1.050 ;
        RECT  1.825 0.350 1.870 0.450 ;
        RECT  1.715 0.520 1.785 0.765 ;
        RECT  1.320 0.695 1.715 0.765 ;
        RECT  1.575 0.205 1.645 0.615 ;
        RECT  1.480 0.545 1.575 0.615 ;
        RECT  0.795 0.995 1.440 1.065 ;
        RECT  1.240 0.330 1.320 0.900 ;
        RECT  0.875 0.195 0.945 0.915 ;
        RECT  0.505 0.195 0.875 0.265 ;
        RECT  0.725 0.340 0.795 1.065 ;
        RECT  0.610 0.340 0.725 0.410 ;
        RECT  0.660 0.915 0.725 1.065 ;
        RECT  0.575 0.490 0.655 0.800 ;
        RECT  0.465 0.730 0.575 0.800 ;
        RECT  0.435 0.195 0.505 0.620 ;
        RECT  0.385 0.730 0.465 0.930 ;
        RECT  0.335 0.540 0.435 0.620 ;
        RECT  0.130 0.860 0.385 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D2BWP40

MACRO XNR3D4BWP40
    CLASS CORE ;
    FOREIGN XNR3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.226500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.185 3.430 0.465 ;
        RECT  3.395 0.715 3.430 1.045 ;
        RECT  3.330 0.185 3.395 1.045 ;
        RECT  3.185 0.350 3.330 0.840 ;
        RECT  3.025 0.350 3.185 0.465 ;
        RECT  3.025 0.715 3.185 0.840 ;
        RECT  2.935 0.185 3.025 0.465 ;
        RECT  2.935 0.715 3.025 1.045 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.060400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.390 0.215 2.495 0.650 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.033000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.495 1.095 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.640 0.115 ;
        RECT  3.510 -0.115 3.590 0.475 ;
        RECT  3.230 -0.115 3.510 0.115 ;
        RECT  3.110 -0.115 3.230 0.250 ;
        RECT  2.845 -0.115 3.110 0.115 ;
        RECT  2.735 -0.115 2.845 0.385 ;
        RECT  2.475 -0.115 2.735 0.115 ;
        RECT  2.355 -0.115 2.475 0.140 ;
        RECT  1.670 -0.115 2.355 0.115 ;
        RECT  1.595 -0.115 1.670 0.435 ;
        RECT  1.120 -0.115 1.595 0.115 ;
        RECT  1.040 -0.115 1.120 0.405 ;
        RECT  0.320 -0.115 1.040 0.115 ;
        RECT  0.240 -0.115 0.320 0.355 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 1.145 3.640 1.375 ;
        RECT  3.510 0.695 3.590 1.375 ;
        RECT  3.230 1.145 3.510 1.375 ;
        RECT  3.110 0.955 3.230 1.375 ;
        RECT  2.845 1.145 3.110 1.375 ;
        RECT  2.725 1.110 2.845 1.375 ;
        RECT  2.475 1.145 2.725 1.375 ;
        RECT  2.355 1.120 2.475 1.375 ;
        RECT  1.790 1.145 2.355 1.375 ;
        RECT  1.710 0.815 1.790 1.375 ;
        RECT  1.580 0.815 1.710 0.895 ;
        RECT  1.140 1.145 1.710 1.375 ;
        RECT  1.020 1.115 1.140 1.375 ;
        RECT  0.340 1.145 1.020 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.025 0.350 3.115 0.465 ;
        RECT  3.025 0.715 3.115 0.840 ;
        RECT  2.935 0.185 3.025 0.465 ;
        RECT  2.935 0.715 3.025 1.045 ;
        RECT  2.820 0.545 3.020 0.630 ;
        RECT  2.725 0.545 2.820 1.020 ;
        RECT  2.105 0.945 2.725 1.020 ;
        RECT  2.565 0.195 2.640 0.855 ;
        RECT  2.260 0.760 2.565 0.855 ;
        RECT  2.175 0.205 2.260 0.855 ;
        RECT  1.815 0.205 2.175 0.275 ;
        RECT  2.035 0.350 2.105 1.020 ;
        RECT  1.935 0.350 2.035 0.435 ;
        RECT  1.960 0.945 2.035 1.020 ;
        RECT  1.895 0.520 1.965 0.745 ;
        RECT  1.490 0.675 1.895 0.745 ;
        RECT  1.740 0.205 1.815 0.605 ;
        RECT  1.630 0.535 1.740 0.605 ;
        RECT  0.790 0.975 1.595 1.045 ;
        RECT  1.410 0.330 1.490 0.900 ;
        RECT  1.235 0.245 1.310 0.905 ;
        RECT  0.930 0.835 1.235 0.905 ;
        RECT  0.860 0.195 0.930 0.905 ;
        RECT  0.480 0.195 0.860 0.265 ;
        RECT  0.720 0.340 0.790 1.045 ;
        RECT  0.590 0.340 0.720 0.410 ;
        RECT  0.640 0.925 0.720 1.045 ;
        RECT  0.555 0.490 0.650 0.800 ;
        RECT  0.465 0.730 0.555 0.800 ;
        RECT  0.400 0.195 0.480 0.620 ;
        RECT  0.385 0.730 0.465 0.930 ;
        RECT  0.340 0.540 0.400 0.620 ;
        RECT  0.130 0.860 0.385 0.930 ;
        RECT  0.105 0.200 0.130 0.360 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.200 0.105 1.040 ;
    END
END XNR3D4BWP40

MACRO XNR4D0BWP40
    CLASS CORE ;
    FOREIGN XNR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.058300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.715 2.540 0.785 ;
        RECT  2.395 0.215 2.485 0.785 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.645 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.520 2.765 0.640 ;
        RECT  2.555 0.355 2.625 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.495 3.605 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.540 -0.115 3.780 0.115 ;
        RECT  3.470 -0.115 3.540 0.415 ;
        RECT  2.710 -0.115 3.470 0.115 ;
        RECT  2.610 -0.115 2.710 0.275 ;
        RECT  1.540 -0.115 2.610 0.115 ;
        RECT  1.470 -0.115 1.540 0.445 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 1.145 3.780 1.375 ;
        RECT  3.430 0.990 3.530 1.375 ;
        RECT  2.720 1.145 3.430 1.375 ;
        RECT  2.600 1.115 2.720 1.375 ;
        RECT  1.580 1.145 2.600 1.375 ;
        RECT  1.500 0.985 1.580 1.375 ;
        RECT  1.230 1.145 1.500 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.290 3.745 1.015 ;
        RECT  3.655 0.290 3.675 0.430 ;
        RECT  3.655 0.850 3.675 1.015 ;
        RECT  3.230 0.850 3.655 0.920 ;
        RECT  3.330 0.200 3.400 0.660 ;
        RECT  2.915 0.200 3.330 0.270 ;
        RECT  3.150 0.530 3.230 0.920 ;
        RECT  3.080 0.350 3.150 0.430 ;
        RECT  3.010 0.350 3.080 1.045 ;
        RECT  2.630 0.975 3.010 1.045 ;
        RECT  2.845 0.200 2.915 0.890 ;
        RECT  2.810 0.785 2.845 0.890 ;
        RECT  2.550 0.855 2.630 1.045 ;
        RECT  2.290 0.855 2.550 0.925 ;
        RECT  2.270 0.995 2.435 1.075 ;
        RECT  2.220 0.195 2.290 0.925 ;
        RECT  2.130 0.995 2.270 1.065 ;
        RECT  1.690 0.195 2.220 0.265 ;
        RECT  2.060 0.335 2.130 1.065 ;
        RECT  1.990 0.335 2.060 0.405 ;
        RECT  1.950 0.995 2.060 1.065 ;
        RECT  1.910 0.500 1.990 0.915 ;
        RECT  1.360 0.845 1.910 0.915 ;
        RECT  1.770 0.335 1.840 0.775 ;
        RECT  1.700 0.705 1.770 0.775 ;
        RECT  1.610 0.195 1.690 0.615 ;
        RECT  1.540 0.545 1.610 0.615 ;
        RECT  1.270 0.995 1.410 1.075 ;
        RECT  1.280 0.305 1.360 0.915 ;
        RECT  0.775 0.995 1.270 1.065 ;
        RECT  1.130 0.355 1.200 0.915 ;
        RECT  0.990 0.355 1.130 0.425 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.910 0.195 0.990 0.425 ;
        RECT  0.340 0.195 0.910 0.265 ;
        RECT  0.690 0.350 0.775 1.065 ;
        RECT  0.525 0.890 0.610 1.075 ;
        RECT  0.455 0.350 0.545 0.820 ;
        RECT  0.130 0.890 0.525 0.960 ;
        RECT  0.105 0.890 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D0BWP40

MACRO XNR4D1BWP40
    CLASS CORE ;
    FOREIGN XNR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.096700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.485 0.715 2.540 0.785 ;
        RECT  2.395 0.215 2.485 0.785 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.645 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.520 2.765 0.640 ;
        RECT  2.555 0.355 2.625 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.515 0.495 3.605 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.540 -0.115 3.780 0.115 ;
        RECT  3.470 -0.115 3.540 0.415 ;
        RECT  2.710 -0.115 3.470 0.115 ;
        RECT  2.610 -0.115 2.710 0.275 ;
        RECT  1.540 -0.115 2.610 0.115 ;
        RECT  1.470 -0.115 1.540 0.445 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.530 1.145 3.780 1.375 ;
        RECT  3.430 0.990 3.530 1.375 ;
        RECT  2.720 1.145 3.430 1.375 ;
        RECT  2.600 1.115 2.720 1.375 ;
        RECT  1.580 1.145 2.600 1.375 ;
        RECT  1.500 0.985 1.580 1.375 ;
        RECT  1.230 1.145 1.500 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.290 3.745 1.015 ;
        RECT  3.655 0.290 3.675 0.430 ;
        RECT  3.655 0.850 3.675 1.015 ;
        RECT  3.230 0.850 3.655 0.920 ;
        RECT  3.330 0.200 3.400 0.660 ;
        RECT  2.915 0.200 3.330 0.270 ;
        RECT  3.150 0.530 3.230 0.920 ;
        RECT  3.080 0.350 3.150 0.430 ;
        RECT  3.010 0.350 3.080 1.045 ;
        RECT  2.630 0.975 3.010 1.045 ;
        RECT  2.845 0.200 2.915 0.890 ;
        RECT  2.810 0.785 2.845 0.890 ;
        RECT  2.550 0.855 2.630 1.045 ;
        RECT  2.290 0.855 2.550 0.925 ;
        RECT  2.270 0.995 2.435 1.075 ;
        RECT  2.220 0.195 2.290 0.925 ;
        RECT  2.130 0.995 2.270 1.065 ;
        RECT  1.690 0.195 2.220 0.265 ;
        RECT  2.060 0.335 2.130 1.065 ;
        RECT  1.990 0.335 2.060 0.405 ;
        RECT  1.950 0.995 2.060 1.065 ;
        RECT  1.910 0.500 1.990 0.915 ;
        RECT  1.360 0.845 1.910 0.915 ;
        RECT  1.770 0.335 1.840 0.775 ;
        RECT  1.700 0.705 1.770 0.775 ;
        RECT  1.610 0.195 1.690 0.615 ;
        RECT  1.540 0.545 1.610 0.615 ;
        RECT  1.270 0.995 1.410 1.075 ;
        RECT  1.280 0.305 1.360 0.915 ;
        RECT  0.775 0.995 1.270 1.065 ;
        RECT  1.130 0.355 1.200 0.915 ;
        RECT  0.990 0.355 1.130 0.425 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.910 0.195 0.990 0.425 ;
        RECT  0.340 0.195 0.910 0.265 ;
        RECT  0.690 0.350 0.775 1.065 ;
        RECT  0.525 0.890 0.610 1.075 ;
        RECT  0.455 0.350 0.545 0.820 ;
        RECT  0.130 0.890 0.525 0.960 ;
        RECT  0.105 0.890 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D1BWP40

MACRO XNR4D2BWP40
    CLASS CORE ;
    FOREIGN XNR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.215 2.660 0.800 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.645 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.355 2.905 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.495 3.745 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.680 -0.115 3.920 0.115 ;
        RECT  3.610 -0.115 3.680 0.415 ;
        RECT  2.850 -0.115 3.610 0.115 ;
        RECT  2.750 -0.115 2.850 0.275 ;
        RECT  2.470 -0.115 2.750 0.115 ;
        RECT  2.380 -0.115 2.470 0.295 ;
        RECT  1.540 -0.115 2.380 0.115 ;
        RECT  1.470 -0.115 1.540 0.430 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.670 1.145 3.920 1.375 ;
        RECT  3.570 0.990 3.670 1.375 ;
        RECT  2.860 1.145 3.570 1.375 ;
        RECT  2.740 1.115 2.860 1.375 ;
        RECT  2.490 1.145 2.740 1.375 ;
        RECT  2.345 1.115 2.490 1.375 ;
        RECT  1.580 1.145 2.345 1.375 ;
        RECT  1.500 0.985 1.580 1.375 ;
        RECT  1.230 1.145 1.500 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.815 0.290 3.885 1.015 ;
        RECT  3.795 0.290 3.815 0.430 ;
        RECT  3.795 0.850 3.815 1.015 ;
        RECT  3.370 0.850 3.795 0.920 ;
        RECT  3.470 0.200 3.540 0.660 ;
        RECT  3.055 0.200 3.470 0.270 ;
        RECT  3.290 0.530 3.370 0.920 ;
        RECT  3.220 0.350 3.290 0.430 ;
        RECT  3.150 0.350 3.220 1.045 ;
        RECT  2.475 0.975 3.150 1.045 ;
        RECT  2.985 0.200 3.055 0.890 ;
        RECT  2.950 0.785 2.985 0.890 ;
        RECT  2.405 0.385 2.475 1.045 ;
        RECT  2.290 0.385 2.405 0.460 ;
        RECT  2.190 0.895 2.405 1.045 ;
        RECT  2.120 0.560 2.335 0.680 ;
        RECT  2.210 0.195 2.290 0.460 ;
        RECT  1.690 0.195 2.210 0.265 ;
        RECT  2.050 0.335 2.120 1.065 ;
        RECT  1.940 0.335 2.050 0.405 ;
        RECT  1.900 0.995 2.050 1.065 ;
        RECT  1.905 0.500 1.975 0.915 ;
        RECT  1.380 0.845 1.905 0.915 ;
        RECT  1.760 0.345 1.830 0.775 ;
        RECT  1.620 0.705 1.760 0.775 ;
        RECT  1.610 0.195 1.690 0.630 ;
        RECT  1.540 0.520 1.610 0.630 ;
        RECT  1.270 0.995 1.410 1.075 ;
        RECT  1.290 0.305 1.380 0.915 ;
        RECT  0.775 0.995 1.270 1.065 ;
        RECT  1.130 0.355 1.200 0.915 ;
        RECT  0.990 0.355 1.130 0.425 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.910 0.195 0.990 0.425 ;
        RECT  0.340 0.195 0.910 0.265 ;
        RECT  0.690 0.350 0.775 1.065 ;
        RECT  0.525 0.890 0.610 1.075 ;
        RECT  0.455 0.350 0.545 0.820 ;
        RECT  0.130 0.890 0.525 0.960 ;
        RECT  0.105 0.890 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D2BWP40

MACRO XNR4D4BWP40
    CLASS CORE ;
    FOREIGN XNR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.180 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN ZN
        ANTENNADIFFAREA 0.234000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.720 3.955 0.850 ;
        RECT  3.845 0.195 3.945 0.490 ;
        RECT  3.815 0.355 3.845 0.490 ;
        RECT  3.605 0.355 3.815 0.850 ;
        RECT  3.555 0.355 3.605 0.490 ;
        RECT  3.480 0.720 3.605 0.850 ;
        RECT  3.480 0.195 3.555 0.490 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.645 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.495 1.405 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.090 0.355 4.190 0.700 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.915 0.495 5.005 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.940 -0.115 5.180 0.115 ;
        RECT  4.870 -0.115 4.940 0.415 ;
        RECT  4.145 -0.115 4.870 0.115 ;
        RECT  4.030 -0.115 4.145 0.270 ;
        RECT  3.750 -0.115 4.030 0.115 ;
        RECT  3.660 -0.115 3.750 0.270 ;
        RECT  3.385 -0.115 3.660 0.115 ;
        RECT  3.280 -0.115 3.385 0.260 ;
        RECT  2.465 -0.115 3.280 0.115 ;
        RECT  2.395 -0.115 2.465 0.430 ;
        RECT  1.920 -0.115 2.395 0.115 ;
        RECT  1.830 -0.115 1.920 0.440 ;
        RECT  1.545 -0.115 1.830 0.115 ;
        RECT  1.445 -0.115 1.545 0.275 ;
        RECT  0.730 -0.115 1.445 0.115 ;
        RECT  0.600 -0.115 0.730 0.125 ;
        RECT  0.270 -0.115 0.600 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 1.145 5.180 1.375 ;
        RECT  4.830 0.990 4.930 1.375 ;
        RECT  4.140 1.145 4.830 1.375 ;
        RECT  4.020 1.115 4.140 1.375 ;
        RECT  3.770 1.145 4.020 1.375 ;
        RECT  3.625 1.115 3.770 1.375 ;
        RECT  3.390 1.145 3.625 1.375 ;
        RECT  3.245 1.115 3.390 1.375 ;
        RECT  2.475 1.145 3.245 1.375 ;
        RECT  2.395 0.985 2.475 1.375 ;
        RECT  1.915 1.145 2.395 1.375 ;
        RECT  1.835 0.985 1.915 1.375 ;
        RECT  1.585 1.145 1.835 1.375 ;
        RECT  1.465 1.135 1.585 1.375 ;
        RECT  0.740 1.145 1.465 1.375 ;
        RECT  0.620 1.030 0.740 1.375 ;
        RECT  0.340 1.145 0.620 1.375 ;
        RECT  0.220 1.030 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.885 0.720 3.955 0.850 ;
        RECT  3.885 0.195 3.945 0.490 ;
        RECT  3.480 0.195 3.535 0.490 ;
        RECT  3.480 0.720 3.535 0.850 ;
        RECT  5.075 0.290 5.145 1.015 ;
        RECT  5.055 0.290 5.075 0.430 ;
        RECT  5.055 0.850 5.075 1.015 ;
        RECT  4.640 0.850 5.055 0.920 ;
        RECT  4.730 0.200 4.800 0.660 ;
        RECT  4.335 0.200 4.730 0.270 ;
        RECT  4.560 0.530 4.640 0.920 ;
        RECT  4.490 0.350 4.560 0.430 ;
        RECT  4.420 0.350 4.490 1.045 ;
        RECT  3.410 0.975 4.420 1.045 ;
        RECT  4.260 0.200 4.335 0.890 ;
        RECT  4.220 0.785 4.260 0.890 ;
        RECT  3.340 0.385 3.410 1.045 ;
        RECT  3.185 0.385 3.340 0.460 ;
        RECT  3.105 0.895 3.340 1.045 ;
        RECT  3.035 0.560 3.240 0.680 ;
        RECT  3.105 0.195 3.185 0.460 ;
        RECT  2.605 0.195 3.105 0.265 ;
        RECT  2.960 0.335 3.035 1.065 ;
        RECT  2.835 0.335 2.960 0.405 ;
        RECT  2.795 0.995 2.960 1.065 ;
        RECT  2.820 0.500 2.890 0.915 ;
        RECT  2.105 0.845 2.820 0.915 ;
        RECT  2.675 0.345 2.750 0.775 ;
        RECT  2.275 0.705 2.675 0.775 ;
        RECT  2.535 0.195 2.605 0.630 ;
        RECT  2.400 0.520 2.535 0.630 ;
        RECT  2.185 0.305 2.275 0.775 ;
        RECT  2.025 0.255 2.105 0.915 ;
        RECT  1.725 0.845 2.025 0.915 ;
        RECT  1.630 0.995 1.755 1.075 ;
        RECT  1.645 0.260 1.725 0.915 ;
        RECT  1.130 0.995 1.630 1.065 ;
        RECT  1.485 0.355 1.560 0.915 ;
        RECT  1.345 0.355 1.485 0.425 ;
        RECT  1.245 0.845 1.485 0.915 ;
        RECT  1.265 0.195 1.345 0.425 ;
        RECT  0.390 0.195 1.265 0.265 ;
        RECT  1.045 0.350 1.130 1.065 ;
        RECT  0.895 0.890 0.965 1.075 ;
        RECT  0.825 0.350 0.900 0.820 ;
        RECT  0.130 0.890 0.895 0.960 ;
        RECT  0.545 0.730 0.825 0.820 ;
        RECT  0.455 0.350 0.545 0.820 ;
        RECT  0.105 0.890 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XNR4D4BWP40

MACRO XOR2D0BWP40
    CLASS CORE ;
    FOREIGN XOR2D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.046000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.215 1.505 1.045 ;
        RECT  1.420 0.215 1.435 0.435 ;
        RECT  1.420 0.895 1.435 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.355 1.225 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 -0.115 1.540 0.115 ;
        RECT  1.185 -0.115 1.265 0.275 ;
        RECT  0.270 -0.115 1.185 0.115 ;
        RECT  0.270 0.345 0.340 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.150 1.135 1.300 1.375 ;
        RECT  0.340 1.145 1.150 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.520 1.365 0.810 ;
        RECT  1.235 0.740 1.295 0.810 ;
        RECT  1.165 0.740 1.235 1.065 ;
        RECT  0.805 0.995 1.165 1.065 ;
        RECT  0.950 0.195 1.020 0.925 ;
        RECT  0.340 0.195 0.950 0.265 ;
        RECT  0.725 0.350 0.805 1.065 ;
        RECT  0.545 0.860 0.635 1.070 ;
        RECT  0.465 0.355 0.565 0.790 ;
        RECT  0.125 0.860 0.545 0.930 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.280 0.120 0.420 ;
        RECT  0.035 0.280 0.105 1.040 ;
    END
END XOR2D0BWP40

MACRO XOR2D1BWP40
    CLASS CORE ;
    FOREIGN XOR2D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.540 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.089700 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.195 1.505 1.045 ;
        RECT  1.415 0.195 1.435 0.460 ;
        RECT  1.420 0.895 1.435 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.355 1.225 0.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.385 0.640 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 -0.115 1.540 0.115 ;
        RECT  1.185 -0.115 1.265 0.275 ;
        RECT  0.270 -0.115 1.185 0.115 ;
        RECT  0.270 0.345 0.340 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.145 1.540 1.375 ;
        RECT  1.150 1.135 1.300 1.375 ;
        RECT  0.340 1.145 1.150 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.295 0.520 1.365 0.810 ;
        RECT  1.235 0.740 1.295 0.810 ;
        RECT  1.165 0.740 1.235 1.065 ;
        RECT  0.805 0.995 1.165 1.065 ;
        RECT  0.950 0.195 1.020 0.925 ;
        RECT  0.340 0.195 0.950 0.265 ;
        RECT  0.725 0.350 0.805 1.065 ;
        RECT  0.545 0.860 0.635 1.070 ;
        RECT  0.465 0.355 0.565 0.790 ;
        RECT  0.125 0.860 0.545 0.930 ;
        RECT  0.105 0.860 0.125 1.040 ;
        RECT  0.105 0.280 0.120 0.420 ;
        RECT  0.035 0.280 0.105 1.040 ;
    END
END XOR2D1BWP40

MACRO XOR2D2BWP40
    CLASS CORE ;
    FOREIGN XOR2D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.117000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 0.355 1.925 0.790 ;
        RECT  1.695 0.355 1.835 0.460 ;
        RECT  1.695 0.690 1.835 0.790 ;
        RECT  1.625 0.195 1.695 0.460 ;
        RECT  1.625 0.690 1.695 1.045 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.245 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.495 1.395 0.765 ;
        RECT  1.155 0.635 1.295 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 -0.115 1.960 0.115 ;
        RECT  1.800 -0.115 1.900 0.275 ;
        RECT  1.530 -0.115 1.800 0.115 ;
        RECT  1.435 -0.115 1.530 0.415 ;
        RECT  0.340 -0.115 1.435 0.115 ;
        RECT  0.220 -0.115 0.340 0.140 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.145 1.960 1.375 ;
        RECT  1.800 0.890 1.900 1.375 ;
        RECT  1.530 1.145 1.800 1.375 ;
        RECT  1.410 1.130 1.530 1.375 ;
        RECT  0.335 1.145 1.410 1.375 ;
        RECT  0.225 1.020 0.335 1.375 ;
        RECT  0.000 1.145 0.225 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.545 0.540 1.745 0.610 ;
        RECT  1.475 0.540 1.545 1.060 ;
        RECT  0.680 0.990 1.475 1.060 ;
        RECT  1.085 0.350 1.350 0.420 ;
        RECT  1.085 0.840 1.340 0.910 ;
        RECT  1.015 0.350 1.085 0.910 ;
        RECT  0.825 0.210 0.905 0.920 ;
        RECT  0.385 0.210 0.825 0.280 ;
        RECT  0.680 0.400 0.735 0.470 ;
        RECT  0.610 0.400 0.680 1.060 ;
        RECT  0.455 0.360 0.525 1.070 ;
        RECT  0.315 0.210 0.385 0.930 ;
        RECT  0.035 0.210 0.315 0.280 ;
        RECT  0.140 0.860 0.315 0.930 ;
        RECT  0.050 0.860 0.140 1.030 ;
    END
END XOR2D2BWP40

MACRO XOR2D3BWP40
    CLASS CORE ;
    FOREIGN XOR2D3BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.380 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.222300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.195 2.345 0.455 ;
        RECT  2.270 0.780 2.345 1.060 ;
        RECT  2.240 0.195 2.270 1.060 ;
        RECT  2.100 0.355 2.240 0.905 ;
        RECT  1.905 0.355 2.100 0.455 ;
        RECT  1.905 0.775 2.100 0.905 ;
        RECT  1.835 0.195 1.905 0.455 ;
        RECT  1.810 0.775 1.905 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.062400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.300 0.625 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.515 0.640 1.590 0.765 ;
        RECT  1.425 0.495 1.515 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 -0.115 2.380 0.115 ;
        RECT  2.020 -0.115 2.120 0.275 ;
        RECT  1.710 -0.115 2.020 0.115 ;
        RECT  1.625 -0.115 1.710 0.430 ;
        RECT  0.560 -0.115 1.625 0.115 ;
        RECT  0.440 -0.115 0.560 0.140 ;
        RECT  0.160 -0.115 0.440 0.115 ;
        RECT  0.060 -0.115 0.160 0.425 ;
        RECT  0.000 -0.115 0.060 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.145 2.380 1.375 ;
        RECT  2.020 0.985 2.120 1.375 ;
        RECT  1.730 1.145 2.020 1.375 ;
        RECT  1.610 1.130 1.730 1.375 ;
        RECT  0.545 1.145 1.610 1.375 ;
        RECT  0.435 0.840 0.545 1.375 ;
        RECT  0.160 1.145 0.435 1.375 ;
        RECT  0.060 0.855 0.160 1.375 ;
        RECT  0.000 1.145 0.060 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 0.540 1.965 0.620 ;
        RECT  1.670 0.540 1.740 1.060 ;
        RECT  0.890 0.990 1.670 1.060 ;
        RECT  1.320 0.310 1.550 0.400 ;
        RECT  1.320 0.850 1.550 0.920 ;
        RECT  1.250 0.310 1.320 0.920 ;
        RECT  1.060 0.210 1.140 0.920 ;
        RECT  0.575 0.210 1.060 0.280 ;
        RECT  0.680 0.360 0.750 0.970 ;
        RECT  0.665 0.360 0.680 0.480 ;
        RECT  0.665 0.800 0.680 0.970 ;
        RECT  0.575 0.510 0.600 0.640 ;
        RECT  0.505 0.210 0.575 0.765 ;
        RECT  0.265 0.210 0.505 0.370 ;
        RECT  0.360 0.695 0.505 0.765 ;
        RECT  0.270 0.695 0.360 1.075 ;
        RECT  0.890 0.400 0.980 0.470 ;
        RECT  0.820 0.400 0.890 1.060 ;
    END
END XOR2D3BWP40

MACRO XOR2D4BWP40
    CLASS CORE ;
    FOREIGN XOR2D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.940 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.231000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.205 2.695 1.065 ;
        RECT  2.615 0.355 2.625 1.065 ;
        RECT  2.485 0.355 2.615 0.915 ;
        RECT  2.315 0.355 2.485 0.485 ;
        RECT  2.315 0.780 2.485 0.915 ;
        RECT  2.245 0.205 2.315 0.485 ;
        RECT  2.245 0.780 2.315 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.061600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.495 0.340 0.645 ;
        RECT  0.035 0.495 0.105 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.965 0.665 2.020 0.765 ;
        RECT  1.855 0.495 1.965 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 -0.115 2.940 0.115 ;
        RECT  2.800 -0.115 2.900 0.480 ;
        RECT  2.520 -0.115 2.800 0.115 ;
        RECT  2.420 -0.115 2.520 0.285 ;
        RECT  2.125 -0.115 2.420 0.115 ;
        RECT  2.045 -0.115 2.125 0.450 ;
        RECT  0.910 -0.115 2.045 0.115 ;
        RECT  0.790 -0.115 0.910 0.140 ;
        RECT  0.530 -0.115 0.790 0.115 ;
        RECT  0.410 -0.115 0.530 0.140 ;
        RECT  0.135 -0.115 0.410 0.115 ;
        RECT  0.050 -0.115 0.135 0.355 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.145 2.940 1.375 ;
        RECT  2.800 0.695 2.900 1.375 ;
        RECT  2.530 1.145 2.800 1.375 ;
        RECT  2.410 0.995 2.530 1.375 ;
        RECT  2.140 1.145 2.410 1.375 ;
        RECT  2.020 1.130 2.140 1.375 ;
        RECT  0.910 1.145 2.020 1.375 ;
        RECT  0.790 1.005 0.910 1.375 ;
        RECT  0.530 1.145 0.790 1.375 ;
        RECT  0.410 1.050 0.530 1.375 ;
        RECT  0.135 1.145 0.410 1.375 ;
        RECT  0.050 0.860 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.315 0.355 2.415 0.485 ;
        RECT  2.315 0.780 2.415 0.915 ;
        RECT  2.245 0.205 2.315 0.485 ;
        RECT  2.245 0.780 2.315 1.065 ;
        RECT  2.165 0.555 2.305 0.625 ;
        RECT  2.095 0.555 2.165 1.060 ;
        RECT  1.215 0.990 2.095 1.060 ;
        RECT  1.730 0.850 1.960 0.920 ;
        RECT  1.730 0.350 1.945 0.420 ;
        RECT  1.660 0.350 1.730 0.920 ;
        RECT  1.410 0.210 1.490 0.920 ;
        RECT  0.500 0.210 1.410 0.280 ;
        RECT  1.215 0.400 1.330 0.470 ;
        RECT  1.145 0.400 1.215 1.060 ;
        RECT  0.985 0.810 1.075 1.065 ;
        RECT  0.835 0.360 1.070 0.490 ;
        RECT  0.835 0.810 0.985 0.880 ;
        RECT  0.750 0.360 0.835 0.880 ;
        RECT  0.600 0.360 0.750 0.460 ;
        RECT  0.715 0.810 0.750 0.880 ;
        RECT  0.615 0.810 0.715 1.015 ;
        RECT  0.500 0.530 0.680 0.660 ;
        RECT  0.330 0.730 0.420 0.800 ;
        RECT  0.240 0.730 0.330 1.075 ;
        RECT  0.420 0.210 0.500 0.800 ;
        RECT  0.240 0.210 0.420 0.370 ;
    END
END XOR2D4BWP40

MACRO XOR2D6BWP40
    CLASS CORE ;
    FOREIGN XOR2D6BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.500 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.346500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.165 0.200 3.275 0.485 ;
        RECT  3.165 0.775 3.275 1.065 ;
        RECT  2.975 0.355 3.165 0.485 ;
        RECT  2.975 0.775 3.165 0.905 ;
        RECT  2.875 0.355 2.975 0.905 ;
        RECT  2.805 0.205 2.875 1.065 ;
        RECT  2.795 0.355 2.805 1.065 ;
        RECT  2.765 0.355 2.795 0.905 ;
        RECT  2.495 0.355 2.765 0.450 ;
        RECT  2.495 0.780 2.765 0.905 ;
        RECT  2.425 0.205 2.495 0.450 ;
        RECT  2.425 0.780 2.495 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.091200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.495 0.390 0.625 ;
        RECT  0.175 0.495 0.245 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.095 0.495 2.205 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 -0.115 3.500 0.115 ;
        RECT  3.360 -0.115 3.460 0.440 ;
        RECT  3.085 -0.115 3.360 0.115 ;
        RECT  2.975 -0.115 3.085 0.275 ;
        RECT  2.700 -0.115 2.975 0.115 ;
        RECT  2.600 -0.115 2.700 0.275 ;
        RECT  2.300 -0.115 2.600 0.115 ;
        RECT  2.225 -0.115 2.300 0.420 ;
        RECT  1.100 -0.115 2.225 0.115 ;
        RECT  0.980 -0.115 1.100 0.140 ;
        RECT  0.720 -0.115 0.980 0.115 ;
        RECT  0.600 -0.115 0.720 0.140 ;
        RECT  0.340 -0.115 0.600 0.115 ;
        RECT  0.220 -0.115 0.340 0.140 ;
        RECT  0.000 -0.115 0.220 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.460 1.145 3.500 1.375 ;
        RECT  3.360 0.705 3.460 1.375 ;
        RECT  3.090 1.145 3.360 1.375 ;
        RECT  2.970 1.005 3.090 1.375 ;
        RECT  2.700 1.145 2.970 1.375 ;
        RECT  2.600 0.985 2.700 1.375 ;
        RECT  2.320 1.145 2.600 1.375 ;
        RECT  2.200 1.130 2.320 1.375 ;
        RECT  1.100 1.145 2.200 1.375 ;
        RECT  0.980 1.050 1.100 1.375 ;
        RECT  0.720 1.145 0.980 1.375 ;
        RECT  0.600 1.050 0.720 1.375 ;
        RECT  0.340 1.145 0.600 1.375 ;
        RECT  0.220 1.050 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.165 0.200 3.275 0.485 ;
        RECT  3.165 0.775 3.275 1.065 ;
        RECT  3.045 0.355 3.165 0.485 ;
        RECT  3.045 0.775 3.165 0.905 ;
        RECT  2.495 0.355 2.695 0.450 ;
        RECT  2.495 0.780 2.695 0.905 ;
        RECT  2.425 0.205 2.495 0.450 ;
        RECT  2.425 0.780 2.495 1.065 ;
        RECT  2.345 0.520 2.605 0.610 ;
        RECT  2.275 0.520 2.345 1.060 ;
        RECT  2.090 0.990 2.275 1.060 ;
        RECT  1.910 0.850 2.140 0.920 ;
        RECT  1.910 0.350 2.125 0.420 ;
        RECT  2.020 0.990 2.090 1.065 ;
        RECT  1.455 0.995 2.020 1.065 ;
        RECT  1.840 0.350 1.910 0.920 ;
        RECT  1.650 0.220 1.730 0.925 ;
        RECT  0.660 0.220 1.650 0.290 ;
        RECT  1.455 0.400 1.570 0.470 ;
        RECT  1.385 0.400 1.455 1.065 ;
        RECT  1.210 0.360 1.290 0.930 ;
        RECT  0.785 0.360 1.210 0.440 ;
        RECT  0.785 0.850 1.210 0.930 ;
        RECT  0.660 0.510 0.890 0.640 ;
        RECT  0.590 0.220 0.660 0.980 ;
        RECT  0.050 0.220 0.590 0.340 ;
        RECT  0.150 0.885 0.590 0.980 ;
        RECT  0.050 0.845 0.150 0.980 ;
    END
END XOR2D6BWP40

MACRO XOR2D8BWP40
    CLASS CORE ;
    FOREIGN XOR2D8BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.468000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.305 0.205 4.375 0.485 ;
        RECT  4.305 0.780 4.375 1.065 ;
        RECT  3.995 0.355 4.305 0.485 ;
        RECT  4.005 0.780 4.305 0.905 ;
        RECT  3.925 0.780 4.005 1.065 ;
        RECT  3.925 0.205 3.995 0.485 ;
        RECT  3.815 0.355 3.925 0.485 ;
        RECT  3.815 0.780 3.925 0.905 ;
        RECT  3.610 0.355 3.815 0.905 ;
        RECT  3.605 0.205 3.610 1.065 ;
        RECT  3.540 0.205 3.605 0.480 ;
        RECT  3.535 0.780 3.605 1.065 ;
        RECT  3.230 0.355 3.540 0.480 ;
        RECT  3.230 0.780 3.535 0.905 ;
        RECT  3.160 0.195 3.230 0.480 ;
        RECT  3.160 0.780 3.230 1.065 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.124800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.495 0.665 0.770 ;
        RECT  0.310 0.495 0.595 0.625 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.048000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.800 0.495 2.915 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 -0.115 4.620 0.115 ;
        RECT  4.480 -0.115 4.580 0.485 ;
        RECT  4.200 -0.115 4.480 0.115 ;
        RECT  4.100 -0.115 4.200 0.275 ;
        RECT  3.820 -0.115 4.100 0.115 ;
        RECT  3.720 -0.115 3.820 0.275 ;
        RECT  3.435 -0.115 3.720 0.115 ;
        RECT  3.335 -0.115 3.435 0.275 ;
        RECT  3.035 -0.115 3.335 0.115 ;
        RECT  2.960 -0.115 3.035 0.415 ;
        RECT  1.650 -0.115 2.960 0.115 ;
        RECT  1.580 -0.115 1.650 0.275 ;
        RECT  1.295 -0.115 1.580 0.115 ;
        RECT  1.170 -0.115 1.295 0.245 ;
        RECT  0.910 -0.115 1.170 0.115 ;
        RECT  0.790 -0.115 0.910 0.215 ;
        RECT  0.535 -0.115 0.790 0.115 ;
        RECT  0.405 -0.115 0.535 0.240 ;
        RECT  0.135 -0.115 0.405 0.115 ;
        RECT  0.050 -0.115 0.135 0.495 ;
        RECT  0.000 -0.115 0.050 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 1.145 4.620 1.375 ;
        RECT  4.480 0.695 4.580 1.375 ;
        RECT  4.200 1.145 4.480 1.375 ;
        RECT  4.100 0.985 4.200 1.375 ;
        RECT  3.820 1.145 4.100 1.375 ;
        RECT  3.720 0.985 3.820 1.375 ;
        RECT  3.435 1.145 3.720 1.375 ;
        RECT  3.335 0.985 3.435 1.375 ;
        RECT  3.055 1.145 3.335 1.375 ;
        RECT  2.935 1.130 3.055 1.375 ;
        RECT  1.670 1.145 2.935 1.375 ;
        RECT  1.560 0.980 1.670 1.375 ;
        RECT  1.285 1.145 1.560 1.375 ;
        RECT  1.175 0.980 1.285 1.375 ;
        RECT  0.905 1.145 1.175 1.375 ;
        RECT  0.795 1.025 0.905 1.375 ;
        RECT  0.535 1.145 0.795 1.375 ;
        RECT  0.405 1.045 0.535 1.375 ;
        RECT  0.135 1.145 0.405 1.375 ;
        RECT  0.050 0.720 0.135 1.375 ;
        RECT  0.000 1.145 0.050 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.305 0.205 4.375 0.485 ;
        RECT  4.305 0.780 4.375 1.065 ;
        RECT  3.995 0.355 4.305 0.485 ;
        RECT  4.005 0.780 4.305 0.905 ;
        RECT  3.925 0.780 4.005 1.065 ;
        RECT  3.925 0.205 3.995 0.485 ;
        RECT  3.885 0.355 3.925 0.485 ;
        RECT  3.885 0.780 3.925 0.905 ;
        RECT  3.230 0.355 3.535 0.480 ;
        RECT  3.230 0.780 3.535 0.905 ;
        RECT  3.160 0.195 3.230 0.480 ;
        RECT  3.160 0.780 3.230 1.065 ;
        RECT  3.080 0.550 3.495 0.625 ;
        RECT  3.010 0.550 3.080 1.060 ;
        RECT  2.555 0.990 3.010 1.060 ;
        RECT  2.705 0.850 2.875 0.920 ;
        RECT  2.705 0.350 2.855 0.420 ;
        RECT  2.635 0.350 2.705 0.920 ;
        RECT  2.555 0.195 2.685 0.265 ;
        RECT  2.485 0.195 2.555 1.060 ;
        RECT  1.735 0.195 2.485 0.265 ;
        RECT  1.740 0.990 2.485 1.060 ;
        RECT  2.325 0.340 2.405 0.920 ;
        RECT  1.350 0.535 2.325 0.605 ;
        RECT  1.230 0.360 2.045 0.430 ;
        RECT  1.230 0.810 2.045 0.880 ;
        RECT  1.145 0.360 1.230 0.880 ;
        RECT  0.975 0.360 1.145 0.430 ;
        RECT  0.975 0.810 1.145 0.880 ;
        RECT  0.855 0.530 1.065 0.620 ;
        RECT  0.775 0.310 0.855 0.955 ;
        RECT  0.320 0.310 0.775 0.380 ;
        RECT  0.220 0.885 0.775 0.955 ;
        RECT  0.250 0.220 0.320 0.380 ;
    END
END XOR2D8BWP40

MACRO XOR3D0BWP40
    CLASS CORE ;
    FOREIGN XOR3D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.050000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.185 2.625 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.285 0.215 2.345 0.485 ;
        RECT  2.205 0.215 2.285 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.120 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 -0.115 2.660 0.115 ;
        RECT  2.275 -0.115 2.395 0.130 ;
        RECT  1.520 -0.115 2.275 0.115 ;
        RECT  1.450 -0.115 1.520 0.465 ;
        RECT  1.170 -0.115 1.450 0.115 ;
        RECT  1.070 -0.115 1.170 0.415 ;
        RECT  0.320 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.320 0.330 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 1.145 2.660 1.375 ;
        RECT  2.275 1.135 2.395 1.375 ;
        RECT  1.620 1.145 2.275 1.375 ;
        RECT  1.540 0.845 1.620 1.375 ;
        RECT  1.430 0.845 1.540 0.915 ;
        RECT  1.210 1.145 1.540 1.375 ;
        RECT  1.090 1.135 1.210 1.375 ;
        RECT  0.340 1.145 1.090 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.395 0.535 2.465 1.055 ;
        RECT  1.970 0.985 2.395 1.055 ;
        RECT  2.120 0.785 2.175 0.905 ;
        RECT  2.050 0.205 2.120 0.905 ;
        RECT  1.670 0.205 2.050 0.275 ;
        RECT  1.900 0.365 1.970 1.055 ;
        RECT  1.780 0.365 1.900 0.435 ;
        RECT  1.850 0.850 1.900 1.055 ;
        RECT  1.750 0.520 1.830 0.765 ;
        RECT  1.365 0.695 1.750 0.765 ;
        RECT  1.590 0.205 1.670 0.615 ;
        RECT  1.480 0.545 1.590 0.615 ;
        RECT  0.790 0.995 1.460 1.065 ;
        RECT  1.360 0.295 1.365 0.765 ;
        RECT  1.295 0.295 1.360 0.900 ;
        RECT  1.265 0.295 1.295 0.435 ;
        RECT  1.260 0.715 1.295 0.900 ;
        RECT  0.870 0.195 0.940 0.915 ;
        RECT  0.495 0.195 0.870 0.265 ;
        RECT  0.715 0.335 0.790 1.065 ;
        RECT  0.640 0.335 0.715 0.415 ;
        RECT  0.670 0.915 0.715 1.065 ;
        RECT  0.565 0.535 0.645 0.835 ;
        RECT  0.445 0.765 0.565 0.835 ;
        RECT  0.425 0.195 0.495 0.640 ;
        RECT  0.355 0.765 0.445 0.930 ;
        RECT  0.365 0.515 0.425 0.640 ;
        RECT  0.130 0.860 0.355 0.930 ;
        RECT  0.105 0.195 0.130 0.355 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END XOR3D0BWP40

MACRO XOR3D1BWP40
    CLASS CORE ;
    FOREIGN XOR3D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.093125 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.535 0.185 2.625 1.045 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.029800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.285 0.215 2.345 0.485 ;
        RECT  2.205 0.215 2.285 0.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.265 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.495 1.130 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 -0.115 2.660 0.115 ;
        RECT  2.275 -0.115 2.395 0.130 ;
        RECT  1.520 -0.115 2.275 0.115 ;
        RECT  1.450 -0.115 1.520 0.465 ;
        RECT  1.170 -0.115 1.450 0.115 ;
        RECT  1.070 -0.115 1.170 0.415 ;
        RECT  0.320 -0.115 1.070 0.115 ;
        RECT  0.240 -0.115 0.320 0.330 ;
        RECT  0.000 -0.115 0.240 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 1.145 2.660 1.375 ;
        RECT  2.275 1.135 2.395 1.375 ;
        RECT  1.620 1.145 2.275 1.375 ;
        RECT  1.540 0.845 1.620 1.375 ;
        RECT  1.430 0.845 1.540 0.915 ;
        RECT  1.210 1.145 1.540 1.375 ;
        RECT  1.090 1.135 1.210 1.375 ;
        RECT  0.340 1.145 1.090 1.375 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.395 0.535 2.465 1.055 ;
        RECT  1.970 0.985 2.395 1.055 ;
        RECT  2.120 0.785 2.175 0.905 ;
        RECT  2.050 0.205 2.120 0.905 ;
        RECT  1.670 0.205 2.050 0.275 ;
        RECT  1.900 0.365 1.970 1.055 ;
        RECT  1.780 0.365 1.900 0.435 ;
        RECT  1.850 0.850 1.900 1.055 ;
        RECT  1.750 0.520 1.830 0.765 ;
        RECT  1.365 0.695 1.750 0.765 ;
        RECT  1.590 0.205 1.670 0.615 ;
        RECT  1.480 0.545 1.590 0.615 ;
        RECT  0.790 0.995 1.460 1.065 ;
        RECT  1.360 0.295 1.365 0.765 ;
        RECT  1.295 0.295 1.360 0.900 ;
        RECT  1.265 0.295 1.295 0.435 ;
        RECT  1.260 0.715 1.295 0.900 ;
        RECT  0.870 0.195 0.940 0.915 ;
        RECT  0.495 0.195 0.870 0.265 ;
        RECT  0.715 0.335 0.790 1.065 ;
        RECT  0.640 0.335 0.715 0.415 ;
        RECT  0.670 0.915 0.715 1.065 ;
        RECT  0.565 0.535 0.645 0.835 ;
        RECT  0.445 0.765 0.565 0.835 ;
        RECT  0.425 0.195 0.495 0.640 ;
        RECT  0.355 0.765 0.445 0.930 ;
        RECT  0.365 0.515 0.425 0.640 ;
        RECT  0.130 0.860 0.355 0.930 ;
        RECT  0.105 0.195 0.130 0.355 ;
        RECT  0.105 0.860 0.130 1.040 ;
        RECT  0.035 0.195 0.105 1.040 ;
    END
END XOR3D1BWP40

MACRO XOR3D2BWP40
    CLASS CORE ;
    FOREIGN XOR3D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.111750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.355 2.765 0.765 ;
        RECT  2.580 0.355 2.695 0.465 ;
        RECT  2.560 0.695 2.695 0.765 ;
        RECT  2.490 0.185 2.580 0.465 ;
        RECT  2.485 0.695 2.560 1.070 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.029800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.735 2.345 1.050 ;
        RECT  2.255 0.520 2.280 1.050 ;
        RECT  2.210 0.520 2.255 0.805 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.770 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.030200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.355 1.105 0.640 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.115 2.800 0.115 ;
        RECT  2.670 -0.115 2.750 0.280 ;
        RECT  2.390 -0.115 2.670 0.115 ;
        RECT  2.270 -0.115 2.390 0.140 ;
        RECT  1.560 -0.115 2.270 0.115 ;
        RECT  1.440 -0.115 1.560 0.265 ;
        RECT  1.165 -0.115 1.440 0.115 ;
        RECT  1.085 -0.115 1.165 0.285 ;
        RECT  0.260 -0.115 1.085 0.115 ;
        RECT  0.260 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.260 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 1.145 2.800 1.375 ;
        RECT  2.670 0.855 2.750 1.375 ;
        RECT  2.390 1.145 2.670 1.375 ;
        RECT  2.270 1.120 2.390 1.375 ;
        RECT  1.545 1.145 2.270 1.375 ;
        RECT  1.460 0.780 1.545 1.375 ;
        RECT  1.215 1.145 1.460 1.375 ;
        RECT  1.095 1.135 1.215 1.375 ;
        RECT  0.340 1.145 1.095 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.420 0.545 2.600 0.615 ;
        RECT  2.350 0.210 2.420 0.615 ;
        RECT  1.990 0.210 2.350 0.280 ;
        RECT  2.140 0.360 2.220 0.430 ;
        RECT  2.140 0.885 2.170 1.065 ;
        RECT  2.070 0.360 2.140 1.065 ;
        RECT  1.720 0.995 2.070 1.065 ;
        RECT  1.880 0.210 1.990 0.925 ;
        RECT  1.720 0.185 1.810 0.415 ;
        RECT  1.360 0.345 1.720 0.415 ;
        RECT  1.640 0.560 1.720 1.065 ;
        RECT  1.510 0.560 1.640 0.635 ;
        RECT  1.280 0.345 1.360 0.900 ;
        RECT  0.765 0.995 1.360 1.065 ;
        RECT  0.945 0.855 0.970 0.925 ;
        RECT  0.860 0.195 0.945 0.925 ;
        RECT  0.340 0.195 0.860 0.265 ;
        RECT  0.695 0.345 0.765 1.065 ;
        RECT  0.560 0.995 0.625 1.065 ;
        RECT  0.490 0.870 0.560 1.065 ;
        RECT  0.125 0.870 0.490 0.940 ;
        RECT  0.105 0.870 0.125 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR3D2BWP40

MACRO XOR3D4BWP40
    CLASS CORE ;
    FOREIGN XOR3D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.228000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.605 0.195 3.675 0.465 ;
        RECT  3.605 0.745 3.675 1.065 ;
        RECT  3.535 0.355 3.605 0.465 ;
        RECT  3.535 0.745 3.605 0.905 ;
        RECT  3.325 0.355 3.535 0.905 ;
        RECT  3.295 0.355 3.325 0.465 ;
        RECT  3.295 0.745 3.325 0.905 ;
        RECT  3.225 0.195 3.295 0.465 ;
        RECT  3.225 0.745 3.295 1.065 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.495 2.775 0.630 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.031400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.635 0.385 0.765 ;
        RECT  0.175 0.555 0.260 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.060800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.355 1.085 0.630 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 -0.115 3.920 0.115 ;
        RECT  3.795 -0.115 3.875 0.485 ;
        RECT  3.500 -0.115 3.795 0.115 ;
        RECT  3.400 -0.115 3.500 0.275 ;
        RECT  3.130 -0.115 3.400 0.115 ;
        RECT  3.010 -0.115 3.130 0.140 ;
        RECT  2.760 -0.115 3.010 0.115 ;
        RECT  2.630 -0.115 2.760 0.140 ;
        RECT  2.020 -0.115 2.630 0.115 ;
        RECT  1.890 -0.115 2.020 0.140 ;
        RECT  1.130 -0.115 1.890 0.115 ;
        RECT  1.030 -0.115 1.130 0.270 ;
        RECT  0.260 -0.115 1.030 0.115 ;
        RECT  0.260 0.380 0.360 0.450 ;
        RECT  0.190 -0.115 0.260 0.450 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.875 1.145 3.920 1.375 ;
        RECT  3.795 0.755 3.875 1.375 ;
        RECT  3.500 1.145 3.795 1.375 ;
        RECT  3.400 0.985 3.500 1.375 ;
        RECT  3.120 1.145 3.400 1.375 ;
        RECT  3.020 1.010 3.120 1.375 ;
        RECT  2.750 1.145 3.020 1.375 ;
        RECT  2.650 1.010 2.750 1.375 ;
        RECT  2.000 1.145 2.650 1.375 ;
        RECT  1.900 0.990 2.000 1.375 ;
        RECT  1.130 1.145 1.900 1.375 ;
        RECT  1.030 1.010 1.130 1.375 ;
        RECT  0.340 1.145 1.030 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.605 0.195 3.675 0.465 ;
        RECT  3.605 0.745 3.675 1.065 ;
        RECT  3.225 0.195 3.255 0.465 ;
        RECT  3.225 0.745 3.255 1.065 ;
        RECT  3.130 0.545 3.255 0.615 ;
        RECT  3.060 0.210 3.130 0.940 ;
        RECT  1.450 0.210 3.060 0.280 ;
        RECT  2.540 0.870 3.060 0.940 ;
        RECT  2.925 0.730 2.960 0.800 ;
        RECT  2.855 0.350 2.925 0.800 ;
        RECT  2.460 0.730 2.855 0.800 ;
        RECT  2.460 0.350 2.585 0.425 ;
        RECT  2.470 0.870 2.540 1.065 ;
        RECT  2.240 0.995 2.470 1.065 ;
        RECT  2.390 0.350 2.460 0.800 ;
        RECT  2.350 0.730 2.390 0.800 ;
        RECT  2.280 0.730 2.350 0.920 ;
        RECT  2.200 0.545 2.320 0.615 ;
        RECT  1.960 0.850 2.280 0.920 ;
        RECT  2.120 0.350 2.200 0.780 ;
        RECT  2.105 0.350 2.120 0.520 ;
        RECT  2.075 0.710 2.120 0.780 ;
        RECT  1.670 0.450 2.105 0.520 ;
        RECT  1.890 0.590 1.960 0.920 ;
        RECT  1.820 0.590 1.890 0.660 ;
        RECT  1.580 0.360 1.670 0.520 ;
        RECT  1.505 0.980 1.665 1.075 ;
        RECT  1.450 0.805 1.520 0.875 ;
        RECT  1.300 0.980 1.505 1.050 ;
        RECT  1.380 0.210 1.450 0.875 ;
        RECT  1.220 0.195 1.310 0.785 ;
        RECT  1.230 0.855 1.300 1.050 ;
        RECT  0.740 0.855 1.230 0.925 ;
        RECT  0.910 0.705 1.220 0.785 ;
        RECT  0.830 0.195 0.910 0.785 ;
        RECT  0.430 0.195 0.830 0.265 ;
        RECT  0.620 0.345 0.740 0.925 ;
        RECT  0.520 0.995 0.640 1.065 ;
        RECT  0.450 0.870 0.520 1.065 ;
        RECT  0.125 0.870 0.450 0.940 ;
        RECT  0.330 0.195 0.430 0.305 ;
        RECT  0.105 0.870 0.125 1.050 ;
        RECT  0.105 0.325 0.120 0.445 ;
        RECT  0.035 0.325 0.105 1.050 ;
    END
END XOR3D4BWP40

MACRO XOR4D0BWP40
    CLASS CORE ;
    FOREIGN XOR4D0BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.082500 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.355 2.485 0.905 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.016000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.440 2.790 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.495 0.495 3.605 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.780 0.115 ;
        RECT  3.520 -0.115 3.590 0.415 ;
        RECT  2.670 -0.115 3.520 0.115 ;
        RECT  3.420 0.345 3.520 0.415 ;
        RECT  2.540 -0.115 2.670 0.140 ;
        RECT  1.540 -0.115 2.540 0.115 ;
        RECT  1.470 -0.115 1.540 0.460 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.145 3.780 1.375 ;
        RECT  3.440 1.010 3.560 1.375 ;
        RECT  2.710 1.145 3.440 1.375 ;
        RECT  2.590 1.120 2.710 1.375 ;
        RECT  1.590 1.145 2.590 1.375 ;
        RECT  1.470 0.995 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.300 3.745 1.050 ;
        RECT  3.660 0.300 3.675 0.440 ;
        RECT  3.650 0.870 3.675 1.050 ;
        RECT  3.260 0.870 3.650 0.940 ;
        RECT  2.940 0.195 3.450 0.265 ;
        RECT  3.160 0.870 3.260 1.070 ;
        RECT  3.090 0.710 3.160 0.790 ;
        RECT  3.020 0.345 3.090 1.050 ;
        RECT  3.010 0.345 3.020 0.535 ;
        RECT  2.625 0.980 3.020 1.050 ;
        RECT  2.870 0.195 2.940 0.910 ;
        RECT  2.780 0.195 2.870 0.360 ;
        RECT  2.760 0.840 2.870 0.910 ;
        RECT  2.555 0.210 2.625 1.050 ;
        RECT  1.680 0.210 2.555 0.280 ;
        RECT  2.270 0.980 2.555 1.050 ;
        RECT  2.120 0.510 2.285 0.630 ;
        RECT  2.200 0.890 2.270 1.050 ;
        RECT  2.050 0.360 2.120 1.065 ;
        RECT  1.910 0.360 2.050 0.440 ;
        RECT  1.910 0.995 2.050 1.065 ;
        RECT  1.900 0.520 1.980 0.925 ;
        RECT  1.360 0.855 1.900 0.925 ;
        RECT  1.760 0.360 1.830 0.785 ;
        RECT  1.660 0.715 1.760 0.785 ;
        RECT  1.610 0.210 1.680 0.640 ;
        RECT  1.270 0.995 1.390 1.075 ;
        RECT  1.280 0.325 1.360 0.925 ;
        RECT  0.795 0.995 1.270 1.065 ;
        RECT  1.130 0.345 1.200 0.915 ;
        RECT  0.990 0.345 1.130 0.415 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.910 0.195 0.990 0.415 ;
        RECT  0.340 0.195 0.910 0.265 ;
        RECT  0.695 0.350 0.795 1.065 ;
        RECT  0.520 0.870 0.600 1.070 ;
        RECT  0.455 0.350 0.545 0.800 ;
        RECT  0.130 0.870 0.520 0.940 ;
        RECT  0.420 0.720 0.455 0.800 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D0BWP40

MACRO XOR4D1BWP40
    CLASS CORE ;
    FOREIGN XOR4D1BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.780 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.111200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.355 2.485 0.905 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.765 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.440 2.790 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.500 0.495 3.605 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.590 -0.115 3.780 0.115 ;
        RECT  3.520 -0.115 3.590 0.415 ;
        RECT  2.670 -0.115 3.520 0.115 ;
        RECT  3.420 0.345 3.520 0.415 ;
        RECT  2.540 -0.115 2.670 0.140 ;
        RECT  1.540 -0.115 2.540 0.115 ;
        RECT  1.470 -0.115 1.540 0.460 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.145 3.780 1.375 ;
        RECT  3.440 1.010 3.560 1.375 ;
        RECT  2.710 1.145 3.440 1.375 ;
        RECT  2.590 1.120 2.710 1.375 ;
        RECT  1.590 1.145 2.590 1.375 ;
        RECT  1.470 0.995 1.590 1.375 ;
        RECT  1.230 1.145 1.470 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.675 0.300 3.745 1.050 ;
        RECT  3.660 0.300 3.675 0.440 ;
        RECT  3.650 0.870 3.675 1.050 ;
        RECT  3.260 0.870 3.650 0.940 ;
        RECT  2.940 0.195 3.450 0.265 ;
        RECT  3.160 0.870 3.260 1.070 ;
        RECT  3.090 0.710 3.160 0.790 ;
        RECT  3.020 0.345 3.090 1.050 ;
        RECT  3.010 0.345 3.020 0.535 ;
        RECT  2.625 0.980 3.020 1.050 ;
        RECT  2.870 0.195 2.940 0.910 ;
        RECT  2.780 0.195 2.870 0.360 ;
        RECT  2.760 0.840 2.870 0.910 ;
        RECT  2.555 0.210 2.625 1.050 ;
        RECT  1.680 0.210 2.555 0.280 ;
        RECT  2.270 0.980 2.555 1.050 ;
        RECT  2.120 0.510 2.285 0.630 ;
        RECT  2.200 0.890 2.270 1.050 ;
        RECT  2.050 0.360 2.120 1.065 ;
        RECT  1.910 0.360 2.050 0.440 ;
        RECT  1.910 0.995 2.050 1.065 ;
        RECT  1.900 0.520 1.980 0.925 ;
        RECT  1.360 0.855 1.900 0.925 ;
        RECT  1.760 0.360 1.830 0.785 ;
        RECT  1.660 0.715 1.760 0.785 ;
        RECT  1.610 0.210 1.680 0.640 ;
        RECT  1.270 0.995 1.390 1.075 ;
        RECT  1.280 0.185 1.360 0.925 ;
        RECT  0.795 0.995 1.270 1.065 ;
        RECT  1.130 0.345 1.200 0.915 ;
        RECT  0.990 0.345 1.130 0.415 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.910 0.195 0.990 0.415 ;
        RECT  0.340 0.195 0.910 0.265 ;
        RECT  0.695 0.350 0.795 1.065 ;
        RECT  0.520 0.870 0.600 1.070 ;
        RECT  0.455 0.350 0.545 0.800 ;
        RECT  0.130 0.870 0.520 0.940 ;
        RECT  0.420 0.720 0.455 0.800 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D1BWP40

MACRO XOR4D2BWP40
    CLASS CORE ;
    FOREIGN XOR4D2BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.114000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.625 0.700 2.665 0.770 ;
        RECT  2.555 0.195 2.625 0.770 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.031800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.031200 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 0.495 1.050 0.640 ;
        RECT  0.875 0.495 0.945 0.765 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.805 0.495 2.905 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.031800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 0.495 3.745 0.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 -0.115 3.920 0.115 ;
        RECT  3.650 -0.115 3.720 0.415 ;
        RECT  2.830 -0.115 3.650 0.115 ;
        RECT  3.570 0.345 3.650 0.415 ;
        RECT  2.750 -0.115 2.830 0.275 ;
        RECT  2.440 -0.115 2.750 0.115 ;
        RECT  2.360 -0.115 2.440 0.290 ;
        RECT  1.540 -0.115 2.360 0.115 ;
        RECT  1.470 -0.115 1.540 0.460 ;
        RECT  1.190 -0.115 1.470 0.115 ;
        RECT  1.090 -0.115 1.190 0.275 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.360 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.700 1.145 3.920 1.375 ;
        RECT  3.580 1.010 3.700 1.375 ;
        RECT  2.870 1.145 3.580 1.375 ;
        RECT  2.750 1.120 2.870 1.375 ;
        RECT  2.460 1.145 2.750 1.375 ;
        RECT  2.380 0.980 2.460 1.375 ;
        RECT  1.600 1.145 2.380 1.375 ;
        RECT  1.480 0.985 1.600 1.375 ;
        RECT  1.230 1.145 1.480 1.375 ;
        RECT  1.110 1.135 1.230 1.375 ;
        RECT  0.340 1.145 1.110 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.815 0.300 3.885 1.050 ;
        RECT  3.800 0.300 3.815 0.440 ;
        RECT  3.790 0.870 3.815 1.050 ;
        RECT  3.425 0.870 3.790 0.940 ;
        RECT  3.070 0.195 3.580 0.265 ;
        RECT  3.355 0.870 3.425 1.055 ;
        RECT  3.280 0.985 3.355 1.055 ;
        RECT  3.210 0.700 3.265 0.830 ;
        RECT  3.140 0.345 3.210 1.050 ;
        RECT  2.620 0.980 3.140 1.050 ;
        RECT  3.000 0.195 3.070 0.910 ;
        RECT  2.955 0.300 3.000 0.420 ;
        RECT  2.950 0.840 3.000 0.910 ;
        RECT  2.550 0.840 2.620 1.050 ;
        RECT  2.480 0.840 2.550 0.910 ;
        RECT  2.410 0.370 2.480 0.910 ;
        RECT  2.280 0.370 2.410 0.440 ;
        RECT  2.270 0.730 2.410 0.800 ;
        RECT  2.120 0.520 2.330 0.640 ;
        RECT  2.210 0.210 2.280 0.440 ;
        RECT  2.200 0.730 2.270 1.050 ;
        RECT  1.690 0.210 2.210 0.280 ;
        RECT  2.050 0.360 2.120 1.055 ;
        RECT  1.950 0.360 2.050 0.440 ;
        RECT  1.945 0.985 2.050 1.055 ;
        RECT  1.900 0.520 1.980 0.915 ;
        RECT  1.360 0.845 1.900 0.915 ;
        RECT  1.760 0.360 1.830 0.775 ;
        RECT  1.695 0.700 1.760 0.775 ;
        RECT  1.610 0.210 1.690 0.620 ;
        RECT  1.545 0.540 1.610 0.620 ;
        RECT  1.270 0.995 1.390 1.075 ;
        RECT  1.280 0.185 1.360 0.915 ;
        RECT  0.805 0.995 1.270 1.065 ;
        RECT  1.130 0.345 1.200 0.915 ;
        RECT  1.000 0.345 1.130 0.415 ;
        RECT  0.890 0.845 1.130 0.915 ;
        RECT  0.900 0.195 1.000 0.415 ;
        RECT  0.340 0.195 0.900 0.265 ;
        RECT  0.735 0.350 0.805 1.065 ;
        RECT  0.720 0.350 0.735 0.830 ;
        RECT  0.675 0.700 0.720 0.830 ;
        RECT  0.510 0.985 0.665 1.055 ;
        RECT  0.450 0.350 0.530 0.800 ;
        RECT  0.440 0.870 0.510 1.055 ;
        RECT  0.130 0.870 0.440 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D2BWP40

MACRO XOR4D4BWP40
    CLASS CORE ;
    FOREIGN XOR4D4BWP40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.620 BY 1.260 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Z
        ANTENNADIFFAREA 0.228000 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.195 0.805 3.305 1.075 ;
        RECT  3.115 0.355 3.285 0.485 ;
        RECT  3.115 0.805 3.195 0.905 ;
        RECT  2.925 0.355 3.115 0.905 ;
        RECT  2.905 0.355 2.925 1.075 ;
        RECT  2.815 0.355 2.905 0.480 ;
        RECT  2.820 0.805 2.905 1.075 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.031600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.175 0.495 0.275 0.770 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.029000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.495 1.225 0.765 ;
        RECT  1.030 0.495 1.135 0.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.030400 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.395 0.495 3.555 0.765 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.032000 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.360 0.495 4.445 0.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.390 -0.115 4.620 0.115 ;
        RECT  4.290 -0.115 4.390 0.315 ;
        RECT  3.510 -0.115 4.290 0.115 ;
        RECT  3.380 -0.115 3.510 0.140 ;
        RECT  3.120 -0.115 3.380 0.115 ;
        RECT  3.000 -0.115 3.120 0.140 ;
        RECT  2.730 -0.115 3.000 0.115 ;
        RECT  2.610 -0.115 2.730 0.140 ;
        RECT  2.360 -0.115 2.610 0.115 ;
        RECT  2.240 -0.115 2.360 0.140 ;
        RECT  1.550 -0.115 2.240 0.115 ;
        RECT  1.465 -0.115 1.550 0.440 ;
        RECT  1.190 -0.115 1.465 0.115 ;
        RECT  1.090 -0.115 1.190 0.420 ;
        RECT  0.270 -0.115 1.090 0.115 ;
        RECT  0.270 0.345 0.350 0.415 ;
        RECT  0.190 -0.115 0.270 0.415 ;
        RECT  0.000 -0.115 0.190 0.115 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.370 1.145 4.620 1.375 ;
        RECT  4.300 0.995 4.370 1.375 ;
        RECT  3.480 1.145 4.300 1.375 ;
        RECT  3.400 0.915 3.480 1.375 ;
        RECT  3.110 1.145 3.400 1.375 ;
        RECT  3.010 0.985 3.110 1.375 ;
        RECT  2.740 1.145 3.010 1.375 ;
        RECT  2.620 1.010 2.740 1.375 ;
        RECT  2.370 1.145 2.620 1.375 ;
        RECT  2.250 1.010 2.370 1.375 ;
        RECT  1.555 1.145 2.250 1.375 ;
        RECT  1.475 0.760 1.555 1.375 ;
        RECT  1.210 1.145 1.475 1.375 ;
        RECT  1.090 1.120 1.210 1.375 ;
        RECT  0.340 1.145 1.090 1.375 ;
        RECT  0.220 1.010 0.340 1.375 ;
        RECT  0.000 1.145 0.220 1.375 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.195 0.805 3.305 1.075 ;
        RECT  3.185 0.355 3.285 0.485 ;
        RECT  3.185 0.805 3.195 0.905 ;
        RECT  2.815 0.355 2.835 0.480 ;
        RECT  2.820 0.805 2.835 1.075 ;
        RECT  4.515 0.195 4.585 1.005 ;
        RECT  4.490 0.195 4.515 0.355 ;
        RECT  4.490 0.845 4.515 1.005 ;
        RECT  4.010 0.845 4.490 0.915 ;
        RECT  3.710 0.990 4.210 1.060 ;
        RECT  3.920 0.530 4.010 0.915 ;
        RECT  3.850 0.210 3.940 0.315 ;
        RECT  3.780 0.210 3.850 0.910 ;
        RECT  2.345 0.210 3.780 0.280 ;
        RECT  3.640 0.350 3.710 1.060 ;
        RECT  3.570 0.350 3.640 0.420 ;
        RECT  3.600 0.905 3.640 1.060 ;
        RECT  2.740 0.550 2.830 0.640 ;
        RECT  2.670 0.550 2.740 0.940 ;
        RECT  1.950 0.870 2.670 0.940 ;
        RECT  2.465 0.350 2.560 0.800 ;
        RECT  2.135 0.730 2.465 0.800 ;
        RECT  2.265 0.210 2.345 0.660 ;
        RECT  1.770 0.210 2.265 0.280 ;
        RECT  2.060 0.350 2.135 0.800 ;
        RECT  1.870 0.350 1.950 0.940 ;
        RECT  1.700 0.210 1.770 0.905 ;
        RECT  1.640 0.210 1.700 0.300 ;
        RECT  1.640 0.835 1.700 0.905 ;
        RECT  1.385 0.530 1.630 0.650 ;
        RECT  1.370 0.530 1.385 0.880 ;
        RECT  0.810 0.980 1.385 1.050 ;
        RECT  1.295 0.350 1.370 0.880 ;
        RECT  0.960 0.840 1.030 0.910 ;
        RECT  0.960 0.310 1.000 0.410 ;
        RECT  0.890 0.195 0.960 0.910 ;
        RECT  0.350 0.195 0.890 0.265 ;
        RECT  0.740 0.350 0.810 1.050 ;
        RECT  0.720 0.350 0.740 0.860 ;
        RECT  0.685 0.730 0.720 0.860 ;
        RECT  0.570 0.995 0.660 1.065 ;
        RECT  0.500 0.870 0.570 1.065 ;
        RECT  0.485 0.350 0.560 0.800 ;
        RECT  0.130 0.870 0.500 0.940 ;
        RECT  0.105 0.870 0.130 1.050 ;
        RECT  0.105 0.300 0.120 0.440 ;
        RECT  0.035 0.300 0.105 1.050 ;
    END
END XOR4D4BWP40

END LIBRARY
